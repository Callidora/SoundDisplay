// Verilog netlist created by TD v5.0.19080
// Sun May 31 12:04:42 2020

`timescale 1ns / 1ps
module VGA_Demo  // source/rtl/VGA_Demo.v(2)
  (
  clk_24m,
  on_off,
  rst_n,
  vga_b,
  vga_clk,
  vga_de,
  vga_g,
  vga_hs,
  vga_r,
  vga_vs
  );

  input clk_24m;  // source/rtl/VGA_Demo.v(4)
  input [7:0] on_off;  // source/rtl/VGA_Demo.v(6)
  input rst_n;  // source/rtl/VGA_Demo.v(5)
  output [7:0] vga_b;  // source/rtl/VGA_Demo.v(17)
  output vga_clk;  // source/rtl/VGA_Demo.v(9)
  output vga_de;  // source/rtl/VGA_Demo.v(13)
  output [7:0] vga_g;  // source/rtl/VGA_Demo.v(16)
  output vga_hs;  // source/rtl/VGA_Demo.v(10)
  output [7:0] vga_r;  // source/rtl/VGA_Demo.v(15)
  output vga_vs;  // source/rtl/VGA_Demo.v(11)

  wire [23:0] lcd_data;  // source/rtl/VGA_Demo.v(23)
  wire [11:0] lcd_xpos;  // source/rtl/VGA_Demo.v(21)
  wire [11:0] lcd_ypos;  // source/rtl/VGA_Demo.v(22)
  wire [11:0] \u1_Driver/hcnt ;  // source/rtl/Driver.v(44)
  wire [11:0] \u1_Driver/n2 ;
  wire [12:0] \u1_Driver/n20 ;
  wire [12:0] \u1_Driver/n21 ;
  wire [11:0] \u1_Driver/n3 ;
  wire [11:0] \u1_Driver/n7 ;
  wire [11:0] \u1_Driver/n8 ;
  wire [11:0] \u1_Driver/vcnt ;  // source/rtl/Driver.v(45)
  wire [31:0] \u2_Display/counta ;  // source/rtl/Display.v(39)
  wire [31:0] \u2_Display/i ;  // source/rtl/Display.v(41)
  wire [31:0] \u2_Display/j ;  // source/rtl/Display.v(42)
  wire [30:0] \u2_Display/n ;  // source/rtl/Display.v(48)
  wire [31:0] \u2_Display/n1014 ;
  wire [31:0] \u2_Display/n102 ;
  wire [31:0] \u2_Display/n1049 ;
  wire [31:0] \u2_Display/n1084 ;
  wire [31:0] \u2_Display/n1119 ;
  wire [31:0] \u2_Display/n1154 ;
  wire [31:0] \u2_Display/n1189 ;
  wire [9:0] \u2_Display/n133 ;
  wire [9:0] \u2_Display/n134 ;
  wire [24:0] \u2_Display/n135 ;
  wire [31:0] \u2_Display/n137 ;
  wire [22:0] \u2_Display/n140 ;
  wire [31:0] \u2_Display/n143 ;
  wire [9:0] \u2_Display/n147 ;
  wire [31:0] \u2_Display/n1542 ;
  wire [31:0] \u2_Display/n1577 ;
  wire [31:0] \u2_Display/n1612 ;
  wire [31:0] \u2_Display/n1647 ;
  wire [31:0] \u2_Display/n1682 ;
  wire [31:0] \u2_Display/n1717 ;
  wire [31:0] \u2_Display/n1752 ;
  wire [31:0] \u2_Display/n1787 ;
  wire [31:0] \u2_Display/n1822 ;
  wire [31:0] \u2_Display/n1857 ;
  wire [31:0] \u2_Display/n1892 ;
  wire [31:0] \u2_Display/n1927 ;
  wire [9:0] \u2_Display/n196 ;
  wire [31:0] \u2_Display/n1962 ;
  wire [31:0] \u2_Display/n1997 ;
  wire [31:0] \u2_Display/n2032 ;
  wire [31:0] \u2_Display/n2067 ;
  wire [31:0] \u2_Display/n2102 ;
  wire [31:0] \u2_Display/n2137 ;
  wire [31:0] \u2_Display/n2172 ;
  wire [31:0] \u2_Display/n2207 ;
  wire [31:0] \u2_Display/n223 ;
  wire [31:0] \u2_Display/n2242 ;
  wire [31:0] \u2_Display/n226 ;
  wire [31:0] \u2_Display/n2277 ;
  wire [31:0] \u2_Display/n230 ;
  wire [31:0] \u2_Display/n231 ;
  wire [31:0] \u2_Display/n2312 ;
  wire [23:0] \u2_Display/n232 ;
  wire [31:0] \u2_Display/n234 ;
  wire [31:0] \u2_Display/n235 ;
  wire [23:0] \u2_Display/n236 ;
  wire [31:0] \u2_Display/n238 ;
  wire [31:0] \u2_Display/n239 ;
  wire [23:0] \u2_Display/n240 ;
  wire [31:0] \u2_Display/n2665 ;
  wire [31:0] \u2_Display/n2700 ;
  wire [31:0] \u2_Display/n2735 ;
  wire [31:0] \u2_Display/n2770 ;
  wire [31:0] \u2_Display/n2805 ;
  wire [31:0] \u2_Display/n2840 ;
  wire [31:0] \u2_Display/n2875 ;
  wire [31:0] \u2_Display/n2910 ;
  wire [31:0] \u2_Display/n2945 ;
  wire [31:0] \u2_Display/n2980 ;
  wire [31:0] \u2_Display/n3015 ;
  wire [31:0] \u2_Display/n3050 ;
  wire [31:0] \u2_Display/n3085 ;
  wire [31:0] \u2_Display/n3120 ;
  wire [31:0] \u2_Display/n3155 ;
  wire [31:0] \u2_Display/n3190 ;
  wire [31:0] \u2_Display/n3225 ;
  wire [31:0] \u2_Display/n3260 ;
  wire [31:0] \u2_Display/n3295 ;
  wire [31:0] \u2_Display/n3330 ;
  wire [31:0] \u2_Display/n3365 ;
  wire [31:0] \u2_Display/n3400 ;
  wire [31:0] \u2_Display/n3435 ;
  wire [30:0] \u2_Display/n37 ;
  wire [31:0] \u2_Display/n3788 ;
  wire [31:0] \u2_Display/n3823 ;
  wire [31:0] \u2_Display/n3858 ;
  wire [31:0] \u2_Display/n3893 ;
  wire [31:0] \u2_Display/n3928 ;
  wire [31:0] \u2_Display/n3963 ;
  wire [31:0] \u2_Display/n3998 ;
  wire [31:0] \u2_Display/n4033 ;
  wire [31:0] \u2_Display/n4068 ;
  wire [31:0] \u2_Display/n41 ;
  wire [31:0] \u2_Display/n4103 ;
  wire [31:0] \u2_Display/n4138 ;
  wire [31:0] \u2_Display/n4173 ;
  wire [31:0] \u2_Display/n419 ;
  wire [10:0] \u2_Display/n42 ;
  wire [31:0] \u2_Display/n4208 ;
  wire [31:0] \u2_Display/n4243 ;
  wire [31:0] \u2_Display/n4278 ;
  wire [23:0] \u2_Display/n43 ;
  wire [31:0] \u2_Display/n4313 ;
  wire [31:0] \u2_Display/n4348 ;
  wire [31:0] \u2_Display/n4383 ;
  wire [31:0] \u2_Display/n4418 ;
  wire [31:0] \u2_Display/n4453 ;
  wire [31:0] \u2_Display/n4488 ;
  wire [31:0] \u2_Display/n4523 ;
  wire [31:0] \u2_Display/n454 ;
  wire [31:0] \u2_Display/n4558 ;
  wire [31:0] \u2_Display/n489 ;
  wire [31:0] \u2_Display/n4911 ;
  wire [31:0] \u2_Display/n4946 ;
  wire [31:0] \u2_Display/n4981 ;
  wire [31:0] \u2_Display/n5016 ;
  wire [31:0] \u2_Display/n5051 ;
  wire [31:0] \u2_Display/n5086 ;
  wire [31:0] \u2_Display/n5121 ;
  wire [31:0] \u2_Display/n5156 ;
  wire [31:0] \u2_Display/n5191 ;
  wire [31:0] \u2_Display/n5226 ;
  wire [31:0] \u2_Display/n524 ;
  wire [31:0] \u2_Display/n5261 ;
  wire [31:0] \u2_Display/n5296 ;
  wire [31:0] \u2_Display/n5331 ;
  wire [31:0] \u2_Display/n5366 ;
  wire [31:0] \u2_Display/n5401 ;
  wire [31:0] \u2_Display/n5436 ;
  wire [31:0] \u2_Display/n5471 ;
  wire [31:0] \u2_Display/n5506 ;
  wire [31:0] \u2_Display/n5541 ;
  wire [31:0] \u2_Display/n5576 ;
  wire [31:0] \u2_Display/n559 ;
  wire [31:0] \u2_Display/n5611 ;
  wire [31:0] \u2_Display/n5646 ;
  wire [31:0] \u2_Display/n5681 ;
  wire [31:0] \u2_Display/n594 ;
  wire [31:0] \u2_Display/n629 ;
  wire [31:0] \u2_Display/n664 ;
  wire [31:0] \u2_Display/n6804 ;
  wire [31:0] \u2_Display/n699 ;
  wire [31:0] \u2_Display/n734 ;
  wire [31:0] \u2_Display/n769 ;
  wire [31:0] \u2_Display/n804 ;
  wire [31:0] \u2_Display/n839 ;
  wire [31:0] \u2_Display/n874 ;
  wire [31:0] \u2_Display/n909 ;
  wire [9:0] \u2_Display/n93 ;
  wire [24:0] \u2_Display/n94 ;
  wire [31:0] \u2_Display/n944 ;
  wire [31:0] \u2_Display/n96 ;
  wire [31:0] \u2_Display/n979 ;
  wire [22:0] \u2_Display/n99 ;
  wire clk_vga;  // source/rtl/VGA_Demo.v(20)
  wire \on_off[0]_neg ;
  wire \on_off[1]_neg ;
  wire \on_off[2]_neg ;
  wire \on_off[3]_neg ;
  wire \on_off[4]_neg ;
  wire \u0_PLL/n0 ;
  wire \u0_PLL/uut/clk0_buf ;  // al_ip/PLL.v(32)
  wire \u1_Driver/lcd_request ;  // source/rtl/Driver.v(46)
  wire \u1_Driver/n1 ;
  wire \u1_Driver/n10 ;
  wire \u1_Driver/n11 ;
  wire \u1_Driver/n12 ;
  wire \u1_Driver/n13 ;
  wire \u1_Driver/n14 ;
  wire \u1_Driver/n15 ;
  wire \u1_Driver/n16 ;
  wire \u1_Driver/n17 ;
  wire \u1_Driver/n18 ;
  wire \u1_Driver/n19 ;
  wire \u1_Driver/n4 ;
  wire \u1_Driver/n5 ;
  wire \u1_Driver/n6 ;
  wire \u2_Display/add2_2_co ;
  wire \u2_Display/add4_2_co ;
  wire \u2_Display/add5_2_co ;
  wire \u2_Display/add6_2_co ;
  wire \u2_Display/add7_2_co ;
  wire \u2_Display/clk1s ;  // source/rtl/Display.v(46)
  wire \u2_Display/mux10_b10_sel_is_2_o ;
  wire \u2_Display/mux11_b0_sel_is_0_o ;
  wire \u2_Display/mux13_b0_sel_is_2_o ;
  wire \u2_Display/mux17_b0_sel_is_2_o ;
  wire \u2_Display/mux17_b0_sel_is_2_o_neg ;
  wire \u2_Display/mux19_b0_sel_is_0_o ;
  wire \u2_Display/mux21_b0_sel_is_0_o ;
  wire \u2_Display/mux5_b0_sel_is_0_o ;
  wire \u2_Display/n100 ;
  wire \u2_Display/n1000 ;
  wire \u2_Display/n1001 ;
  wire \u2_Display/n1002 ;
  wire \u2_Display/n1003 ;
  wire \u2_Display/n1004 ;
  wire \u2_Display/n1005 ;
  wire \u2_Display/n1006 ;
  wire \u2_Display/n1007 ;
  wire \u2_Display/n1008 ;
  wire \u2_Display/n1009 ;
  wire \u2_Display/n101 ;
  wire \u2_Display/n1010 ;
  wire \u2_Display/n1011 ;
  wire \u2_Display/n1012 ;
  wire \u2_Display/n1013 ;
  wire \u2_Display/n1015 ;
  wire \u2_Display/n1016 ;
  wire \u2_Display/n1017 ;
  wire \u2_Display/n1018 ;
  wire \u2_Display/n1019 ;
  wire \u2_Display/n1020 ;
  wire \u2_Display/n1021 ;
  wire \u2_Display/n1022 ;
  wire \u2_Display/n1023 ;
  wire \u2_Display/n1024 ;
  wire \u2_Display/n1025 ;
  wire \u2_Display/n1026 ;
  wire \u2_Display/n1027 ;
  wire \u2_Display/n1028 ;
  wire \u2_Display/n1029 ;
  wire \u2_Display/n103 ;
  wire \u2_Display/n1030 ;
  wire \u2_Display/n1031 ;
  wire \u2_Display/n1032 ;
  wire \u2_Display/n1033 ;
  wire \u2_Display/n1034 ;
  wire \u2_Display/n1035 ;
  wire \u2_Display/n1036 ;
  wire \u2_Display/n1037 ;
  wire \u2_Display/n1038 ;
  wire \u2_Display/n1039 ;
  wire \u2_Display/n104 ;
  wire \u2_Display/n1040 ;
  wire \u2_Display/n1041 ;
  wire \u2_Display/n1042 ;
  wire \u2_Display/n1043 ;
  wire \u2_Display/n1044 ;
  wire \u2_Display/n1045 ;
  wire \u2_Display/n1046 ;
  wire \u2_Display/n1047 ;
  wire \u2_Display/n1048 ;
  wire \u2_Display/n1050 ;
  wire \u2_Display/n1051 ;
  wire \u2_Display/n1052 ;
  wire \u2_Display/n1053 ;
  wire \u2_Display/n1054 ;
  wire \u2_Display/n1055 ;
  wire \u2_Display/n1056 ;
  wire \u2_Display/n1057 ;
  wire \u2_Display/n1058 ;
  wire \u2_Display/n1059 ;
  wire \u2_Display/n1060 ;
  wire \u2_Display/n1061 ;
  wire \u2_Display/n1062 ;
  wire \u2_Display/n1063 ;
  wire \u2_Display/n1064 ;
  wire \u2_Display/n1065 ;
  wire \u2_Display/n1066 ;
  wire \u2_Display/n1067 ;
  wire \u2_Display/n1068 ;
  wire \u2_Display/n1069 ;
  wire \u2_Display/n1070 ;
  wire \u2_Display/n1071 ;
  wire \u2_Display/n1072 ;
  wire \u2_Display/n1073 ;
  wire \u2_Display/n1074 ;
  wire \u2_Display/n1075 ;
  wire \u2_Display/n1076 ;
  wire \u2_Display/n1077 ;
  wire \u2_Display/n1078 ;
  wire \u2_Display/n1079 ;
  wire \u2_Display/n1080 ;
  wire \u2_Display/n1081 ;
  wire \u2_Display/n1082 ;
  wire \u2_Display/n1083 ;
  wire \u2_Display/n1085 ;
  wire \u2_Display/n1086 ;
  wire \u2_Display/n1087 ;
  wire \u2_Display/n1088 ;
  wire \u2_Display/n1089 ;
  wire \u2_Display/n1090 ;
  wire \u2_Display/n1091 ;
  wire \u2_Display/n1092 ;
  wire \u2_Display/n1093 ;
  wire \u2_Display/n1094 ;
  wire \u2_Display/n1095 ;
  wire \u2_Display/n1096 ;
  wire \u2_Display/n1097 ;
  wire \u2_Display/n1098 ;
  wire \u2_Display/n1099 ;
  wire \u2_Display/n1100 ;
  wire \u2_Display/n1101 ;
  wire \u2_Display/n1102 ;
  wire \u2_Display/n1103 ;
  wire \u2_Display/n1104 ;
  wire \u2_Display/n1105 ;
  wire \u2_Display/n1106 ;
  wire \u2_Display/n1107 ;
  wire \u2_Display/n1108 ;
  wire \u2_Display/n1109 ;
  wire \u2_Display/n1110 ;
  wire \u2_Display/n1111 ;
  wire \u2_Display/n1112 ;
  wire \u2_Display/n1113 ;
  wire \u2_Display/n1114 ;
  wire \u2_Display/n1115 ;
  wire \u2_Display/n1116 ;
  wire \u2_Display/n1117 ;
  wire \u2_Display/n1118 ;
  wire \u2_Display/n1120 ;
  wire \u2_Display/n1121 ;
  wire \u2_Display/n1122 ;
  wire \u2_Display/n1123 ;
  wire \u2_Display/n1124 ;
  wire \u2_Display/n1125 ;
  wire \u2_Display/n1126 ;
  wire \u2_Display/n1127 ;
  wire \u2_Display/n1128 ;
  wire \u2_Display/n1129 ;
  wire \u2_Display/n1130 ;
  wire \u2_Display/n1131 ;
  wire \u2_Display/n1132 ;
  wire \u2_Display/n1133 ;
  wire \u2_Display/n1134 ;
  wire \u2_Display/n1135 ;
  wire \u2_Display/n1136 ;
  wire \u2_Display/n1137 ;
  wire \u2_Display/n1138 ;
  wire \u2_Display/n1139 ;
  wire \u2_Display/n1140 ;
  wire \u2_Display/n1141 ;
  wire \u2_Display/n1142 ;
  wire \u2_Display/n1143 ;
  wire \u2_Display/n1144 ;
  wire \u2_Display/n1145 ;
  wire \u2_Display/n1146 ;
  wire \u2_Display/n1147 ;
  wire \u2_Display/n1148 ;
  wire \u2_Display/n1149 ;
  wire \u2_Display/n1150 ;
  wire \u2_Display/n1151 ;
  wire \u2_Display/n1152 ;
  wire \u2_Display/n1153 ;
  wire \u2_Display/n1155 ;
  wire \u2_Display/n1156 ;
  wire \u2_Display/n1157 ;
  wire \u2_Display/n1158 ;
  wire \u2_Display/n1159 ;
  wire \u2_Display/n1160 ;
  wire \u2_Display/n1161 ;
  wire \u2_Display/n1162 ;
  wire \u2_Display/n1163 ;
  wire \u2_Display/n1164 ;
  wire \u2_Display/n1165 ;
  wire \u2_Display/n1166 ;
  wire \u2_Display/n1167 ;
  wire \u2_Display/n1168 ;
  wire \u2_Display/n1169 ;
  wire \u2_Display/n1170 ;
  wire \u2_Display/n1171 ;
  wire \u2_Display/n1172 ;
  wire \u2_Display/n1173 ;
  wire \u2_Display/n1174 ;
  wire \u2_Display/n1175 ;
  wire \u2_Display/n1176 ;
  wire \u2_Display/n1177 ;
  wire \u2_Display/n1178 ;
  wire \u2_Display/n1179 ;
  wire \u2_Display/n1180 ;
  wire \u2_Display/n1181 ;
  wire \u2_Display/n1182 ;
  wire \u2_Display/n1183 ;
  wire \u2_Display/n1184 ;
  wire \u2_Display/n1185 ;
  wire \u2_Display/n1186 ;
  wire \u2_Display/n1187 ;
  wire \u2_Display/n1188 ;
  wire \u2_Display/n136 ;
  wire \u2_Display/n138 ;
  wire \u2_Display/n139 ;
  wire \u2_Display/n141 ;
  wire \u2_Display/n142 ;
  wire \u2_Display/n144 ;
  wire \u2_Display/n145 ;
  wire \u2_Display/n1540 ;
  wire \u2_Display/n1541 ;
  wire \u2_Display/n1543 ;
  wire \u2_Display/n1544 ;
  wire \u2_Display/n1545 ;
  wire \u2_Display/n1546 ;
  wire \u2_Display/n1547 ;
  wire \u2_Display/n1548 ;
  wire \u2_Display/n1549 ;
  wire \u2_Display/n1550 ;
  wire \u2_Display/n1551 ;
  wire \u2_Display/n1552 ;
  wire \u2_Display/n1553 ;
  wire \u2_Display/n1554 ;
  wire \u2_Display/n1555 ;
  wire \u2_Display/n1556 ;
  wire \u2_Display/n1557 ;
  wire \u2_Display/n1558 ;
  wire \u2_Display/n1559 ;
  wire \u2_Display/n1560 ;
  wire \u2_Display/n1561 ;
  wire \u2_Display/n1562 ;
  wire \u2_Display/n1563 ;
  wire \u2_Display/n1564 ;
  wire \u2_Display/n1565 ;
  wire \u2_Display/n1566 ;
  wire \u2_Display/n1567 ;
  wire \u2_Display/n1568 ;
  wire \u2_Display/n1569 ;
  wire \u2_Display/n1570 ;
  wire \u2_Display/n1571 ;
  wire \u2_Display/n1572 ;
  wire \u2_Display/n1573 ;
  wire \u2_Display/n1574 ;
  wire \u2_Display/n1575 ;
  wire \u2_Display/n1576 ;
  wire \u2_Display/n1578 ;
  wire \u2_Display/n1579 ;
  wire \u2_Display/n1580 ;
  wire \u2_Display/n1581 ;
  wire \u2_Display/n1582 ;
  wire \u2_Display/n1583 ;
  wire \u2_Display/n1584 ;
  wire \u2_Display/n1585 ;
  wire \u2_Display/n1586 ;
  wire \u2_Display/n1587 ;
  wire \u2_Display/n1588 ;
  wire \u2_Display/n1589 ;
  wire \u2_Display/n1590 ;
  wire \u2_Display/n1591 ;
  wire \u2_Display/n1592 ;
  wire \u2_Display/n1593 ;
  wire \u2_Display/n1594 ;
  wire \u2_Display/n1595 ;
  wire \u2_Display/n1596 ;
  wire \u2_Display/n1597 ;
  wire \u2_Display/n1598 ;
  wire \u2_Display/n1599 ;
  wire \u2_Display/n1600 ;
  wire \u2_Display/n1601 ;
  wire \u2_Display/n1602 ;
  wire \u2_Display/n1603 ;
  wire \u2_Display/n1604 ;
  wire \u2_Display/n1605 ;
  wire \u2_Display/n1606 ;
  wire \u2_Display/n1607 ;
  wire \u2_Display/n1608 ;
  wire \u2_Display/n1609 ;
  wire \u2_Display/n1610 ;
  wire \u2_Display/n1611 ;
  wire \u2_Display/n1613 ;
  wire \u2_Display/n1614 ;
  wire \u2_Display/n1615 ;
  wire \u2_Display/n1616 ;
  wire \u2_Display/n1617 ;
  wire \u2_Display/n1618 ;
  wire \u2_Display/n1619 ;
  wire \u2_Display/n1620 ;
  wire \u2_Display/n1621 ;
  wire \u2_Display/n1622 ;
  wire \u2_Display/n1623 ;
  wire \u2_Display/n1624 ;
  wire \u2_Display/n1625 ;
  wire \u2_Display/n1626 ;
  wire \u2_Display/n1627 ;
  wire \u2_Display/n1628 ;
  wire \u2_Display/n1629 ;
  wire \u2_Display/n1630 ;
  wire \u2_Display/n1631 ;
  wire \u2_Display/n1632 ;
  wire \u2_Display/n1633 ;
  wire \u2_Display/n1634 ;
  wire \u2_Display/n1635 ;
  wire \u2_Display/n1636 ;
  wire \u2_Display/n1637 ;
  wire \u2_Display/n1638 ;
  wire \u2_Display/n1639 ;
  wire \u2_Display/n1640 ;
  wire \u2_Display/n1641 ;
  wire \u2_Display/n1642 ;
  wire \u2_Display/n1643 ;
  wire \u2_Display/n1644 ;
  wire \u2_Display/n1645 ;
  wire \u2_Display/n1646 ;
  wire \u2_Display/n1648 ;
  wire \u2_Display/n1649 ;
  wire \u2_Display/n1650 ;
  wire \u2_Display/n1651 ;
  wire \u2_Display/n1652 ;
  wire \u2_Display/n1653 ;
  wire \u2_Display/n1654 ;
  wire \u2_Display/n1655 ;
  wire \u2_Display/n1656 ;
  wire \u2_Display/n1657 ;
  wire \u2_Display/n1658 ;
  wire \u2_Display/n1659 ;
  wire \u2_Display/n1660 ;
  wire \u2_Display/n1661 ;
  wire \u2_Display/n1662 ;
  wire \u2_Display/n1663 ;
  wire \u2_Display/n1664 ;
  wire \u2_Display/n1665 ;
  wire \u2_Display/n1666 ;
  wire \u2_Display/n1667 ;
  wire \u2_Display/n1668 ;
  wire \u2_Display/n1669 ;
  wire \u2_Display/n1670 ;
  wire \u2_Display/n1671 ;
  wire \u2_Display/n1672 ;
  wire \u2_Display/n1673 ;
  wire \u2_Display/n1674 ;
  wire \u2_Display/n1675 ;
  wire \u2_Display/n1676 ;
  wire \u2_Display/n1677 ;
  wire \u2_Display/n1678 ;
  wire \u2_Display/n1679 ;
  wire \u2_Display/n1680 ;
  wire \u2_Display/n1681 ;
  wire \u2_Display/n1683 ;
  wire \u2_Display/n1684 ;
  wire \u2_Display/n1685 ;
  wire \u2_Display/n1686 ;
  wire \u2_Display/n1687 ;
  wire \u2_Display/n1688 ;
  wire \u2_Display/n1689 ;
  wire \u2_Display/n1690 ;
  wire \u2_Display/n1691 ;
  wire \u2_Display/n1692 ;
  wire \u2_Display/n1693 ;
  wire \u2_Display/n1694 ;
  wire \u2_Display/n1695 ;
  wire \u2_Display/n1696 ;
  wire \u2_Display/n1697 ;
  wire \u2_Display/n1698 ;
  wire \u2_Display/n1699 ;
  wire \u2_Display/n1700 ;
  wire \u2_Display/n1701 ;
  wire \u2_Display/n1702 ;
  wire \u2_Display/n1703 ;
  wire \u2_Display/n1704 ;
  wire \u2_Display/n1705 ;
  wire \u2_Display/n1706 ;
  wire \u2_Display/n1707 ;
  wire \u2_Display/n1708 ;
  wire \u2_Display/n1709 ;
  wire \u2_Display/n1710 ;
  wire \u2_Display/n1711 ;
  wire \u2_Display/n1712 ;
  wire \u2_Display/n1713 ;
  wire \u2_Display/n1714 ;
  wire \u2_Display/n1715 ;
  wire \u2_Display/n1716 ;
  wire \u2_Display/n1718 ;
  wire \u2_Display/n1719 ;
  wire \u2_Display/n1720 ;
  wire \u2_Display/n1721 ;
  wire \u2_Display/n1722 ;
  wire \u2_Display/n1723 ;
  wire \u2_Display/n1724 ;
  wire \u2_Display/n1725 ;
  wire \u2_Display/n1726 ;
  wire \u2_Display/n1727 ;
  wire \u2_Display/n1728 ;
  wire \u2_Display/n1729 ;
  wire \u2_Display/n1730 ;
  wire \u2_Display/n1731 ;
  wire \u2_Display/n1732 ;
  wire \u2_Display/n1733 ;
  wire \u2_Display/n1734 ;
  wire \u2_Display/n1735 ;
  wire \u2_Display/n1736 ;
  wire \u2_Display/n1737 ;
  wire \u2_Display/n1738 ;
  wire \u2_Display/n1739 ;
  wire \u2_Display/n1740 ;
  wire \u2_Display/n1741 ;
  wire \u2_Display/n1742 ;
  wire \u2_Display/n1743 ;
  wire \u2_Display/n1744 ;
  wire \u2_Display/n1745 ;
  wire \u2_Display/n1746 ;
  wire \u2_Display/n1747 ;
  wire \u2_Display/n1748 ;
  wire \u2_Display/n1749 ;
  wire \u2_Display/n1750 ;
  wire \u2_Display/n1751 ;
  wire \u2_Display/n1753 ;
  wire \u2_Display/n1754 ;
  wire \u2_Display/n1755 ;
  wire \u2_Display/n1756 ;
  wire \u2_Display/n1757 ;
  wire \u2_Display/n1758 ;
  wire \u2_Display/n1759 ;
  wire \u2_Display/n1760 ;
  wire \u2_Display/n1761 ;
  wire \u2_Display/n1762 ;
  wire \u2_Display/n1763 ;
  wire \u2_Display/n1764 ;
  wire \u2_Display/n1765 ;
  wire \u2_Display/n1766 ;
  wire \u2_Display/n1767 ;
  wire \u2_Display/n1768 ;
  wire \u2_Display/n1769 ;
  wire \u2_Display/n1770 ;
  wire \u2_Display/n1771 ;
  wire \u2_Display/n1772 ;
  wire \u2_Display/n1773 ;
  wire \u2_Display/n1774 ;
  wire \u2_Display/n1775 ;
  wire \u2_Display/n1776 ;
  wire \u2_Display/n1777 ;
  wire \u2_Display/n1778 ;
  wire \u2_Display/n1779 ;
  wire \u2_Display/n1780 ;
  wire \u2_Display/n1781 ;
  wire \u2_Display/n1782 ;
  wire \u2_Display/n1783 ;
  wire \u2_Display/n1784 ;
  wire \u2_Display/n1785 ;
  wire \u2_Display/n1786 ;
  wire \u2_Display/n1788 ;
  wire \u2_Display/n1789 ;
  wire \u2_Display/n1790 ;
  wire \u2_Display/n1791 ;
  wire \u2_Display/n1792 ;
  wire \u2_Display/n1793 ;
  wire \u2_Display/n1794 ;
  wire \u2_Display/n1795 ;
  wire \u2_Display/n1796 ;
  wire \u2_Display/n1797 ;
  wire \u2_Display/n1798 ;
  wire \u2_Display/n1799 ;
  wire \u2_Display/n1800 ;
  wire \u2_Display/n1801 ;
  wire \u2_Display/n1802 ;
  wire \u2_Display/n1803 ;
  wire \u2_Display/n1804 ;
  wire \u2_Display/n1805 ;
  wire \u2_Display/n1806 ;
  wire \u2_Display/n1807 ;
  wire \u2_Display/n1808 ;
  wire \u2_Display/n1809 ;
  wire \u2_Display/n1810 ;
  wire \u2_Display/n1811 ;
  wire \u2_Display/n1812 ;
  wire \u2_Display/n1813 ;
  wire \u2_Display/n1814 ;
  wire \u2_Display/n1815 ;
  wire \u2_Display/n1816 ;
  wire \u2_Display/n1817 ;
  wire \u2_Display/n1818 ;
  wire \u2_Display/n1819 ;
  wire \u2_Display/n1820 ;
  wire \u2_Display/n1821 ;
  wire \u2_Display/n1823 ;
  wire \u2_Display/n1824 ;
  wire \u2_Display/n1825 ;
  wire \u2_Display/n1826 ;
  wire \u2_Display/n1827 ;
  wire \u2_Display/n1828 ;
  wire \u2_Display/n1829 ;
  wire \u2_Display/n1830 ;
  wire \u2_Display/n1831 ;
  wire \u2_Display/n1832 ;
  wire \u2_Display/n1833 ;
  wire \u2_Display/n1834 ;
  wire \u2_Display/n1835 ;
  wire \u2_Display/n1836 ;
  wire \u2_Display/n1837 ;
  wire \u2_Display/n1838 ;
  wire \u2_Display/n1839 ;
  wire \u2_Display/n1840 ;
  wire \u2_Display/n1841 ;
  wire \u2_Display/n1842 ;
  wire \u2_Display/n1843 ;
  wire \u2_Display/n1844 ;
  wire \u2_Display/n1845 ;
  wire \u2_Display/n1846 ;
  wire \u2_Display/n1847 ;
  wire \u2_Display/n1848 ;
  wire \u2_Display/n1849 ;
  wire \u2_Display/n1850 ;
  wire \u2_Display/n1851 ;
  wire \u2_Display/n1852 ;
  wire \u2_Display/n1853 ;
  wire \u2_Display/n1854 ;
  wire \u2_Display/n1855 ;
  wire \u2_Display/n1856 ;
  wire \u2_Display/n1858 ;
  wire \u2_Display/n1859 ;
  wire \u2_Display/n1860 ;
  wire \u2_Display/n1861 ;
  wire \u2_Display/n1862 ;
  wire \u2_Display/n1863 ;
  wire \u2_Display/n1864 ;
  wire \u2_Display/n1865 ;
  wire \u2_Display/n1866 ;
  wire \u2_Display/n1867 ;
  wire \u2_Display/n1868 ;
  wire \u2_Display/n1869 ;
  wire \u2_Display/n1870 ;
  wire \u2_Display/n1871 ;
  wire \u2_Display/n1872 ;
  wire \u2_Display/n1873 ;
  wire \u2_Display/n1874 ;
  wire \u2_Display/n1875 ;
  wire \u2_Display/n1876 ;
  wire \u2_Display/n1877 ;
  wire \u2_Display/n1878 ;
  wire \u2_Display/n1879 ;
  wire \u2_Display/n1880 ;
  wire \u2_Display/n1881 ;
  wire \u2_Display/n1882 ;
  wire \u2_Display/n1883 ;
  wire \u2_Display/n1884 ;
  wire \u2_Display/n1885 ;
  wire \u2_Display/n1886 ;
  wire \u2_Display/n1887 ;
  wire \u2_Display/n1888 ;
  wire \u2_Display/n1889 ;
  wire \u2_Display/n1890 ;
  wire \u2_Display/n1891 ;
  wire \u2_Display/n1893 ;
  wire \u2_Display/n1894 ;
  wire \u2_Display/n1895 ;
  wire \u2_Display/n1896 ;
  wire \u2_Display/n1897 ;
  wire \u2_Display/n1898 ;
  wire \u2_Display/n1899 ;
  wire \u2_Display/n1900 ;
  wire \u2_Display/n1901 ;
  wire \u2_Display/n1902 ;
  wire \u2_Display/n1903 ;
  wire \u2_Display/n1904 ;
  wire \u2_Display/n1905 ;
  wire \u2_Display/n1906 ;
  wire \u2_Display/n1907 ;
  wire \u2_Display/n1908 ;
  wire \u2_Display/n1909 ;
  wire \u2_Display/n1910 ;
  wire \u2_Display/n1911 ;
  wire \u2_Display/n1912 ;
  wire \u2_Display/n1913 ;
  wire \u2_Display/n1914 ;
  wire \u2_Display/n1915 ;
  wire \u2_Display/n1916 ;
  wire \u2_Display/n1917 ;
  wire \u2_Display/n1918 ;
  wire \u2_Display/n1919 ;
  wire \u2_Display/n1920 ;
  wire \u2_Display/n1921 ;
  wire \u2_Display/n1922 ;
  wire \u2_Display/n1923 ;
  wire \u2_Display/n1924 ;
  wire \u2_Display/n1925 ;
  wire \u2_Display/n1926 ;
  wire \u2_Display/n1928 ;
  wire \u2_Display/n1929 ;
  wire \u2_Display/n1930 ;
  wire \u2_Display/n1931 ;
  wire \u2_Display/n1932 ;
  wire \u2_Display/n1933 ;
  wire \u2_Display/n1934 ;
  wire \u2_Display/n1935 ;
  wire \u2_Display/n1936 ;
  wire \u2_Display/n1937 ;
  wire \u2_Display/n1938 ;
  wire \u2_Display/n1939 ;
  wire \u2_Display/n1940 ;
  wire \u2_Display/n1941 ;
  wire \u2_Display/n1942 ;
  wire \u2_Display/n1943 ;
  wire \u2_Display/n1944 ;
  wire \u2_Display/n1945 ;
  wire \u2_Display/n1946 ;
  wire \u2_Display/n1947 ;
  wire \u2_Display/n1948 ;
  wire \u2_Display/n1949 ;
  wire \u2_Display/n1950 ;
  wire \u2_Display/n1951 ;
  wire \u2_Display/n1952 ;
  wire \u2_Display/n1953 ;
  wire \u2_Display/n1954 ;
  wire \u2_Display/n1955 ;
  wire \u2_Display/n1956 ;
  wire \u2_Display/n1957 ;
  wire \u2_Display/n1958 ;
  wire \u2_Display/n1959 ;
  wire \u2_Display/n1960 ;
  wire \u2_Display/n1961 ;
  wire \u2_Display/n1963 ;
  wire \u2_Display/n1964 ;
  wire \u2_Display/n1965 ;
  wire \u2_Display/n1966 ;
  wire \u2_Display/n1967 ;
  wire \u2_Display/n1968 ;
  wire \u2_Display/n1969 ;
  wire \u2_Display/n1970 ;
  wire \u2_Display/n1971 ;
  wire \u2_Display/n1972 ;
  wire \u2_Display/n1973 ;
  wire \u2_Display/n1974 ;
  wire \u2_Display/n1975 ;
  wire \u2_Display/n1976 ;
  wire \u2_Display/n1977 ;
  wire \u2_Display/n1978 ;
  wire \u2_Display/n1979 ;
  wire \u2_Display/n1980 ;
  wire \u2_Display/n1981 ;
  wire \u2_Display/n1982 ;
  wire \u2_Display/n1983 ;
  wire \u2_Display/n1984 ;
  wire \u2_Display/n1985 ;
  wire \u2_Display/n1986 ;
  wire \u2_Display/n1987 ;
  wire \u2_Display/n1988 ;
  wire \u2_Display/n1989 ;
  wire \u2_Display/n1990 ;
  wire \u2_Display/n1991 ;
  wire \u2_Display/n1992 ;
  wire \u2_Display/n1993 ;
  wire \u2_Display/n1994 ;
  wire \u2_Display/n1995 ;
  wire \u2_Display/n1996 ;
  wire \u2_Display/n1998 ;
  wire \u2_Display/n1999 ;
  wire \u2_Display/n2000 ;
  wire \u2_Display/n2001 ;
  wire \u2_Display/n2002 ;
  wire \u2_Display/n2003 ;
  wire \u2_Display/n2004 ;
  wire \u2_Display/n2005 ;
  wire \u2_Display/n2006 ;
  wire \u2_Display/n2007 ;
  wire \u2_Display/n2008 ;
  wire \u2_Display/n2009 ;
  wire \u2_Display/n2010 ;
  wire \u2_Display/n2011 ;
  wire \u2_Display/n2012 ;
  wire \u2_Display/n2013 ;
  wire \u2_Display/n2014 ;
  wire \u2_Display/n2015 ;
  wire \u2_Display/n2016 ;
  wire \u2_Display/n2017 ;
  wire \u2_Display/n2018 ;
  wire \u2_Display/n2019 ;
  wire \u2_Display/n2020 ;
  wire \u2_Display/n2021 ;
  wire \u2_Display/n2022 ;
  wire \u2_Display/n2023 ;
  wire \u2_Display/n2024 ;
  wire \u2_Display/n2025 ;
  wire \u2_Display/n2026 ;
  wire \u2_Display/n2027 ;
  wire \u2_Display/n2028 ;
  wire \u2_Display/n2029 ;
  wire \u2_Display/n2030 ;
  wire \u2_Display/n2031 ;
  wire \u2_Display/n2033 ;
  wire \u2_Display/n2034 ;
  wire \u2_Display/n2035 ;
  wire \u2_Display/n2036 ;
  wire \u2_Display/n2037 ;
  wire \u2_Display/n2038 ;
  wire \u2_Display/n2039 ;
  wire \u2_Display/n2040 ;
  wire \u2_Display/n2041 ;
  wire \u2_Display/n2042 ;
  wire \u2_Display/n2043 ;
  wire \u2_Display/n2044 ;
  wire \u2_Display/n2045 ;
  wire \u2_Display/n2046 ;
  wire \u2_Display/n2047 ;
  wire \u2_Display/n2048 ;
  wire \u2_Display/n2049 ;
  wire \u2_Display/n2050 ;
  wire \u2_Display/n2051 ;
  wire \u2_Display/n2052 ;
  wire \u2_Display/n2053 ;
  wire \u2_Display/n2054 ;
  wire \u2_Display/n2055 ;
  wire \u2_Display/n2056 ;
  wire \u2_Display/n2057 ;
  wire \u2_Display/n2058 ;
  wire \u2_Display/n2059 ;
  wire \u2_Display/n2060 ;
  wire \u2_Display/n2061 ;
  wire \u2_Display/n2062 ;
  wire \u2_Display/n2063 ;
  wire \u2_Display/n2064 ;
  wire \u2_Display/n2065 ;
  wire \u2_Display/n2066 ;
  wire \u2_Display/n2068 ;
  wire \u2_Display/n2069 ;
  wire \u2_Display/n2070 ;
  wire \u2_Display/n2071 ;
  wire \u2_Display/n2072 ;
  wire \u2_Display/n2073 ;
  wire \u2_Display/n2074 ;
  wire \u2_Display/n2075 ;
  wire \u2_Display/n2076 ;
  wire \u2_Display/n2077 ;
  wire \u2_Display/n2078 ;
  wire \u2_Display/n2079 ;
  wire \u2_Display/n2080 ;
  wire \u2_Display/n2081 ;
  wire \u2_Display/n2082 ;
  wire \u2_Display/n2083 ;
  wire \u2_Display/n2084 ;
  wire \u2_Display/n2085 ;
  wire \u2_Display/n2086 ;
  wire \u2_Display/n2087 ;
  wire \u2_Display/n2088 ;
  wire \u2_Display/n2089 ;
  wire \u2_Display/n2090 ;
  wire \u2_Display/n2091 ;
  wire \u2_Display/n2092 ;
  wire \u2_Display/n2093 ;
  wire \u2_Display/n2094 ;
  wire \u2_Display/n2095 ;
  wire \u2_Display/n2096 ;
  wire \u2_Display/n2097 ;
  wire \u2_Display/n2098 ;
  wire \u2_Display/n2099 ;
  wire \u2_Display/n2100 ;
  wire \u2_Display/n2101 ;
  wire \u2_Display/n2103 ;
  wire \u2_Display/n2104 ;
  wire \u2_Display/n2105 ;
  wire \u2_Display/n2106 ;
  wire \u2_Display/n2107 ;
  wire \u2_Display/n2108 ;
  wire \u2_Display/n2109 ;
  wire \u2_Display/n2110 ;
  wire \u2_Display/n2111 ;
  wire \u2_Display/n2112 ;
  wire \u2_Display/n2113 ;
  wire \u2_Display/n2114 ;
  wire \u2_Display/n2115 ;
  wire \u2_Display/n2116 ;
  wire \u2_Display/n2117 ;
  wire \u2_Display/n2118 ;
  wire \u2_Display/n2119 ;
  wire \u2_Display/n2120 ;
  wire \u2_Display/n2121 ;
  wire \u2_Display/n2122 ;
  wire \u2_Display/n2123 ;
  wire \u2_Display/n2124 ;
  wire \u2_Display/n2125 ;
  wire \u2_Display/n2126 ;
  wire \u2_Display/n2127 ;
  wire \u2_Display/n2128 ;
  wire \u2_Display/n2129 ;
  wire \u2_Display/n2130 ;
  wire \u2_Display/n2131 ;
  wire \u2_Display/n2132 ;
  wire \u2_Display/n2133 ;
  wire \u2_Display/n2134 ;
  wire \u2_Display/n2135 ;
  wire \u2_Display/n2136 ;
  wire \u2_Display/n2138 ;
  wire \u2_Display/n2139 ;
  wire \u2_Display/n2140 ;
  wire \u2_Display/n2141 ;
  wire \u2_Display/n2142 ;
  wire \u2_Display/n2143 ;
  wire \u2_Display/n2144 ;
  wire \u2_Display/n2145 ;
  wire \u2_Display/n2146 ;
  wire \u2_Display/n2147 ;
  wire \u2_Display/n2148 ;
  wire \u2_Display/n2149 ;
  wire \u2_Display/n2150 ;
  wire \u2_Display/n2151 ;
  wire \u2_Display/n2152 ;
  wire \u2_Display/n2153 ;
  wire \u2_Display/n2154 ;
  wire \u2_Display/n2155 ;
  wire \u2_Display/n2156 ;
  wire \u2_Display/n2157 ;
  wire \u2_Display/n2158 ;
  wire \u2_Display/n2159 ;
  wire \u2_Display/n2160 ;
  wire \u2_Display/n2161 ;
  wire \u2_Display/n2162 ;
  wire \u2_Display/n2163 ;
  wire \u2_Display/n2164 ;
  wire \u2_Display/n2165 ;
  wire \u2_Display/n2166 ;
  wire \u2_Display/n2167 ;
  wire \u2_Display/n2168 ;
  wire \u2_Display/n2169 ;
  wire \u2_Display/n2170 ;
  wire \u2_Display/n2171 ;
  wire \u2_Display/n2173 ;
  wire \u2_Display/n2174 ;
  wire \u2_Display/n2175 ;
  wire \u2_Display/n2176 ;
  wire \u2_Display/n2177 ;
  wire \u2_Display/n2178 ;
  wire \u2_Display/n2179 ;
  wire \u2_Display/n2180 ;
  wire \u2_Display/n2181 ;
  wire \u2_Display/n2182 ;
  wire \u2_Display/n2183 ;
  wire \u2_Display/n2184 ;
  wire \u2_Display/n2185 ;
  wire \u2_Display/n2186 ;
  wire \u2_Display/n2187 ;
  wire \u2_Display/n2188 ;
  wire \u2_Display/n2189 ;
  wire \u2_Display/n2190 ;
  wire \u2_Display/n2191 ;
  wire \u2_Display/n2192 ;
  wire \u2_Display/n2193 ;
  wire \u2_Display/n2194 ;
  wire \u2_Display/n2195 ;
  wire \u2_Display/n2196 ;
  wire \u2_Display/n2197 ;
  wire \u2_Display/n2198 ;
  wire \u2_Display/n2199 ;
  wire \u2_Display/n2200 ;
  wire \u2_Display/n2201 ;
  wire \u2_Display/n2202 ;
  wire \u2_Display/n2203 ;
  wire \u2_Display/n2204 ;
  wire \u2_Display/n2205 ;
  wire \u2_Display/n2206 ;
  wire \u2_Display/n2208 ;
  wire \u2_Display/n2209 ;
  wire \u2_Display/n2210 ;
  wire \u2_Display/n2211 ;
  wire \u2_Display/n2212 ;
  wire \u2_Display/n2213 ;
  wire \u2_Display/n2214 ;
  wire \u2_Display/n2215 ;
  wire \u2_Display/n2216 ;
  wire \u2_Display/n2217 ;
  wire \u2_Display/n2218 ;
  wire \u2_Display/n2219 ;
  wire \u2_Display/n2220 ;
  wire \u2_Display/n2221 ;
  wire \u2_Display/n2222 ;
  wire \u2_Display/n2223 ;
  wire \u2_Display/n2224 ;
  wire \u2_Display/n2225 ;
  wire \u2_Display/n2226 ;
  wire \u2_Display/n2227 ;
  wire \u2_Display/n2228 ;
  wire \u2_Display/n2229 ;
  wire \u2_Display/n2230 ;
  wire \u2_Display/n2231 ;
  wire \u2_Display/n2232 ;
  wire \u2_Display/n2233 ;
  wire \u2_Display/n2234 ;
  wire \u2_Display/n2235 ;
  wire \u2_Display/n2236 ;
  wire \u2_Display/n2237 ;
  wire \u2_Display/n2238 ;
  wire \u2_Display/n2239 ;
  wire \u2_Display/n2240 ;
  wire \u2_Display/n2241 ;
  wire \u2_Display/n2243 ;
  wire \u2_Display/n2244 ;
  wire \u2_Display/n2245 ;
  wire \u2_Display/n2246 ;
  wire \u2_Display/n2247 ;
  wire \u2_Display/n2248 ;
  wire \u2_Display/n2249 ;
  wire \u2_Display/n2250 ;
  wire \u2_Display/n2251 ;
  wire \u2_Display/n2252 ;
  wire \u2_Display/n2253 ;
  wire \u2_Display/n2254 ;
  wire \u2_Display/n2255 ;
  wire \u2_Display/n2256 ;
  wire \u2_Display/n2257 ;
  wire \u2_Display/n2258 ;
  wire \u2_Display/n2259 ;
  wire \u2_Display/n2260 ;
  wire \u2_Display/n2261 ;
  wire \u2_Display/n2262 ;
  wire \u2_Display/n2263 ;
  wire \u2_Display/n2264 ;
  wire \u2_Display/n2265 ;
  wire \u2_Display/n2266 ;
  wire \u2_Display/n2267 ;
  wire \u2_Display/n2268 ;
  wire \u2_Display/n2269 ;
  wire \u2_Display/n2270 ;
  wire \u2_Display/n2271 ;
  wire \u2_Display/n2272 ;
  wire \u2_Display/n2273 ;
  wire \u2_Display/n2274 ;
  wire \u2_Display/n2275 ;
  wire \u2_Display/n2276 ;
  wire \u2_Display/n2278 ;
  wire \u2_Display/n2279 ;
  wire \u2_Display/n2280 ;
  wire \u2_Display/n2281 ;
  wire \u2_Display/n2282 ;
  wire \u2_Display/n2283 ;
  wire \u2_Display/n2284 ;
  wire \u2_Display/n2285 ;
  wire \u2_Display/n2286 ;
  wire \u2_Display/n2287 ;
  wire \u2_Display/n2288 ;
  wire \u2_Display/n2289 ;
  wire \u2_Display/n2290 ;
  wire \u2_Display/n2291 ;
  wire \u2_Display/n2292 ;
  wire \u2_Display/n2293 ;
  wire \u2_Display/n2294 ;
  wire \u2_Display/n2295 ;
  wire \u2_Display/n2296 ;
  wire \u2_Display/n2297 ;
  wire \u2_Display/n2298 ;
  wire \u2_Display/n2299 ;
  wire \u2_Display/n2300 ;
  wire \u2_Display/n2301 ;
  wire \u2_Display/n2302 ;
  wire \u2_Display/n2303 ;
  wire \u2_Display/n2304 ;
  wire \u2_Display/n2305 ;
  wire \u2_Display/n2306 ;
  wire \u2_Display/n2307 ;
  wire \u2_Display/n2308 ;
  wire \u2_Display/n2309 ;
  wire \u2_Display/n2310 ;
  wire \u2_Display/n2311 ;
  wire \u2_Display/n2663 ;
  wire \u2_Display/n2664 ;
  wire \u2_Display/n2666 ;
  wire \u2_Display/n2667 ;
  wire \u2_Display/n2668 ;
  wire \u2_Display/n2669 ;
  wire \u2_Display/n2670 ;
  wire \u2_Display/n2671 ;
  wire \u2_Display/n2672 ;
  wire \u2_Display/n2673 ;
  wire \u2_Display/n2674 ;
  wire \u2_Display/n2675 ;
  wire \u2_Display/n2676 ;
  wire \u2_Display/n2677 ;
  wire \u2_Display/n2678 ;
  wire \u2_Display/n2679 ;
  wire \u2_Display/n2680 ;
  wire \u2_Display/n2681 ;
  wire \u2_Display/n2682 ;
  wire \u2_Display/n2683 ;
  wire \u2_Display/n2684 ;
  wire \u2_Display/n2685 ;
  wire \u2_Display/n2686 ;
  wire \u2_Display/n2687 ;
  wire \u2_Display/n2688 ;
  wire \u2_Display/n2689 ;
  wire \u2_Display/n2690 ;
  wire \u2_Display/n2691 ;
  wire \u2_Display/n2692 ;
  wire \u2_Display/n2693 ;
  wire \u2_Display/n2694 ;
  wire \u2_Display/n2695 ;
  wire \u2_Display/n2696 ;
  wire \u2_Display/n2697 ;
  wire \u2_Display/n2698 ;
  wire \u2_Display/n2699 ;
  wire \u2_Display/n2701 ;
  wire \u2_Display/n2702 ;
  wire \u2_Display/n2703 ;
  wire \u2_Display/n2704 ;
  wire \u2_Display/n2705 ;
  wire \u2_Display/n2706 ;
  wire \u2_Display/n2707 ;
  wire \u2_Display/n2708 ;
  wire \u2_Display/n2709 ;
  wire \u2_Display/n2710 ;
  wire \u2_Display/n2711 ;
  wire \u2_Display/n2712 ;
  wire \u2_Display/n2713 ;
  wire \u2_Display/n2714 ;
  wire \u2_Display/n2715 ;
  wire \u2_Display/n2716 ;
  wire \u2_Display/n2717 ;
  wire \u2_Display/n2718 ;
  wire \u2_Display/n2719 ;
  wire \u2_Display/n2720 ;
  wire \u2_Display/n2721 ;
  wire \u2_Display/n2722 ;
  wire \u2_Display/n2723 ;
  wire \u2_Display/n2724 ;
  wire \u2_Display/n2725 ;
  wire \u2_Display/n2726 ;
  wire \u2_Display/n2727 ;
  wire \u2_Display/n2728 ;
  wire \u2_Display/n2729 ;
  wire \u2_Display/n2730 ;
  wire \u2_Display/n2731 ;
  wire \u2_Display/n2732 ;
  wire \u2_Display/n2733 ;
  wire \u2_Display/n2734 ;
  wire \u2_Display/n2736 ;
  wire \u2_Display/n2737 ;
  wire \u2_Display/n2738 ;
  wire \u2_Display/n2739 ;
  wire \u2_Display/n2740 ;
  wire \u2_Display/n2741 ;
  wire \u2_Display/n2742 ;
  wire \u2_Display/n2743 ;
  wire \u2_Display/n2744 ;
  wire \u2_Display/n2745 ;
  wire \u2_Display/n2746 ;
  wire \u2_Display/n2747 ;
  wire \u2_Display/n2748 ;
  wire \u2_Display/n2749 ;
  wire \u2_Display/n2750 ;
  wire \u2_Display/n2751 ;
  wire \u2_Display/n2752 ;
  wire \u2_Display/n2753 ;
  wire \u2_Display/n2754 ;
  wire \u2_Display/n2755 ;
  wire \u2_Display/n2756 ;
  wire \u2_Display/n2757 ;
  wire \u2_Display/n2758 ;
  wire \u2_Display/n2759 ;
  wire \u2_Display/n2760 ;
  wire \u2_Display/n2761 ;
  wire \u2_Display/n2762 ;
  wire \u2_Display/n2763 ;
  wire \u2_Display/n2764 ;
  wire \u2_Display/n2765 ;
  wire \u2_Display/n2766 ;
  wire \u2_Display/n2767 ;
  wire \u2_Display/n2768 ;
  wire \u2_Display/n2769 ;
  wire \u2_Display/n2771 ;
  wire \u2_Display/n2772 ;
  wire \u2_Display/n2773 ;
  wire \u2_Display/n2774 ;
  wire \u2_Display/n2775 ;
  wire \u2_Display/n2776 ;
  wire \u2_Display/n2777 ;
  wire \u2_Display/n2778 ;
  wire \u2_Display/n2779 ;
  wire \u2_Display/n2780 ;
  wire \u2_Display/n2781 ;
  wire \u2_Display/n2782 ;
  wire \u2_Display/n2783 ;
  wire \u2_Display/n2784 ;
  wire \u2_Display/n2785 ;
  wire \u2_Display/n2786 ;
  wire \u2_Display/n2787 ;
  wire \u2_Display/n2788 ;
  wire \u2_Display/n2789 ;
  wire \u2_Display/n2790 ;
  wire \u2_Display/n2791 ;
  wire \u2_Display/n2792 ;
  wire \u2_Display/n2793 ;
  wire \u2_Display/n2794 ;
  wire \u2_Display/n2795 ;
  wire \u2_Display/n2796 ;
  wire \u2_Display/n2797 ;
  wire \u2_Display/n2798 ;
  wire \u2_Display/n2799 ;
  wire \u2_Display/n2800 ;
  wire \u2_Display/n2801 ;
  wire \u2_Display/n2802 ;
  wire \u2_Display/n2803 ;
  wire \u2_Display/n2804 ;
  wire \u2_Display/n2806 ;
  wire \u2_Display/n2807 ;
  wire \u2_Display/n2808 ;
  wire \u2_Display/n2809 ;
  wire \u2_Display/n2810 ;
  wire \u2_Display/n2811 ;
  wire \u2_Display/n2812 ;
  wire \u2_Display/n2813 ;
  wire \u2_Display/n2814 ;
  wire \u2_Display/n2815 ;
  wire \u2_Display/n2816 ;
  wire \u2_Display/n2817 ;
  wire \u2_Display/n2818 ;
  wire \u2_Display/n2819 ;
  wire \u2_Display/n2820 ;
  wire \u2_Display/n2821 ;
  wire \u2_Display/n2822 ;
  wire \u2_Display/n2823 ;
  wire \u2_Display/n2824 ;
  wire \u2_Display/n2825 ;
  wire \u2_Display/n2826 ;
  wire \u2_Display/n2827 ;
  wire \u2_Display/n2828 ;
  wire \u2_Display/n2829 ;
  wire \u2_Display/n2830 ;
  wire \u2_Display/n2831 ;
  wire \u2_Display/n2832 ;
  wire \u2_Display/n2833 ;
  wire \u2_Display/n2834 ;
  wire \u2_Display/n2835 ;
  wire \u2_Display/n2836 ;
  wire \u2_Display/n2837 ;
  wire \u2_Display/n2838 ;
  wire \u2_Display/n2839 ;
  wire \u2_Display/n2841 ;
  wire \u2_Display/n2842 ;
  wire \u2_Display/n2843 ;
  wire \u2_Display/n2844 ;
  wire \u2_Display/n2845 ;
  wire \u2_Display/n2846 ;
  wire \u2_Display/n2847 ;
  wire \u2_Display/n2848 ;
  wire \u2_Display/n2849 ;
  wire \u2_Display/n2850 ;
  wire \u2_Display/n2851 ;
  wire \u2_Display/n2852 ;
  wire \u2_Display/n2853 ;
  wire \u2_Display/n2854 ;
  wire \u2_Display/n2855 ;
  wire \u2_Display/n2856 ;
  wire \u2_Display/n2857 ;
  wire \u2_Display/n2858 ;
  wire \u2_Display/n2859 ;
  wire \u2_Display/n2860 ;
  wire \u2_Display/n2861 ;
  wire \u2_Display/n2862 ;
  wire \u2_Display/n2863 ;
  wire \u2_Display/n2864 ;
  wire \u2_Display/n2865 ;
  wire \u2_Display/n2866 ;
  wire \u2_Display/n2867 ;
  wire \u2_Display/n2868 ;
  wire \u2_Display/n2869 ;
  wire \u2_Display/n2870 ;
  wire \u2_Display/n2871 ;
  wire \u2_Display/n2872 ;
  wire \u2_Display/n2873 ;
  wire \u2_Display/n2874 ;
  wire \u2_Display/n2876 ;
  wire \u2_Display/n2877 ;
  wire \u2_Display/n2878 ;
  wire \u2_Display/n2879 ;
  wire \u2_Display/n2880 ;
  wire \u2_Display/n2881 ;
  wire \u2_Display/n2882 ;
  wire \u2_Display/n2883 ;
  wire \u2_Display/n2884 ;
  wire \u2_Display/n2885 ;
  wire \u2_Display/n2886 ;
  wire \u2_Display/n2887 ;
  wire \u2_Display/n2888 ;
  wire \u2_Display/n2889 ;
  wire \u2_Display/n2890 ;
  wire \u2_Display/n2891 ;
  wire \u2_Display/n2892 ;
  wire \u2_Display/n2893 ;
  wire \u2_Display/n2894 ;
  wire \u2_Display/n2895 ;
  wire \u2_Display/n2896 ;
  wire \u2_Display/n2897 ;
  wire \u2_Display/n2898 ;
  wire \u2_Display/n2899 ;
  wire \u2_Display/n2900 ;
  wire \u2_Display/n2901 ;
  wire \u2_Display/n2902 ;
  wire \u2_Display/n2903 ;
  wire \u2_Display/n2904 ;
  wire \u2_Display/n2905 ;
  wire \u2_Display/n2906 ;
  wire \u2_Display/n2907 ;
  wire \u2_Display/n2908 ;
  wire \u2_Display/n2909 ;
  wire \u2_Display/n2911 ;
  wire \u2_Display/n2912 ;
  wire \u2_Display/n2913 ;
  wire \u2_Display/n2914 ;
  wire \u2_Display/n2915 ;
  wire \u2_Display/n2916 ;
  wire \u2_Display/n2917 ;
  wire \u2_Display/n2918 ;
  wire \u2_Display/n2919 ;
  wire \u2_Display/n2920 ;
  wire \u2_Display/n2921 ;
  wire \u2_Display/n2922 ;
  wire \u2_Display/n2923 ;
  wire \u2_Display/n2924 ;
  wire \u2_Display/n2925 ;
  wire \u2_Display/n2926 ;
  wire \u2_Display/n2927 ;
  wire \u2_Display/n2928 ;
  wire \u2_Display/n2929 ;
  wire \u2_Display/n2930 ;
  wire \u2_Display/n2931 ;
  wire \u2_Display/n2932 ;
  wire \u2_Display/n2933 ;
  wire \u2_Display/n2934 ;
  wire \u2_Display/n2935 ;
  wire \u2_Display/n2936 ;
  wire \u2_Display/n2937 ;
  wire \u2_Display/n2938 ;
  wire \u2_Display/n2939 ;
  wire \u2_Display/n2940 ;
  wire \u2_Display/n2941 ;
  wire \u2_Display/n2942 ;
  wire \u2_Display/n2943 ;
  wire \u2_Display/n2944 ;
  wire \u2_Display/n2946 ;
  wire \u2_Display/n2947 ;
  wire \u2_Display/n2948 ;
  wire \u2_Display/n2949 ;
  wire \u2_Display/n2950 ;
  wire \u2_Display/n2951 ;
  wire \u2_Display/n2952 ;
  wire \u2_Display/n2953 ;
  wire \u2_Display/n2954 ;
  wire \u2_Display/n2955 ;
  wire \u2_Display/n2956 ;
  wire \u2_Display/n2957 ;
  wire \u2_Display/n2958 ;
  wire \u2_Display/n2959 ;
  wire \u2_Display/n2960 ;
  wire \u2_Display/n2961 ;
  wire \u2_Display/n2962 ;
  wire \u2_Display/n2963 ;
  wire \u2_Display/n2964 ;
  wire \u2_Display/n2965 ;
  wire \u2_Display/n2966 ;
  wire \u2_Display/n2967 ;
  wire \u2_Display/n2968 ;
  wire \u2_Display/n2969 ;
  wire \u2_Display/n2970 ;
  wire \u2_Display/n2971 ;
  wire \u2_Display/n2972 ;
  wire \u2_Display/n2973 ;
  wire \u2_Display/n2974 ;
  wire \u2_Display/n2975 ;
  wire \u2_Display/n2976 ;
  wire \u2_Display/n2977 ;
  wire \u2_Display/n2978 ;
  wire \u2_Display/n2979 ;
  wire \u2_Display/n2981 ;
  wire \u2_Display/n2982 ;
  wire \u2_Display/n2983 ;
  wire \u2_Display/n2984 ;
  wire \u2_Display/n2985 ;
  wire \u2_Display/n2986 ;
  wire \u2_Display/n2987 ;
  wire \u2_Display/n2988 ;
  wire \u2_Display/n2989 ;
  wire \u2_Display/n2990 ;
  wire \u2_Display/n2991 ;
  wire \u2_Display/n2992 ;
  wire \u2_Display/n2993 ;
  wire \u2_Display/n2994 ;
  wire \u2_Display/n2995 ;
  wire \u2_Display/n2996 ;
  wire \u2_Display/n2997 ;
  wire \u2_Display/n2998 ;
  wire \u2_Display/n2999 ;
  wire \u2_Display/n3000 ;
  wire \u2_Display/n3001 ;
  wire \u2_Display/n3002 ;
  wire \u2_Display/n3003 ;
  wire \u2_Display/n3004 ;
  wire \u2_Display/n3005 ;
  wire \u2_Display/n3006 ;
  wire \u2_Display/n3007 ;
  wire \u2_Display/n3008 ;
  wire \u2_Display/n3009 ;
  wire \u2_Display/n3010 ;
  wire \u2_Display/n3011 ;
  wire \u2_Display/n3012 ;
  wire \u2_Display/n3013 ;
  wire \u2_Display/n3014 ;
  wire \u2_Display/n3016 ;
  wire \u2_Display/n3017 ;
  wire \u2_Display/n3018 ;
  wire \u2_Display/n3019 ;
  wire \u2_Display/n3020 ;
  wire \u2_Display/n3021 ;
  wire \u2_Display/n3022 ;
  wire \u2_Display/n3023 ;
  wire \u2_Display/n3024 ;
  wire \u2_Display/n3025 ;
  wire \u2_Display/n3026 ;
  wire \u2_Display/n3027 ;
  wire \u2_Display/n3028 ;
  wire \u2_Display/n3029 ;
  wire \u2_Display/n3030 ;
  wire \u2_Display/n3031 ;
  wire \u2_Display/n3032 ;
  wire \u2_Display/n3033 ;
  wire \u2_Display/n3034 ;
  wire \u2_Display/n3035 ;
  wire \u2_Display/n3036 ;
  wire \u2_Display/n3037 ;
  wire \u2_Display/n3038 ;
  wire \u2_Display/n3039 ;
  wire \u2_Display/n3040 ;
  wire \u2_Display/n3041 ;
  wire \u2_Display/n3042 ;
  wire \u2_Display/n3043 ;
  wire \u2_Display/n3044 ;
  wire \u2_Display/n3045 ;
  wire \u2_Display/n3046 ;
  wire \u2_Display/n3047 ;
  wire \u2_Display/n3048 ;
  wire \u2_Display/n3049 ;
  wire \u2_Display/n3051 ;
  wire \u2_Display/n3052 ;
  wire \u2_Display/n3053 ;
  wire \u2_Display/n3054 ;
  wire \u2_Display/n3055 ;
  wire \u2_Display/n3056 ;
  wire \u2_Display/n3057 ;
  wire \u2_Display/n3058 ;
  wire \u2_Display/n3059 ;
  wire \u2_Display/n3060 ;
  wire \u2_Display/n3061 ;
  wire \u2_Display/n3062 ;
  wire \u2_Display/n3063 ;
  wire \u2_Display/n3064 ;
  wire \u2_Display/n3065 ;
  wire \u2_Display/n3066 ;
  wire \u2_Display/n3067 ;
  wire \u2_Display/n3068 ;
  wire \u2_Display/n3069 ;
  wire \u2_Display/n3070 ;
  wire \u2_Display/n3071 ;
  wire \u2_Display/n3072 ;
  wire \u2_Display/n3073 ;
  wire \u2_Display/n3074 ;
  wire \u2_Display/n3075 ;
  wire \u2_Display/n3076 ;
  wire \u2_Display/n3077 ;
  wire \u2_Display/n3078 ;
  wire \u2_Display/n3079 ;
  wire \u2_Display/n3080 ;
  wire \u2_Display/n3081 ;
  wire \u2_Display/n3082 ;
  wire \u2_Display/n3083 ;
  wire \u2_Display/n3084 ;
  wire \u2_Display/n3086 ;
  wire \u2_Display/n3087 ;
  wire \u2_Display/n3088 ;
  wire \u2_Display/n3089 ;
  wire \u2_Display/n3090 ;
  wire \u2_Display/n3091 ;
  wire \u2_Display/n3092 ;
  wire \u2_Display/n3093 ;
  wire \u2_Display/n3094 ;
  wire \u2_Display/n3095 ;
  wire \u2_Display/n3096 ;
  wire \u2_Display/n3097 ;
  wire \u2_Display/n3098 ;
  wire \u2_Display/n3099 ;
  wire \u2_Display/n3100 ;
  wire \u2_Display/n3101 ;
  wire \u2_Display/n3102 ;
  wire \u2_Display/n3103 ;
  wire \u2_Display/n3104 ;
  wire \u2_Display/n3105 ;
  wire \u2_Display/n3106 ;
  wire \u2_Display/n3107 ;
  wire \u2_Display/n3108 ;
  wire \u2_Display/n3109 ;
  wire \u2_Display/n3110 ;
  wire \u2_Display/n3111 ;
  wire \u2_Display/n3112 ;
  wire \u2_Display/n3113 ;
  wire \u2_Display/n3114 ;
  wire \u2_Display/n3115 ;
  wire \u2_Display/n3116 ;
  wire \u2_Display/n3117 ;
  wire \u2_Display/n3118 ;
  wire \u2_Display/n3119 ;
  wire \u2_Display/n3121 ;
  wire \u2_Display/n3122 ;
  wire \u2_Display/n3123 ;
  wire \u2_Display/n3124 ;
  wire \u2_Display/n3125 ;
  wire \u2_Display/n3126 ;
  wire \u2_Display/n3127 ;
  wire \u2_Display/n3128 ;
  wire \u2_Display/n3129 ;
  wire \u2_Display/n3130 ;
  wire \u2_Display/n3131 ;
  wire \u2_Display/n3132 ;
  wire \u2_Display/n3133 ;
  wire \u2_Display/n3134 ;
  wire \u2_Display/n3135 ;
  wire \u2_Display/n3136 ;
  wire \u2_Display/n3137 ;
  wire \u2_Display/n3138 ;
  wire \u2_Display/n3139 ;
  wire \u2_Display/n3140 ;
  wire \u2_Display/n3141 ;
  wire \u2_Display/n3142 ;
  wire \u2_Display/n3143 ;
  wire \u2_Display/n3144 ;
  wire \u2_Display/n3145 ;
  wire \u2_Display/n3146 ;
  wire \u2_Display/n3147 ;
  wire \u2_Display/n3148 ;
  wire \u2_Display/n3149 ;
  wire \u2_Display/n3150 ;
  wire \u2_Display/n3151 ;
  wire \u2_Display/n3152 ;
  wire \u2_Display/n3153 ;
  wire \u2_Display/n3154 ;
  wire \u2_Display/n3156 ;
  wire \u2_Display/n3157 ;
  wire \u2_Display/n3158 ;
  wire \u2_Display/n3159 ;
  wire \u2_Display/n3160 ;
  wire \u2_Display/n3161 ;
  wire \u2_Display/n3162 ;
  wire \u2_Display/n3163 ;
  wire \u2_Display/n3164 ;
  wire \u2_Display/n3165 ;
  wire \u2_Display/n3166 ;
  wire \u2_Display/n3167 ;
  wire \u2_Display/n3168 ;
  wire \u2_Display/n3169 ;
  wire \u2_Display/n3170 ;
  wire \u2_Display/n3171 ;
  wire \u2_Display/n3172 ;
  wire \u2_Display/n3173 ;
  wire \u2_Display/n3174 ;
  wire \u2_Display/n3175 ;
  wire \u2_Display/n3176 ;
  wire \u2_Display/n3177 ;
  wire \u2_Display/n3178 ;
  wire \u2_Display/n3179 ;
  wire \u2_Display/n3180 ;
  wire \u2_Display/n3181 ;
  wire \u2_Display/n3182 ;
  wire \u2_Display/n3183 ;
  wire \u2_Display/n3184 ;
  wire \u2_Display/n3185 ;
  wire \u2_Display/n3186 ;
  wire \u2_Display/n3187 ;
  wire \u2_Display/n3188 ;
  wire \u2_Display/n3189 ;
  wire \u2_Display/n3191 ;
  wire \u2_Display/n3192 ;
  wire \u2_Display/n3193 ;
  wire \u2_Display/n3194 ;
  wire \u2_Display/n3195 ;
  wire \u2_Display/n3196 ;
  wire \u2_Display/n3197 ;
  wire \u2_Display/n3198 ;
  wire \u2_Display/n3199 ;
  wire \u2_Display/n3200 ;
  wire \u2_Display/n3201 ;
  wire \u2_Display/n3202 ;
  wire \u2_Display/n3203 ;
  wire \u2_Display/n3204 ;
  wire \u2_Display/n3205 ;
  wire \u2_Display/n3206 ;
  wire \u2_Display/n3207 ;
  wire \u2_Display/n3208 ;
  wire \u2_Display/n3209 ;
  wire \u2_Display/n3210 ;
  wire \u2_Display/n3211 ;
  wire \u2_Display/n3212 ;
  wire \u2_Display/n3213 ;
  wire \u2_Display/n3214 ;
  wire \u2_Display/n3215 ;
  wire \u2_Display/n3216 ;
  wire \u2_Display/n3217 ;
  wire \u2_Display/n3218 ;
  wire \u2_Display/n3219 ;
  wire \u2_Display/n3220 ;
  wire \u2_Display/n3221 ;
  wire \u2_Display/n3222 ;
  wire \u2_Display/n3223 ;
  wire \u2_Display/n3224 ;
  wire \u2_Display/n3226 ;
  wire \u2_Display/n3227 ;
  wire \u2_Display/n3228 ;
  wire \u2_Display/n3229 ;
  wire \u2_Display/n3230 ;
  wire \u2_Display/n3231 ;
  wire \u2_Display/n3232 ;
  wire \u2_Display/n3233 ;
  wire \u2_Display/n3234 ;
  wire \u2_Display/n3235 ;
  wire \u2_Display/n3236 ;
  wire \u2_Display/n3237 ;
  wire \u2_Display/n3238 ;
  wire \u2_Display/n3239 ;
  wire \u2_Display/n3240 ;
  wire \u2_Display/n3241 ;
  wire \u2_Display/n3242 ;
  wire \u2_Display/n3243 ;
  wire \u2_Display/n3244 ;
  wire \u2_Display/n3245 ;
  wire \u2_Display/n3246 ;
  wire \u2_Display/n3247 ;
  wire \u2_Display/n3248 ;
  wire \u2_Display/n3249 ;
  wire \u2_Display/n3250 ;
  wire \u2_Display/n3251 ;
  wire \u2_Display/n3252 ;
  wire \u2_Display/n3253 ;
  wire \u2_Display/n3254 ;
  wire \u2_Display/n3255 ;
  wire \u2_Display/n3256 ;
  wire \u2_Display/n3257 ;
  wire \u2_Display/n3258 ;
  wire \u2_Display/n3259 ;
  wire \u2_Display/n3261 ;
  wire \u2_Display/n3262 ;
  wire \u2_Display/n3263 ;
  wire \u2_Display/n3264 ;
  wire \u2_Display/n3265 ;
  wire \u2_Display/n3266 ;
  wire \u2_Display/n3267 ;
  wire \u2_Display/n3268 ;
  wire \u2_Display/n3269 ;
  wire \u2_Display/n3270 ;
  wire \u2_Display/n3271 ;
  wire \u2_Display/n3272 ;
  wire \u2_Display/n3273 ;
  wire \u2_Display/n3274 ;
  wire \u2_Display/n3275 ;
  wire \u2_Display/n3276 ;
  wire \u2_Display/n3277 ;
  wire \u2_Display/n3278 ;
  wire \u2_Display/n3279 ;
  wire \u2_Display/n3280 ;
  wire \u2_Display/n3281 ;
  wire \u2_Display/n3282 ;
  wire \u2_Display/n3283 ;
  wire \u2_Display/n3284 ;
  wire \u2_Display/n3285 ;
  wire \u2_Display/n3286 ;
  wire \u2_Display/n3287 ;
  wire \u2_Display/n3288 ;
  wire \u2_Display/n3289 ;
  wire \u2_Display/n3290 ;
  wire \u2_Display/n3291 ;
  wire \u2_Display/n3292 ;
  wire \u2_Display/n3293 ;
  wire \u2_Display/n3294 ;
  wire \u2_Display/n3296 ;
  wire \u2_Display/n3297 ;
  wire \u2_Display/n3298 ;
  wire \u2_Display/n3299 ;
  wire \u2_Display/n3300 ;
  wire \u2_Display/n3301 ;
  wire \u2_Display/n3302 ;
  wire \u2_Display/n3303 ;
  wire \u2_Display/n3304 ;
  wire \u2_Display/n3305 ;
  wire \u2_Display/n3306 ;
  wire \u2_Display/n3307 ;
  wire \u2_Display/n3308 ;
  wire \u2_Display/n3309 ;
  wire \u2_Display/n3310 ;
  wire \u2_Display/n3311 ;
  wire \u2_Display/n3312 ;
  wire \u2_Display/n3313 ;
  wire \u2_Display/n3314 ;
  wire \u2_Display/n3315 ;
  wire \u2_Display/n3316 ;
  wire \u2_Display/n3317 ;
  wire \u2_Display/n3318 ;
  wire \u2_Display/n3319 ;
  wire \u2_Display/n3320 ;
  wire \u2_Display/n3321 ;
  wire \u2_Display/n3322 ;
  wire \u2_Display/n3323 ;
  wire \u2_Display/n3324 ;
  wire \u2_Display/n3325 ;
  wire \u2_Display/n3326 ;
  wire \u2_Display/n3327 ;
  wire \u2_Display/n3328 ;
  wire \u2_Display/n3329 ;
  wire \u2_Display/n3331 ;
  wire \u2_Display/n3332 ;
  wire \u2_Display/n3333 ;
  wire \u2_Display/n3334 ;
  wire \u2_Display/n3335 ;
  wire \u2_Display/n3336 ;
  wire \u2_Display/n3337 ;
  wire \u2_Display/n3338 ;
  wire \u2_Display/n3339 ;
  wire \u2_Display/n3340 ;
  wire \u2_Display/n3341 ;
  wire \u2_Display/n3342 ;
  wire \u2_Display/n3343 ;
  wire \u2_Display/n3344 ;
  wire \u2_Display/n3345 ;
  wire \u2_Display/n3346 ;
  wire \u2_Display/n3347 ;
  wire \u2_Display/n3348 ;
  wire \u2_Display/n3349 ;
  wire \u2_Display/n3350 ;
  wire \u2_Display/n3351 ;
  wire \u2_Display/n3352 ;
  wire \u2_Display/n3353 ;
  wire \u2_Display/n3354 ;
  wire \u2_Display/n3355 ;
  wire \u2_Display/n3356 ;
  wire \u2_Display/n3357 ;
  wire \u2_Display/n3358 ;
  wire \u2_Display/n3359 ;
  wire \u2_Display/n3360 ;
  wire \u2_Display/n3361 ;
  wire \u2_Display/n3362 ;
  wire \u2_Display/n3363 ;
  wire \u2_Display/n3364 ;
  wire \u2_Display/n3366 ;
  wire \u2_Display/n3367 ;
  wire \u2_Display/n3368 ;
  wire \u2_Display/n3369 ;
  wire \u2_Display/n3370 ;
  wire \u2_Display/n3371 ;
  wire \u2_Display/n3372 ;
  wire \u2_Display/n3373 ;
  wire \u2_Display/n3374 ;
  wire \u2_Display/n3375 ;
  wire \u2_Display/n3376 ;
  wire \u2_Display/n3377 ;
  wire \u2_Display/n3378 ;
  wire \u2_Display/n3379 ;
  wire \u2_Display/n3380 ;
  wire \u2_Display/n3381 ;
  wire \u2_Display/n3382 ;
  wire \u2_Display/n3383 ;
  wire \u2_Display/n3384 ;
  wire \u2_Display/n3385 ;
  wire \u2_Display/n3386 ;
  wire \u2_Display/n3387 ;
  wire \u2_Display/n3388 ;
  wire \u2_Display/n3389 ;
  wire \u2_Display/n3390 ;
  wire \u2_Display/n3391 ;
  wire \u2_Display/n3392 ;
  wire \u2_Display/n3393 ;
  wire \u2_Display/n3394 ;
  wire \u2_Display/n3395 ;
  wire \u2_Display/n3396 ;
  wire \u2_Display/n3397 ;
  wire \u2_Display/n3398 ;
  wire \u2_Display/n3399 ;
  wire \u2_Display/n3401 ;
  wire \u2_Display/n3402 ;
  wire \u2_Display/n3403 ;
  wire \u2_Display/n3404 ;
  wire \u2_Display/n3405 ;
  wire \u2_Display/n3406 ;
  wire \u2_Display/n3407 ;
  wire \u2_Display/n3408 ;
  wire \u2_Display/n3409 ;
  wire \u2_Display/n3410 ;
  wire \u2_Display/n3411 ;
  wire \u2_Display/n3412 ;
  wire \u2_Display/n3413 ;
  wire \u2_Display/n3414 ;
  wire \u2_Display/n3415 ;
  wire \u2_Display/n3416 ;
  wire \u2_Display/n3417 ;
  wire \u2_Display/n3418 ;
  wire \u2_Display/n3419 ;
  wire \u2_Display/n3420 ;
  wire \u2_Display/n3421 ;
  wire \u2_Display/n3422 ;
  wire \u2_Display/n3423 ;
  wire \u2_Display/n3424 ;
  wire \u2_Display/n3425 ;
  wire \u2_Display/n3426 ;
  wire \u2_Display/n3427 ;
  wire \u2_Display/n3428 ;
  wire \u2_Display/n3429 ;
  wire \u2_Display/n3430 ;
  wire \u2_Display/n3431 ;
  wire \u2_Display/n3432 ;
  wire \u2_Display/n3433 ;
  wire \u2_Display/n3434 ;
  wire \u2_Display/n35 ;
  wire \u2_Display/n36 ;
  wire \u2_Display/n3786 ;
  wire \u2_Display/n3787 ;
  wire \u2_Display/n3789 ;
  wire \u2_Display/n3790 ;
  wire \u2_Display/n3791 ;
  wire \u2_Display/n3792 ;
  wire \u2_Display/n3793 ;
  wire \u2_Display/n3794 ;
  wire \u2_Display/n3795 ;
  wire \u2_Display/n3796 ;
  wire \u2_Display/n3797 ;
  wire \u2_Display/n3798 ;
  wire \u2_Display/n3799 ;
  wire \u2_Display/n3800 ;
  wire \u2_Display/n3801 ;
  wire \u2_Display/n3802 ;
  wire \u2_Display/n3803 ;
  wire \u2_Display/n3804 ;
  wire \u2_Display/n3805 ;
  wire \u2_Display/n3806 ;
  wire \u2_Display/n3807 ;
  wire \u2_Display/n3808 ;
  wire \u2_Display/n3809 ;
  wire \u2_Display/n3810 ;
  wire \u2_Display/n3811 ;
  wire \u2_Display/n3812 ;
  wire \u2_Display/n3813 ;
  wire \u2_Display/n3814 ;
  wire \u2_Display/n3815 ;
  wire \u2_Display/n3816 ;
  wire \u2_Display/n3817 ;
  wire \u2_Display/n3818 ;
  wire \u2_Display/n3819 ;
  wire \u2_Display/n3820 ;
  wire \u2_Display/n3821 ;
  wire \u2_Display/n3822 ;
  wire \u2_Display/n3824 ;
  wire \u2_Display/n3825 ;
  wire \u2_Display/n3826 ;
  wire \u2_Display/n3827 ;
  wire \u2_Display/n3828 ;
  wire \u2_Display/n3829 ;
  wire \u2_Display/n3830 ;
  wire \u2_Display/n3831 ;
  wire \u2_Display/n3832 ;
  wire \u2_Display/n3833 ;
  wire \u2_Display/n3834 ;
  wire \u2_Display/n3835 ;
  wire \u2_Display/n3836 ;
  wire \u2_Display/n3837 ;
  wire \u2_Display/n3838 ;
  wire \u2_Display/n3839 ;
  wire \u2_Display/n3840 ;
  wire \u2_Display/n3841 ;
  wire \u2_Display/n3842 ;
  wire \u2_Display/n3843 ;
  wire \u2_Display/n3844 ;
  wire \u2_Display/n3845 ;
  wire \u2_Display/n3846 ;
  wire \u2_Display/n3847 ;
  wire \u2_Display/n3848 ;
  wire \u2_Display/n3849 ;
  wire \u2_Display/n3850 ;
  wire \u2_Display/n3851 ;
  wire \u2_Display/n3852 ;
  wire \u2_Display/n3853 ;
  wire \u2_Display/n3854 ;
  wire \u2_Display/n3855 ;
  wire \u2_Display/n3856 ;
  wire \u2_Display/n3857 ;
  wire \u2_Display/n3859 ;
  wire \u2_Display/n3860 ;
  wire \u2_Display/n3861 ;
  wire \u2_Display/n3862 ;
  wire \u2_Display/n3863 ;
  wire \u2_Display/n3864 ;
  wire \u2_Display/n3865 ;
  wire \u2_Display/n3866 ;
  wire \u2_Display/n3867 ;
  wire \u2_Display/n3868 ;
  wire \u2_Display/n3869 ;
  wire \u2_Display/n3870 ;
  wire \u2_Display/n3871 ;
  wire \u2_Display/n3872 ;
  wire \u2_Display/n3873 ;
  wire \u2_Display/n3874 ;
  wire \u2_Display/n3875 ;
  wire \u2_Display/n3876 ;
  wire \u2_Display/n3877 ;
  wire \u2_Display/n3878 ;
  wire \u2_Display/n3879 ;
  wire \u2_Display/n3880 ;
  wire \u2_Display/n3881 ;
  wire \u2_Display/n3882 ;
  wire \u2_Display/n3883 ;
  wire \u2_Display/n3884 ;
  wire \u2_Display/n3885 ;
  wire \u2_Display/n3886 ;
  wire \u2_Display/n3887 ;
  wire \u2_Display/n3888 ;
  wire \u2_Display/n3889 ;
  wire \u2_Display/n3890 ;
  wire \u2_Display/n3891 ;
  wire \u2_Display/n3892 ;
  wire \u2_Display/n3894 ;
  wire \u2_Display/n3895 ;
  wire \u2_Display/n3896 ;
  wire \u2_Display/n3897 ;
  wire \u2_Display/n3898 ;
  wire \u2_Display/n3899 ;
  wire \u2_Display/n3900 ;
  wire \u2_Display/n3901 ;
  wire \u2_Display/n3902 ;
  wire \u2_Display/n3903 ;
  wire \u2_Display/n3904 ;
  wire \u2_Display/n3905 ;
  wire \u2_Display/n3906 ;
  wire \u2_Display/n3907 ;
  wire \u2_Display/n3908 ;
  wire \u2_Display/n3909 ;
  wire \u2_Display/n3910 ;
  wire \u2_Display/n3911 ;
  wire \u2_Display/n3912 ;
  wire \u2_Display/n3913 ;
  wire \u2_Display/n3914 ;
  wire \u2_Display/n3915 ;
  wire \u2_Display/n3916 ;
  wire \u2_Display/n3917 ;
  wire \u2_Display/n3918 ;
  wire \u2_Display/n3919 ;
  wire \u2_Display/n3920 ;
  wire \u2_Display/n3921 ;
  wire \u2_Display/n3922 ;
  wire \u2_Display/n3923 ;
  wire \u2_Display/n3924 ;
  wire \u2_Display/n3925 ;
  wire \u2_Display/n3926 ;
  wire \u2_Display/n3927 ;
  wire \u2_Display/n3929 ;
  wire \u2_Display/n3930 ;
  wire \u2_Display/n3931 ;
  wire \u2_Display/n3932 ;
  wire \u2_Display/n3933 ;
  wire \u2_Display/n3934 ;
  wire \u2_Display/n3935 ;
  wire \u2_Display/n3936 ;
  wire \u2_Display/n3937 ;
  wire \u2_Display/n3938 ;
  wire \u2_Display/n3939 ;
  wire \u2_Display/n3940 ;
  wire \u2_Display/n3941 ;
  wire \u2_Display/n3942 ;
  wire \u2_Display/n3943 ;
  wire \u2_Display/n3944 ;
  wire \u2_Display/n3945 ;
  wire \u2_Display/n3946 ;
  wire \u2_Display/n3947 ;
  wire \u2_Display/n3948 ;
  wire \u2_Display/n3949 ;
  wire \u2_Display/n3950 ;
  wire \u2_Display/n3951 ;
  wire \u2_Display/n3952 ;
  wire \u2_Display/n3953 ;
  wire \u2_Display/n3954 ;
  wire \u2_Display/n3955 ;
  wire \u2_Display/n3956 ;
  wire \u2_Display/n3957 ;
  wire \u2_Display/n3958 ;
  wire \u2_Display/n3959 ;
  wire \u2_Display/n3960 ;
  wire \u2_Display/n3961 ;
  wire \u2_Display/n3962 ;
  wire \u2_Display/n3964 ;
  wire \u2_Display/n3965 ;
  wire \u2_Display/n3966 ;
  wire \u2_Display/n3967 ;
  wire \u2_Display/n3968 ;
  wire \u2_Display/n3969 ;
  wire \u2_Display/n3970 ;
  wire \u2_Display/n3971 ;
  wire \u2_Display/n3972 ;
  wire \u2_Display/n3973 ;
  wire \u2_Display/n3974 ;
  wire \u2_Display/n3975 ;
  wire \u2_Display/n3976 ;
  wire \u2_Display/n3977 ;
  wire \u2_Display/n3978 ;
  wire \u2_Display/n3979 ;
  wire \u2_Display/n3980 ;
  wire \u2_Display/n3981 ;
  wire \u2_Display/n3982 ;
  wire \u2_Display/n3983 ;
  wire \u2_Display/n3984 ;
  wire \u2_Display/n3985 ;
  wire \u2_Display/n3986 ;
  wire \u2_Display/n3987 ;
  wire \u2_Display/n3988 ;
  wire \u2_Display/n3989 ;
  wire \u2_Display/n3990 ;
  wire \u2_Display/n3991 ;
  wire \u2_Display/n3992 ;
  wire \u2_Display/n3993 ;
  wire \u2_Display/n3994 ;
  wire \u2_Display/n3995 ;
  wire \u2_Display/n3996 ;
  wire \u2_Display/n3997 ;
  wire \u2_Display/n3999 ;
  wire \u2_Display/n4000 ;
  wire \u2_Display/n4001 ;
  wire \u2_Display/n4002 ;
  wire \u2_Display/n4003 ;
  wire \u2_Display/n4004 ;
  wire \u2_Display/n4005 ;
  wire \u2_Display/n4006 ;
  wire \u2_Display/n4007 ;
  wire \u2_Display/n4008 ;
  wire \u2_Display/n4009 ;
  wire \u2_Display/n4010 ;
  wire \u2_Display/n4011 ;
  wire \u2_Display/n4012 ;
  wire \u2_Display/n4013 ;
  wire \u2_Display/n4014 ;
  wire \u2_Display/n4015 ;
  wire \u2_Display/n4016 ;
  wire \u2_Display/n4017 ;
  wire \u2_Display/n4018 ;
  wire \u2_Display/n4019 ;
  wire \u2_Display/n4020 ;
  wire \u2_Display/n4021 ;
  wire \u2_Display/n4022 ;
  wire \u2_Display/n4023 ;
  wire \u2_Display/n4024 ;
  wire \u2_Display/n4025 ;
  wire \u2_Display/n4026 ;
  wire \u2_Display/n4027 ;
  wire \u2_Display/n4028 ;
  wire \u2_Display/n4029 ;
  wire \u2_Display/n4030 ;
  wire \u2_Display/n4031 ;
  wire \u2_Display/n4032 ;
  wire \u2_Display/n4034 ;
  wire \u2_Display/n4035 ;
  wire \u2_Display/n4036 ;
  wire \u2_Display/n4037 ;
  wire \u2_Display/n4038 ;
  wire \u2_Display/n4039 ;
  wire \u2_Display/n4040 ;
  wire \u2_Display/n4041 ;
  wire \u2_Display/n4042 ;
  wire \u2_Display/n4043 ;
  wire \u2_Display/n4044 ;
  wire \u2_Display/n4045 ;
  wire \u2_Display/n4046 ;
  wire \u2_Display/n4047 ;
  wire \u2_Display/n4048 ;
  wire \u2_Display/n4049 ;
  wire \u2_Display/n4050 ;
  wire \u2_Display/n4051 ;
  wire \u2_Display/n4052 ;
  wire \u2_Display/n4053 ;
  wire \u2_Display/n4054 ;
  wire \u2_Display/n4055 ;
  wire \u2_Display/n4056 ;
  wire \u2_Display/n4057 ;
  wire \u2_Display/n4058 ;
  wire \u2_Display/n4059 ;
  wire \u2_Display/n4060 ;
  wire \u2_Display/n4061 ;
  wire \u2_Display/n4062 ;
  wire \u2_Display/n4063 ;
  wire \u2_Display/n4064 ;
  wire \u2_Display/n4065 ;
  wire \u2_Display/n4066 ;
  wire \u2_Display/n4067 ;
  wire \u2_Display/n4069 ;
  wire \u2_Display/n4070 ;
  wire \u2_Display/n4071 ;
  wire \u2_Display/n4072 ;
  wire \u2_Display/n4073 ;
  wire \u2_Display/n4074 ;
  wire \u2_Display/n4075 ;
  wire \u2_Display/n4076 ;
  wire \u2_Display/n4077 ;
  wire \u2_Display/n4078 ;
  wire \u2_Display/n4079 ;
  wire \u2_Display/n4080 ;
  wire \u2_Display/n4081 ;
  wire \u2_Display/n4082 ;
  wire \u2_Display/n4083 ;
  wire \u2_Display/n4084 ;
  wire \u2_Display/n4085 ;
  wire \u2_Display/n4086 ;
  wire \u2_Display/n4087 ;
  wire \u2_Display/n4088 ;
  wire \u2_Display/n4089 ;
  wire \u2_Display/n4090 ;
  wire \u2_Display/n4091 ;
  wire \u2_Display/n4092 ;
  wire \u2_Display/n4093 ;
  wire \u2_Display/n4094 ;
  wire \u2_Display/n4095 ;
  wire \u2_Display/n4096 ;
  wire \u2_Display/n4097 ;
  wire \u2_Display/n4098 ;
  wire \u2_Display/n4099 ;
  wire \u2_Display/n4100 ;
  wire \u2_Display/n4101 ;
  wire \u2_Display/n4102 ;
  wire \u2_Display/n4104 ;
  wire \u2_Display/n4105 ;
  wire \u2_Display/n4106 ;
  wire \u2_Display/n4107 ;
  wire \u2_Display/n4108 ;
  wire \u2_Display/n4109 ;
  wire \u2_Display/n4110 ;
  wire \u2_Display/n4111 ;
  wire \u2_Display/n4112 ;
  wire \u2_Display/n4113 ;
  wire \u2_Display/n4114 ;
  wire \u2_Display/n4115 ;
  wire \u2_Display/n4116 ;
  wire \u2_Display/n4117 ;
  wire \u2_Display/n4118 ;
  wire \u2_Display/n4119 ;
  wire \u2_Display/n4120 ;
  wire \u2_Display/n4121 ;
  wire \u2_Display/n4122 ;
  wire \u2_Display/n4123 ;
  wire \u2_Display/n4124 ;
  wire \u2_Display/n4125 ;
  wire \u2_Display/n4126 ;
  wire \u2_Display/n4127 ;
  wire \u2_Display/n4128 ;
  wire \u2_Display/n4129 ;
  wire \u2_Display/n4130 ;
  wire \u2_Display/n4131 ;
  wire \u2_Display/n4132 ;
  wire \u2_Display/n4133 ;
  wire \u2_Display/n4134 ;
  wire \u2_Display/n4135 ;
  wire \u2_Display/n4136 ;
  wire \u2_Display/n4137 ;
  wire \u2_Display/n4139 ;
  wire \u2_Display/n4140 ;
  wire \u2_Display/n4141 ;
  wire \u2_Display/n4142 ;
  wire \u2_Display/n4143 ;
  wire \u2_Display/n4144 ;
  wire \u2_Display/n4145 ;
  wire \u2_Display/n4146 ;
  wire \u2_Display/n4147 ;
  wire \u2_Display/n4148 ;
  wire \u2_Display/n4149 ;
  wire \u2_Display/n4150 ;
  wire \u2_Display/n4151 ;
  wire \u2_Display/n4152 ;
  wire \u2_Display/n4153 ;
  wire \u2_Display/n4154 ;
  wire \u2_Display/n4155 ;
  wire \u2_Display/n4156 ;
  wire \u2_Display/n4157 ;
  wire \u2_Display/n4158 ;
  wire \u2_Display/n4159 ;
  wire \u2_Display/n4160 ;
  wire \u2_Display/n4161 ;
  wire \u2_Display/n4162 ;
  wire \u2_Display/n4163 ;
  wire \u2_Display/n4164 ;
  wire \u2_Display/n4165 ;
  wire \u2_Display/n4166 ;
  wire \u2_Display/n4167 ;
  wire \u2_Display/n4168 ;
  wire \u2_Display/n4169 ;
  wire \u2_Display/n417 ;
  wire \u2_Display/n4170 ;
  wire \u2_Display/n4171 ;
  wire \u2_Display/n4172 ;
  wire \u2_Display/n4174 ;
  wire \u2_Display/n4175 ;
  wire \u2_Display/n4176 ;
  wire \u2_Display/n4177 ;
  wire \u2_Display/n4178 ;
  wire \u2_Display/n4179 ;
  wire \u2_Display/n418 ;
  wire \u2_Display/n4180 ;
  wire \u2_Display/n4181 ;
  wire \u2_Display/n4182 ;
  wire \u2_Display/n4183 ;
  wire \u2_Display/n4184 ;
  wire \u2_Display/n4185 ;
  wire \u2_Display/n4186 ;
  wire \u2_Display/n4187 ;
  wire \u2_Display/n4188 ;
  wire \u2_Display/n4189 ;
  wire \u2_Display/n4190 ;
  wire \u2_Display/n4191 ;
  wire \u2_Display/n4192 ;
  wire \u2_Display/n4193 ;
  wire \u2_Display/n4194 ;
  wire \u2_Display/n4195 ;
  wire \u2_Display/n4196 ;
  wire \u2_Display/n4197 ;
  wire \u2_Display/n4198 ;
  wire \u2_Display/n4199 ;
  wire \u2_Display/n420 ;
  wire \u2_Display/n4200 ;
  wire \u2_Display/n4201 ;
  wire \u2_Display/n4202 ;
  wire \u2_Display/n4203 ;
  wire \u2_Display/n4204 ;
  wire \u2_Display/n4205 ;
  wire \u2_Display/n4206 ;
  wire \u2_Display/n4207 ;
  wire \u2_Display/n4209 ;
  wire \u2_Display/n421 ;
  wire \u2_Display/n4210 ;
  wire \u2_Display/n4211 ;
  wire \u2_Display/n4212 ;
  wire \u2_Display/n4213 ;
  wire \u2_Display/n4214 ;
  wire \u2_Display/n4215 ;
  wire \u2_Display/n4216 ;
  wire \u2_Display/n4217 ;
  wire \u2_Display/n4218 ;
  wire \u2_Display/n4219 ;
  wire \u2_Display/n422 ;
  wire \u2_Display/n4220 ;
  wire \u2_Display/n4221 ;
  wire \u2_Display/n4222 ;
  wire \u2_Display/n4223 ;
  wire \u2_Display/n4224 ;
  wire \u2_Display/n4225 ;
  wire \u2_Display/n4226 ;
  wire \u2_Display/n4227 ;
  wire \u2_Display/n4228 ;
  wire \u2_Display/n4229 ;
  wire \u2_Display/n423 ;
  wire \u2_Display/n4230 ;
  wire \u2_Display/n4231 ;
  wire \u2_Display/n4232 ;
  wire \u2_Display/n4233 ;
  wire \u2_Display/n4234 ;
  wire \u2_Display/n4235 ;
  wire \u2_Display/n4236 ;
  wire \u2_Display/n4237 ;
  wire \u2_Display/n4238 ;
  wire \u2_Display/n4239 ;
  wire \u2_Display/n424 ;
  wire \u2_Display/n4240 ;
  wire \u2_Display/n4241 ;
  wire \u2_Display/n4242 ;
  wire \u2_Display/n4244 ;
  wire \u2_Display/n4245 ;
  wire \u2_Display/n4246 ;
  wire \u2_Display/n4247 ;
  wire \u2_Display/n4248 ;
  wire \u2_Display/n4249 ;
  wire \u2_Display/n425 ;
  wire \u2_Display/n4250 ;
  wire \u2_Display/n4251 ;
  wire \u2_Display/n4252 ;
  wire \u2_Display/n4253 ;
  wire \u2_Display/n4254 ;
  wire \u2_Display/n4255 ;
  wire \u2_Display/n4256 ;
  wire \u2_Display/n4257 ;
  wire \u2_Display/n4258 ;
  wire \u2_Display/n4259 ;
  wire \u2_Display/n426 ;
  wire \u2_Display/n4260 ;
  wire \u2_Display/n4261 ;
  wire \u2_Display/n4262 ;
  wire \u2_Display/n4263 ;
  wire \u2_Display/n4264 ;
  wire \u2_Display/n4265 ;
  wire \u2_Display/n4266 ;
  wire \u2_Display/n4267 ;
  wire \u2_Display/n4268 ;
  wire \u2_Display/n4269 ;
  wire \u2_Display/n427 ;
  wire \u2_Display/n4270 ;
  wire \u2_Display/n4271 ;
  wire \u2_Display/n4272 ;
  wire \u2_Display/n4273 ;
  wire \u2_Display/n4274 ;
  wire \u2_Display/n4275 ;
  wire \u2_Display/n4276 ;
  wire \u2_Display/n4277 ;
  wire \u2_Display/n4279 ;
  wire \u2_Display/n428 ;
  wire \u2_Display/n4280 ;
  wire \u2_Display/n4281 ;
  wire \u2_Display/n4282 ;
  wire \u2_Display/n4283 ;
  wire \u2_Display/n4284 ;
  wire \u2_Display/n4285 ;
  wire \u2_Display/n4286 ;
  wire \u2_Display/n4287 ;
  wire \u2_Display/n4288 ;
  wire \u2_Display/n4289 ;
  wire \u2_Display/n429 ;
  wire \u2_Display/n4290 ;
  wire \u2_Display/n4291 ;
  wire \u2_Display/n4292 ;
  wire \u2_Display/n4293 ;
  wire \u2_Display/n4294 ;
  wire \u2_Display/n4295 ;
  wire \u2_Display/n4296 ;
  wire \u2_Display/n4297 ;
  wire \u2_Display/n4298 ;
  wire \u2_Display/n4299 ;
  wire \u2_Display/n430 ;
  wire \u2_Display/n4300 ;
  wire \u2_Display/n4301 ;
  wire \u2_Display/n4302 ;
  wire \u2_Display/n4303 ;
  wire \u2_Display/n4304 ;
  wire \u2_Display/n4305 ;
  wire \u2_Display/n4306 ;
  wire \u2_Display/n4307 ;
  wire \u2_Display/n4308 ;
  wire \u2_Display/n4309 ;
  wire \u2_Display/n431 ;
  wire \u2_Display/n4310 ;
  wire \u2_Display/n4311 ;
  wire \u2_Display/n4312 ;
  wire \u2_Display/n4314 ;
  wire \u2_Display/n4315 ;
  wire \u2_Display/n4316 ;
  wire \u2_Display/n4317 ;
  wire \u2_Display/n4318 ;
  wire \u2_Display/n4319 ;
  wire \u2_Display/n432 ;
  wire \u2_Display/n4320 ;
  wire \u2_Display/n4321 ;
  wire \u2_Display/n4322 ;
  wire \u2_Display/n4323 ;
  wire \u2_Display/n4324 ;
  wire \u2_Display/n4325 ;
  wire \u2_Display/n4326 ;
  wire \u2_Display/n4327 ;
  wire \u2_Display/n4328 ;
  wire \u2_Display/n4329 ;
  wire \u2_Display/n433 ;
  wire \u2_Display/n4330 ;
  wire \u2_Display/n4331 ;
  wire \u2_Display/n4332 ;
  wire \u2_Display/n4333 ;
  wire \u2_Display/n4334 ;
  wire \u2_Display/n4335 ;
  wire \u2_Display/n4336 ;
  wire \u2_Display/n4337 ;
  wire \u2_Display/n4338 ;
  wire \u2_Display/n4339 ;
  wire \u2_Display/n434 ;
  wire \u2_Display/n4340 ;
  wire \u2_Display/n4341 ;
  wire \u2_Display/n4342 ;
  wire \u2_Display/n4343 ;
  wire \u2_Display/n4344 ;
  wire \u2_Display/n4345 ;
  wire \u2_Display/n4346 ;
  wire \u2_Display/n4347 ;
  wire \u2_Display/n4349 ;
  wire \u2_Display/n435 ;
  wire \u2_Display/n4350 ;
  wire \u2_Display/n4351 ;
  wire \u2_Display/n4352 ;
  wire \u2_Display/n4353 ;
  wire \u2_Display/n4354 ;
  wire \u2_Display/n4355 ;
  wire \u2_Display/n4356 ;
  wire \u2_Display/n4357 ;
  wire \u2_Display/n4358 ;
  wire \u2_Display/n4359 ;
  wire \u2_Display/n436 ;
  wire \u2_Display/n4360 ;
  wire \u2_Display/n4361 ;
  wire \u2_Display/n4362 ;
  wire \u2_Display/n4363 ;
  wire \u2_Display/n4364 ;
  wire \u2_Display/n4365 ;
  wire \u2_Display/n4366 ;
  wire \u2_Display/n4367 ;
  wire \u2_Display/n4368 ;
  wire \u2_Display/n4369 ;
  wire \u2_Display/n437 ;
  wire \u2_Display/n4370 ;
  wire \u2_Display/n4371 ;
  wire \u2_Display/n4372 ;
  wire \u2_Display/n4373 ;
  wire \u2_Display/n4374 ;
  wire \u2_Display/n4375 ;
  wire \u2_Display/n4376 ;
  wire \u2_Display/n4377 ;
  wire \u2_Display/n4378 ;
  wire \u2_Display/n4379 ;
  wire \u2_Display/n438 ;
  wire \u2_Display/n4380 ;
  wire \u2_Display/n4381 ;
  wire \u2_Display/n4382 ;
  wire \u2_Display/n4384 ;
  wire \u2_Display/n4385 ;
  wire \u2_Display/n4386 ;
  wire \u2_Display/n4387 ;
  wire \u2_Display/n4388 ;
  wire \u2_Display/n4389 ;
  wire \u2_Display/n439 ;
  wire \u2_Display/n4390 ;
  wire \u2_Display/n4391 ;
  wire \u2_Display/n4392 ;
  wire \u2_Display/n4393 ;
  wire \u2_Display/n4394 ;
  wire \u2_Display/n4395 ;
  wire \u2_Display/n4396 ;
  wire \u2_Display/n4397 ;
  wire \u2_Display/n4398 ;
  wire \u2_Display/n4399 ;
  wire \u2_Display/n44 ;
  wire \u2_Display/n440 ;
  wire \u2_Display/n4400 ;
  wire \u2_Display/n4401 ;
  wire \u2_Display/n4402 ;
  wire \u2_Display/n4403 ;
  wire \u2_Display/n4404 ;
  wire \u2_Display/n4405 ;
  wire \u2_Display/n4406 ;
  wire \u2_Display/n4407 ;
  wire \u2_Display/n4408 ;
  wire \u2_Display/n4409 ;
  wire \u2_Display/n441 ;
  wire \u2_Display/n4410 ;
  wire \u2_Display/n4411 ;
  wire \u2_Display/n4412 ;
  wire \u2_Display/n4413 ;
  wire \u2_Display/n4414 ;
  wire \u2_Display/n4415 ;
  wire \u2_Display/n4416 ;
  wire \u2_Display/n4417 ;
  wire \u2_Display/n4419 ;
  wire \u2_Display/n442 ;
  wire \u2_Display/n4420 ;
  wire \u2_Display/n4421 ;
  wire \u2_Display/n4422 ;
  wire \u2_Display/n4423 ;
  wire \u2_Display/n4424 ;
  wire \u2_Display/n4425 ;
  wire \u2_Display/n4426 ;
  wire \u2_Display/n4427 ;
  wire \u2_Display/n4428 ;
  wire \u2_Display/n4429 ;
  wire \u2_Display/n443 ;
  wire \u2_Display/n4430 ;
  wire \u2_Display/n4431 ;
  wire \u2_Display/n4432 ;
  wire \u2_Display/n4433 ;
  wire \u2_Display/n4434 ;
  wire \u2_Display/n4435 ;
  wire \u2_Display/n4436 ;
  wire \u2_Display/n4437 ;
  wire \u2_Display/n4438 ;
  wire \u2_Display/n4439 ;
  wire \u2_Display/n444 ;
  wire \u2_Display/n4440 ;
  wire \u2_Display/n4441 ;
  wire \u2_Display/n4442 ;
  wire \u2_Display/n4443 ;
  wire \u2_Display/n4444 ;
  wire \u2_Display/n4445 ;
  wire \u2_Display/n4446 ;
  wire \u2_Display/n4447 ;
  wire \u2_Display/n4448 ;
  wire \u2_Display/n4449 ;
  wire \u2_Display/n445 ;
  wire \u2_Display/n4450 ;
  wire \u2_Display/n4451 ;
  wire \u2_Display/n4452 ;
  wire \u2_Display/n4454 ;
  wire \u2_Display/n4455 ;
  wire \u2_Display/n4456 ;
  wire \u2_Display/n4457 ;
  wire \u2_Display/n4458 ;
  wire \u2_Display/n4459 ;
  wire \u2_Display/n446 ;
  wire \u2_Display/n4460 ;
  wire \u2_Display/n4461 ;
  wire \u2_Display/n4462 ;
  wire \u2_Display/n4463 ;
  wire \u2_Display/n4464 ;
  wire \u2_Display/n4465 ;
  wire \u2_Display/n4466 ;
  wire \u2_Display/n4467 ;
  wire \u2_Display/n4468 ;
  wire \u2_Display/n4469 ;
  wire \u2_Display/n447 ;
  wire \u2_Display/n4470 ;
  wire \u2_Display/n4471 ;
  wire \u2_Display/n4472 ;
  wire \u2_Display/n4473 ;
  wire \u2_Display/n4474 ;
  wire \u2_Display/n4475 ;
  wire \u2_Display/n4476 ;
  wire \u2_Display/n4477 ;
  wire \u2_Display/n4478 ;
  wire \u2_Display/n4479 ;
  wire \u2_Display/n448 ;
  wire \u2_Display/n4480 ;
  wire \u2_Display/n4481 ;
  wire \u2_Display/n4482 ;
  wire \u2_Display/n4483 ;
  wire \u2_Display/n4484 ;
  wire \u2_Display/n4485 ;
  wire \u2_Display/n4486 ;
  wire \u2_Display/n4487 ;
  wire \u2_Display/n4489 ;
  wire \u2_Display/n449 ;
  wire \u2_Display/n4490 ;
  wire \u2_Display/n4491 ;
  wire \u2_Display/n4492 ;
  wire \u2_Display/n4493 ;
  wire \u2_Display/n4494 ;
  wire \u2_Display/n4495 ;
  wire \u2_Display/n4496 ;
  wire \u2_Display/n4497 ;
  wire \u2_Display/n4498 ;
  wire \u2_Display/n4499 ;
  wire \u2_Display/n45 ;
  wire \u2_Display/n450 ;
  wire \u2_Display/n4500 ;
  wire \u2_Display/n4501 ;
  wire \u2_Display/n4502 ;
  wire \u2_Display/n4503 ;
  wire \u2_Display/n4504 ;
  wire \u2_Display/n4505 ;
  wire \u2_Display/n4506 ;
  wire \u2_Display/n4507 ;
  wire \u2_Display/n4508 ;
  wire \u2_Display/n4509 ;
  wire \u2_Display/n451 ;
  wire \u2_Display/n4510 ;
  wire \u2_Display/n4511 ;
  wire \u2_Display/n4512 ;
  wire \u2_Display/n4513 ;
  wire \u2_Display/n4514 ;
  wire \u2_Display/n4515 ;
  wire \u2_Display/n4516 ;
  wire \u2_Display/n4517 ;
  wire \u2_Display/n4518 ;
  wire \u2_Display/n4519 ;
  wire \u2_Display/n452 ;
  wire \u2_Display/n4520 ;
  wire \u2_Display/n4521 ;
  wire \u2_Display/n4522 ;
  wire \u2_Display/n4524 ;
  wire \u2_Display/n4525 ;
  wire \u2_Display/n4526 ;
  wire \u2_Display/n4527 ;
  wire \u2_Display/n4528 ;
  wire \u2_Display/n4529 ;
  wire \u2_Display/n453 ;
  wire \u2_Display/n4530 ;
  wire \u2_Display/n4531 ;
  wire \u2_Display/n4532 ;
  wire \u2_Display/n4533 ;
  wire \u2_Display/n4534 ;
  wire \u2_Display/n4535 ;
  wire \u2_Display/n4536 ;
  wire \u2_Display/n4537 ;
  wire \u2_Display/n4538 ;
  wire \u2_Display/n4539 ;
  wire \u2_Display/n4540 ;
  wire \u2_Display/n4541 ;
  wire \u2_Display/n4542 ;
  wire \u2_Display/n4543 ;
  wire \u2_Display/n4544 ;
  wire \u2_Display/n4545 ;
  wire \u2_Display/n4546 ;
  wire \u2_Display/n4547 ;
  wire \u2_Display/n4548 ;
  wire \u2_Display/n4549 ;
  wire \u2_Display/n455 ;
  wire \u2_Display/n4550 ;
  wire \u2_Display/n4551 ;
  wire \u2_Display/n4552 ;
  wire \u2_Display/n4553 ;
  wire \u2_Display/n4554 ;
  wire \u2_Display/n4555 ;
  wire \u2_Display/n4556 ;
  wire \u2_Display/n4557 ;
  wire \u2_Display/n456 ;
  wire \u2_Display/n457 ;
  wire \u2_Display/n458 ;
  wire \u2_Display/n459 ;
  wire \u2_Display/n46 ;
  wire \u2_Display/n460 ;
  wire \u2_Display/n461 ;
  wire \u2_Display/n462 ;
  wire \u2_Display/n463 ;
  wire \u2_Display/n464 ;
  wire \u2_Display/n465 ;
  wire \u2_Display/n466 ;
  wire \u2_Display/n467 ;
  wire \u2_Display/n468 ;
  wire \u2_Display/n469 ;
  wire \u2_Display/n470 ;
  wire \u2_Display/n471 ;
  wire \u2_Display/n472 ;
  wire \u2_Display/n473 ;
  wire \u2_Display/n474 ;
  wire \u2_Display/n475 ;
  wire \u2_Display/n476 ;
  wire \u2_Display/n477 ;
  wire \u2_Display/n478 ;
  wire \u2_Display/n479 ;
  wire \u2_Display/n48 ;
  wire \u2_Display/n480 ;
  wire \u2_Display/n481 ;
  wire \u2_Display/n482 ;
  wire \u2_Display/n483 ;
  wire \u2_Display/n484 ;
  wire \u2_Display/n485 ;
  wire \u2_Display/n486 ;
  wire \u2_Display/n487 ;
  wire \u2_Display/n488 ;
  wire \u2_Display/n49 ;
  wire \u2_Display/n490 ;
  wire \u2_Display/n4909 ;
  wire \u2_Display/n491 ;
  wire \u2_Display/n492 ;
  wire \u2_Display/n493 ;
  wire \u2_Display/n494 ;
  wire \u2_Display/n4944 ;
  wire \u2_Display/n495 ;
  wire \u2_Display/n496 ;
  wire \u2_Display/n497 ;
  wire \u2_Display/n4979 ;
  wire \u2_Display/n498 ;
  wire \u2_Display/n499 ;
  wire \u2_Display/n50 ;
  wire \u2_Display/n500 ;
  wire \u2_Display/n501 ;
  wire \u2_Display/n5014 ;
  wire \u2_Display/n502 ;
  wire \u2_Display/n503 ;
  wire \u2_Display/n504 ;
  wire \u2_Display/n5049 ;
  wire \u2_Display/n505 ;
  wire \u2_Display/n506 ;
  wire \u2_Display/n507 ;
  wire \u2_Display/n508 ;
  wire \u2_Display/n5084 ;
  wire \u2_Display/n509 ;
  wire \u2_Display/n51 ;
  wire \u2_Display/n510 ;
  wire \u2_Display/n511 ;
  wire \u2_Display/n5119 ;
  wire \u2_Display/n512 ;
  wire \u2_Display/n513 ;
  wire \u2_Display/n514 ;
  wire \u2_Display/n515 ;
  wire \u2_Display/n5154 ;
  wire \u2_Display/n516 ;
  wire \u2_Display/n517 ;
  wire \u2_Display/n518 ;
  wire \u2_Display/n5189 ;
  wire \u2_Display/n519 ;
  wire \u2_Display/n5196 ;
  wire \u2_Display/n5197 ;
  wire \u2_Display/n5198 ;
  wire \u2_Display/n5199 ;
  wire \u2_Display/n520 ;
  wire \u2_Display/n5200 ;
  wire \u2_Display/n5201 ;
  wire \u2_Display/n5202 ;
  wire \u2_Display/n5203 ;
  wire \u2_Display/n5204 ;
  wire \u2_Display/n5205 ;
  wire \u2_Display/n5206 ;
  wire \u2_Display/n5207 ;
  wire \u2_Display/n5208 ;
  wire \u2_Display/n5209 ;
  wire \u2_Display/n521 ;
  wire \u2_Display/n5210 ;
  wire \u2_Display/n5211 ;
  wire \u2_Display/n5212 ;
  wire \u2_Display/n5213 ;
  wire \u2_Display/n5214 ;
  wire \u2_Display/n5215 ;
  wire \u2_Display/n5216 ;
  wire \u2_Display/n5217 ;
  wire \u2_Display/n5218 ;
  wire \u2_Display/n5219 ;
  wire \u2_Display/n522 ;
  wire \u2_Display/n5220 ;
  wire \u2_Display/n5221 ;
  wire \u2_Display/n5222 ;
  wire \u2_Display/n5223 ;
  wire \u2_Display/n5224 ;
  wire \u2_Display/n5225 ;
  wire \u2_Display/n5227 ;
  wire \u2_Display/n5228 ;
  wire \u2_Display/n5229 ;
  wire \u2_Display/n523 ;
  wire \u2_Display/n5230 ;
  wire \u2_Display/n5231 ;
  wire \u2_Display/n5232 ;
  wire \u2_Display/n5233 ;
  wire \u2_Display/n5234 ;
  wire \u2_Display/n5235 ;
  wire \u2_Display/n5236 ;
  wire \u2_Display/n5237 ;
  wire \u2_Display/n5238 ;
  wire \u2_Display/n5239 ;
  wire \u2_Display/n5240 ;
  wire \u2_Display/n5241 ;
  wire \u2_Display/n5242 ;
  wire \u2_Display/n5243 ;
  wire \u2_Display/n5244 ;
  wire \u2_Display/n5245 ;
  wire \u2_Display/n5246 ;
  wire \u2_Display/n5247 ;
  wire \u2_Display/n5248 ;
  wire \u2_Display/n5249 ;
  wire \u2_Display/n525 ;
  wire \u2_Display/n5250 ;
  wire \u2_Display/n5251 ;
  wire \u2_Display/n5252 ;
  wire \u2_Display/n5253 ;
  wire \u2_Display/n5254 ;
  wire \u2_Display/n5255 ;
  wire \u2_Display/n5256 ;
  wire \u2_Display/n5257 ;
  wire \u2_Display/n5258 ;
  wire \u2_Display/n5259 ;
  wire \u2_Display/n526 ;
  wire \u2_Display/n5260 ;
  wire \u2_Display/n5262 ;
  wire \u2_Display/n5263 ;
  wire \u2_Display/n5264 ;
  wire \u2_Display/n5265 ;
  wire \u2_Display/n5266 ;
  wire \u2_Display/n5267 ;
  wire \u2_Display/n5268 ;
  wire \u2_Display/n5269 ;
  wire \u2_Display/n527 ;
  wire \u2_Display/n5270 ;
  wire \u2_Display/n5271 ;
  wire \u2_Display/n5272 ;
  wire \u2_Display/n5273 ;
  wire \u2_Display/n5274 ;
  wire \u2_Display/n5275 ;
  wire \u2_Display/n5276 ;
  wire \u2_Display/n5277 ;
  wire \u2_Display/n5278 ;
  wire \u2_Display/n5279 ;
  wire \u2_Display/n528 ;
  wire \u2_Display/n5280 ;
  wire \u2_Display/n5281 ;
  wire \u2_Display/n5282 ;
  wire \u2_Display/n5283 ;
  wire \u2_Display/n5284 ;
  wire \u2_Display/n5285 ;
  wire \u2_Display/n5286 ;
  wire \u2_Display/n5287 ;
  wire \u2_Display/n5288 ;
  wire \u2_Display/n5289 ;
  wire \u2_Display/n529 ;
  wire \u2_Display/n5290 ;
  wire \u2_Display/n5291 ;
  wire \u2_Display/n5292 ;
  wire \u2_Display/n5293 ;
  wire \u2_Display/n5294 ;
  wire \u2_Display/n5295 ;
  wire \u2_Display/n5297 ;
  wire \u2_Display/n5298 ;
  wire \u2_Display/n5299 ;
  wire \u2_Display/n530 ;
  wire \u2_Display/n5300 ;
  wire \u2_Display/n5301 ;
  wire \u2_Display/n5302 ;
  wire \u2_Display/n5303 ;
  wire \u2_Display/n5304 ;
  wire \u2_Display/n5305 ;
  wire \u2_Display/n5306 ;
  wire \u2_Display/n5307 ;
  wire \u2_Display/n5308 ;
  wire \u2_Display/n5309 ;
  wire \u2_Display/n531 ;
  wire \u2_Display/n5310 ;
  wire \u2_Display/n5311 ;
  wire \u2_Display/n5312 ;
  wire \u2_Display/n5313 ;
  wire \u2_Display/n5314 ;
  wire \u2_Display/n5315 ;
  wire \u2_Display/n5316 ;
  wire \u2_Display/n5317 ;
  wire \u2_Display/n5318 ;
  wire \u2_Display/n5319 ;
  wire \u2_Display/n532 ;
  wire \u2_Display/n5320 ;
  wire \u2_Display/n5321 ;
  wire \u2_Display/n5322 ;
  wire \u2_Display/n5323 ;
  wire \u2_Display/n5324 ;
  wire \u2_Display/n5325 ;
  wire \u2_Display/n5326 ;
  wire \u2_Display/n5327 ;
  wire \u2_Display/n5328 ;
  wire \u2_Display/n5329 ;
  wire \u2_Display/n533 ;
  wire \u2_Display/n5330 ;
  wire \u2_Display/n5332 ;
  wire \u2_Display/n5333 ;
  wire \u2_Display/n5334 ;
  wire \u2_Display/n5335 ;
  wire \u2_Display/n5336 ;
  wire \u2_Display/n5337 ;
  wire \u2_Display/n5338 ;
  wire \u2_Display/n5339 ;
  wire \u2_Display/n534 ;
  wire \u2_Display/n5340 ;
  wire \u2_Display/n5341 ;
  wire \u2_Display/n5342 ;
  wire \u2_Display/n5343 ;
  wire \u2_Display/n5344 ;
  wire \u2_Display/n5345 ;
  wire \u2_Display/n5346 ;
  wire \u2_Display/n5347 ;
  wire \u2_Display/n5348 ;
  wire \u2_Display/n5349 ;
  wire \u2_Display/n535 ;
  wire \u2_Display/n5350 ;
  wire \u2_Display/n5351 ;
  wire \u2_Display/n5352 ;
  wire \u2_Display/n5353 ;
  wire \u2_Display/n5354 ;
  wire \u2_Display/n5355 ;
  wire \u2_Display/n5356 ;
  wire \u2_Display/n5357 ;
  wire \u2_Display/n5358 ;
  wire \u2_Display/n5359 ;
  wire \u2_Display/n536 ;
  wire \u2_Display/n5360 ;
  wire \u2_Display/n5361 ;
  wire \u2_Display/n5362 ;
  wire \u2_Display/n5363 ;
  wire \u2_Display/n5364 ;
  wire \u2_Display/n5365 ;
  wire \u2_Display/n5367 ;
  wire \u2_Display/n5368 ;
  wire \u2_Display/n5369 ;
  wire \u2_Display/n537 ;
  wire \u2_Display/n5370 ;
  wire \u2_Display/n5371 ;
  wire \u2_Display/n5372 ;
  wire \u2_Display/n5373 ;
  wire \u2_Display/n5374 ;
  wire \u2_Display/n5375 ;
  wire \u2_Display/n5376 ;
  wire \u2_Display/n5377 ;
  wire \u2_Display/n5378 ;
  wire \u2_Display/n5379 ;
  wire \u2_Display/n538 ;
  wire \u2_Display/n5380 ;
  wire \u2_Display/n5381 ;
  wire \u2_Display/n5382 ;
  wire \u2_Display/n5383 ;
  wire \u2_Display/n5384 ;
  wire \u2_Display/n5385 ;
  wire \u2_Display/n5386 ;
  wire \u2_Display/n5387 ;
  wire \u2_Display/n5388 ;
  wire \u2_Display/n5389 ;
  wire \u2_Display/n539 ;
  wire \u2_Display/n5390 ;
  wire \u2_Display/n5391 ;
  wire \u2_Display/n5392 ;
  wire \u2_Display/n5393 ;
  wire \u2_Display/n5394 ;
  wire \u2_Display/n5395 ;
  wire \u2_Display/n5396 ;
  wire \u2_Display/n5397 ;
  wire \u2_Display/n5398 ;
  wire \u2_Display/n5399 ;
  wire \u2_Display/n540 ;
  wire \u2_Display/n5400 ;
  wire \u2_Display/n5402 ;
  wire \u2_Display/n5403 ;
  wire \u2_Display/n5404 ;
  wire \u2_Display/n5405 ;
  wire \u2_Display/n5406 ;
  wire \u2_Display/n5407 ;
  wire \u2_Display/n5408 ;
  wire \u2_Display/n5409 ;
  wire \u2_Display/n541 ;
  wire \u2_Display/n5410 ;
  wire \u2_Display/n5411 ;
  wire \u2_Display/n5412 ;
  wire \u2_Display/n5413 ;
  wire \u2_Display/n5414 ;
  wire \u2_Display/n5415 ;
  wire \u2_Display/n5416 ;
  wire \u2_Display/n5417 ;
  wire \u2_Display/n5418 ;
  wire \u2_Display/n5419 ;
  wire \u2_Display/n542 ;
  wire \u2_Display/n5420 ;
  wire \u2_Display/n5421 ;
  wire \u2_Display/n5422 ;
  wire \u2_Display/n5423 ;
  wire \u2_Display/n5424 ;
  wire \u2_Display/n5425 ;
  wire \u2_Display/n5426 ;
  wire \u2_Display/n5427 ;
  wire \u2_Display/n5428 ;
  wire \u2_Display/n5429 ;
  wire \u2_Display/n543 ;
  wire \u2_Display/n5430 ;
  wire \u2_Display/n5431 ;
  wire \u2_Display/n5432 ;
  wire \u2_Display/n5433 ;
  wire \u2_Display/n5434 ;
  wire \u2_Display/n5435 ;
  wire \u2_Display/n5437 ;
  wire \u2_Display/n5438 ;
  wire \u2_Display/n5439 ;
  wire \u2_Display/n544 ;
  wire \u2_Display/n5440 ;
  wire \u2_Display/n5441 ;
  wire \u2_Display/n5442 ;
  wire \u2_Display/n5443 ;
  wire \u2_Display/n5444 ;
  wire \u2_Display/n5445 ;
  wire \u2_Display/n5446 ;
  wire \u2_Display/n5447 ;
  wire \u2_Display/n5448 ;
  wire \u2_Display/n5449 ;
  wire \u2_Display/n545 ;
  wire \u2_Display/n5450 ;
  wire \u2_Display/n5451 ;
  wire \u2_Display/n5452 ;
  wire \u2_Display/n5453 ;
  wire \u2_Display/n5454 ;
  wire \u2_Display/n5455 ;
  wire \u2_Display/n5456 ;
  wire \u2_Display/n5457 ;
  wire \u2_Display/n5458 ;
  wire \u2_Display/n5459 ;
  wire \u2_Display/n546 ;
  wire \u2_Display/n5460 ;
  wire \u2_Display/n5461 ;
  wire \u2_Display/n5462 ;
  wire \u2_Display/n5463 ;
  wire \u2_Display/n5464 ;
  wire \u2_Display/n5465 ;
  wire \u2_Display/n5466 ;
  wire \u2_Display/n5467 ;
  wire \u2_Display/n5468 ;
  wire \u2_Display/n5469 ;
  wire \u2_Display/n547 ;
  wire \u2_Display/n5470 ;
  wire \u2_Display/n5472 ;
  wire \u2_Display/n5473 ;
  wire \u2_Display/n5474 ;
  wire \u2_Display/n5475 ;
  wire \u2_Display/n5476 ;
  wire \u2_Display/n5477 ;
  wire \u2_Display/n5478 ;
  wire \u2_Display/n5479 ;
  wire \u2_Display/n548 ;
  wire \u2_Display/n5480 ;
  wire \u2_Display/n5481 ;
  wire \u2_Display/n5482 ;
  wire \u2_Display/n5483 ;
  wire \u2_Display/n5484 ;
  wire \u2_Display/n5485 ;
  wire \u2_Display/n5486 ;
  wire \u2_Display/n5487 ;
  wire \u2_Display/n5488 ;
  wire \u2_Display/n5489 ;
  wire \u2_Display/n549 ;
  wire \u2_Display/n5490 ;
  wire \u2_Display/n5491 ;
  wire \u2_Display/n5492 ;
  wire \u2_Display/n5493 ;
  wire \u2_Display/n5494 ;
  wire \u2_Display/n5495 ;
  wire \u2_Display/n5496 ;
  wire \u2_Display/n5497 ;
  wire \u2_Display/n5498 ;
  wire \u2_Display/n5499 ;
  wire \u2_Display/n550 ;
  wire \u2_Display/n5500 ;
  wire \u2_Display/n5501 ;
  wire \u2_Display/n5502 ;
  wire \u2_Display/n5503 ;
  wire \u2_Display/n5504 ;
  wire \u2_Display/n5505 ;
  wire \u2_Display/n5507 ;
  wire \u2_Display/n5508 ;
  wire \u2_Display/n5509 ;
  wire \u2_Display/n551 ;
  wire \u2_Display/n5510 ;
  wire \u2_Display/n5511 ;
  wire \u2_Display/n5512 ;
  wire \u2_Display/n5513 ;
  wire \u2_Display/n5514 ;
  wire \u2_Display/n5515 ;
  wire \u2_Display/n5516 ;
  wire \u2_Display/n5517 ;
  wire \u2_Display/n5518 ;
  wire \u2_Display/n5519 ;
  wire \u2_Display/n552 ;
  wire \u2_Display/n5520 ;
  wire \u2_Display/n5521 ;
  wire \u2_Display/n5522 ;
  wire \u2_Display/n5523 ;
  wire \u2_Display/n5524 ;
  wire \u2_Display/n5525 ;
  wire \u2_Display/n5526 ;
  wire \u2_Display/n5527 ;
  wire \u2_Display/n5528 ;
  wire \u2_Display/n5529 ;
  wire \u2_Display/n553 ;
  wire \u2_Display/n5530 ;
  wire \u2_Display/n5531 ;
  wire \u2_Display/n5532 ;
  wire \u2_Display/n5533 ;
  wire \u2_Display/n5534 ;
  wire \u2_Display/n5535 ;
  wire \u2_Display/n5536 ;
  wire \u2_Display/n5537 ;
  wire \u2_Display/n5538 ;
  wire \u2_Display/n5539 ;
  wire \u2_Display/n554 ;
  wire \u2_Display/n5540 ;
  wire \u2_Display/n5542 ;
  wire \u2_Display/n5543 ;
  wire \u2_Display/n5544 ;
  wire \u2_Display/n5545 ;
  wire \u2_Display/n5546 ;
  wire \u2_Display/n5547 ;
  wire \u2_Display/n5548 ;
  wire \u2_Display/n5549 ;
  wire \u2_Display/n555 ;
  wire \u2_Display/n5550 ;
  wire \u2_Display/n5551 ;
  wire \u2_Display/n5552 ;
  wire \u2_Display/n5553 ;
  wire \u2_Display/n5554 ;
  wire \u2_Display/n5555 ;
  wire \u2_Display/n5556 ;
  wire \u2_Display/n5557 ;
  wire \u2_Display/n5558 ;
  wire \u2_Display/n5559 ;
  wire \u2_Display/n556 ;
  wire \u2_Display/n5560 ;
  wire \u2_Display/n5561 ;
  wire \u2_Display/n5562 ;
  wire \u2_Display/n5563 ;
  wire \u2_Display/n5564 ;
  wire \u2_Display/n5565 ;
  wire \u2_Display/n5566 ;
  wire \u2_Display/n5567 ;
  wire \u2_Display/n5568 ;
  wire \u2_Display/n5569 ;
  wire \u2_Display/n557 ;
  wire \u2_Display/n5570 ;
  wire \u2_Display/n5571 ;
  wire \u2_Display/n5572 ;
  wire \u2_Display/n5573 ;
  wire \u2_Display/n5574 ;
  wire \u2_Display/n5575 ;
  wire \u2_Display/n5577 ;
  wire \u2_Display/n5578 ;
  wire \u2_Display/n5579 ;
  wire \u2_Display/n558 ;
  wire \u2_Display/n5580 ;
  wire \u2_Display/n5581 ;
  wire \u2_Display/n5582 ;
  wire \u2_Display/n5583 ;
  wire \u2_Display/n5584 ;
  wire \u2_Display/n5585 ;
  wire \u2_Display/n5586 ;
  wire \u2_Display/n5587 ;
  wire \u2_Display/n5588 ;
  wire \u2_Display/n5589 ;
  wire \u2_Display/n5590 ;
  wire \u2_Display/n5591 ;
  wire \u2_Display/n5592 ;
  wire \u2_Display/n5593 ;
  wire \u2_Display/n5594 ;
  wire \u2_Display/n5595 ;
  wire \u2_Display/n5596 ;
  wire \u2_Display/n5597 ;
  wire \u2_Display/n5598 ;
  wire \u2_Display/n5599 ;
  wire \u2_Display/n560 ;
  wire \u2_Display/n5600 ;
  wire \u2_Display/n5601 ;
  wire \u2_Display/n5602 ;
  wire \u2_Display/n5603 ;
  wire \u2_Display/n5604 ;
  wire \u2_Display/n5605 ;
  wire \u2_Display/n5606 ;
  wire \u2_Display/n5607 ;
  wire \u2_Display/n5608 ;
  wire \u2_Display/n5609 ;
  wire \u2_Display/n561 ;
  wire \u2_Display/n5610 ;
  wire \u2_Display/n5612 ;
  wire \u2_Display/n5613 ;
  wire \u2_Display/n5614 ;
  wire \u2_Display/n5615 ;
  wire \u2_Display/n5616 ;
  wire \u2_Display/n5617 ;
  wire \u2_Display/n5618 ;
  wire \u2_Display/n5619 ;
  wire \u2_Display/n562 ;
  wire \u2_Display/n5620 ;
  wire \u2_Display/n5621 ;
  wire \u2_Display/n5622 ;
  wire \u2_Display/n5623 ;
  wire \u2_Display/n5624 ;
  wire \u2_Display/n5625 ;
  wire \u2_Display/n5626 ;
  wire \u2_Display/n5627 ;
  wire \u2_Display/n5628 ;
  wire \u2_Display/n5629 ;
  wire \u2_Display/n563 ;
  wire \u2_Display/n5630 ;
  wire \u2_Display/n5631 ;
  wire \u2_Display/n5632 ;
  wire \u2_Display/n5633 ;
  wire \u2_Display/n5634 ;
  wire \u2_Display/n5635 ;
  wire \u2_Display/n5636 ;
  wire \u2_Display/n5637 ;
  wire \u2_Display/n5638 ;
  wire \u2_Display/n5639 ;
  wire \u2_Display/n564 ;
  wire \u2_Display/n5640 ;
  wire \u2_Display/n5641 ;
  wire \u2_Display/n5642 ;
  wire \u2_Display/n5643 ;
  wire \u2_Display/n5644 ;
  wire \u2_Display/n5645 ;
  wire \u2_Display/n5647 ;
  wire \u2_Display/n5648 ;
  wire \u2_Display/n5649 ;
  wire \u2_Display/n565 ;
  wire \u2_Display/n5650 ;
  wire \u2_Display/n5651 ;
  wire \u2_Display/n5652 ;
  wire \u2_Display/n5653 ;
  wire \u2_Display/n5654 ;
  wire \u2_Display/n5655 ;
  wire \u2_Display/n5656 ;
  wire \u2_Display/n5657 ;
  wire \u2_Display/n5658 ;
  wire \u2_Display/n5659 ;
  wire \u2_Display/n566 ;
  wire \u2_Display/n5660 ;
  wire \u2_Display/n5661 ;
  wire \u2_Display/n5662 ;
  wire \u2_Display/n5663 ;
  wire \u2_Display/n5664 ;
  wire \u2_Display/n5665 ;
  wire \u2_Display/n5666 ;
  wire \u2_Display/n5667 ;
  wire \u2_Display/n5668 ;
  wire \u2_Display/n5669 ;
  wire \u2_Display/n567 ;
  wire \u2_Display/n5670 ;
  wire \u2_Display/n5671 ;
  wire \u2_Display/n5672 ;
  wire \u2_Display/n5673 ;
  wire \u2_Display/n5674 ;
  wire \u2_Display/n5675 ;
  wire \u2_Display/n5676 ;
  wire \u2_Display/n5677 ;
  wire \u2_Display/n5678 ;
  wire \u2_Display/n5679 ;
  wire \u2_Display/n568 ;
  wire \u2_Display/n5680 ;
  wire \u2_Display/n569 ;
  wire \u2_Display/n570 ;
  wire \u2_Display/n571 ;
  wire \u2_Display/n572 ;
  wire \u2_Display/n573 ;
  wire \u2_Display/n574 ;
  wire \u2_Display/n575 ;
  wire \u2_Display/n576 ;
  wire \u2_Display/n577 ;
  wire \u2_Display/n578 ;
  wire \u2_Display/n579 ;
  wire \u2_Display/n580 ;
  wire \u2_Display/n581 ;
  wire \u2_Display/n582 ;
  wire \u2_Display/n583 ;
  wire \u2_Display/n584 ;
  wire \u2_Display/n585 ;
  wire \u2_Display/n586 ;
  wire \u2_Display/n587 ;
  wire \u2_Display/n588 ;
  wire \u2_Display/n589 ;
  wire \u2_Display/n590 ;
  wire \u2_Display/n591 ;
  wire \u2_Display/n592 ;
  wire \u2_Display/n593 ;
  wire \u2_Display/n595 ;
  wire \u2_Display/n596 ;
  wire \u2_Display/n597 ;
  wire \u2_Display/n598 ;
  wire \u2_Display/n599 ;
  wire \u2_Display/n600 ;
  wire \u2_Display/n601 ;
  wire \u2_Display/n602 ;
  wire \u2_Display/n603 ;
  wire \u2_Display/n604 ;
  wire \u2_Display/n605 ;
  wire \u2_Display/n606 ;
  wire \u2_Display/n6068 ;
  wire \u2_Display/n607 ;
  wire \u2_Display/n6070 ;
  wire \u2_Display/n6071 ;
  wire \u2_Display/n6072 ;
  wire \u2_Display/n6073 ;
  wire \u2_Display/n6074 ;
  wire \u2_Display/n6075 ;
  wire \u2_Display/n6076 ;
  wire \u2_Display/n6077 ;
  wire \u2_Display/n6078 ;
  wire \u2_Display/n6079 ;
  wire \u2_Display/n608 ;
  wire \u2_Display/n6080 ;
  wire \u2_Display/n6081 ;
  wire \u2_Display/n6082 ;
  wire \u2_Display/n6083 ;
  wire \u2_Display/n6084 ;
  wire \u2_Display/n6085 ;
  wire \u2_Display/n6086 ;
  wire \u2_Display/n6087 ;
  wire \u2_Display/n6088 ;
  wire \u2_Display/n6089 ;
  wire \u2_Display/n609 ;
  wire \u2_Display/n6090 ;
  wire \u2_Display/n6091 ;
  wire \u2_Display/n6092 ;
  wire \u2_Display/n6093 ;
  wire \u2_Display/n6094 ;
  wire \u2_Display/n6095 ;
  wire \u2_Display/n6096 ;
  wire \u2_Display/n6097 ;
  wire \u2_Display/n6098 ;
  wire \u2_Display/n6099 ;
  wire \u2_Display/n610 ;
  wire \u2_Display/n6100 ;
  wire \u2_Display/n6101 ;
  wire \u2_Display/n6103 ;
  wire \u2_Display/n6105 ;
  wire \u2_Display/n6106 ;
  wire \u2_Display/n6107 ;
  wire \u2_Display/n6108 ;
  wire \u2_Display/n6109 ;
  wire \u2_Display/n611 ;
  wire \u2_Display/n6110 ;
  wire \u2_Display/n6111 ;
  wire \u2_Display/n6112 ;
  wire \u2_Display/n6113 ;
  wire \u2_Display/n6114 ;
  wire \u2_Display/n6115 ;
  wire \u2_Display/n6116 ;
  wire \u2_Display/n6117 ;
  wire \u2_Display/n6118 ;
  wire \u2_Display/n6119 ;
  wire \u2_Display/n612 ;
  wire \u2_Display/n6120 ;
  wire \u2_Display/n6121 ;
  wire \u2_Display/n6122 ;
  wire \u2_Display/n6123 ;
  wire \u2_Display/n6124 ;
  wire \u2_Display/n6125 ;
  wire \u2_Display/n6126 ;
  wire \u2_Display/n6127 ;
  wire \u2_Display/n6128 ;
  wire \u2_Display/n6129 ;
  wire \u2_Display/n613 ;
  wire \u2_Display/n6130 ;
  wire \u2_Display/n6131 ;
  wire \u2_Display/n6132 ;
  wire \u2_Display/n6133 ;
  wire \u2_Display/n6134 ;
  wire \u2_Display/n6135 ;
  wire \u2_Display/n6136 ;
  wire \u2_Display/n6138 ;
  wire \u2_Display/n614 ;
  wire \u2_Display/n6140 ;
  wire \u2_Display/n6141 ;
  wire \u2_Display/n6142 ;
  wire \u2_Display/n6143 ;
  wire \u2_Display/n6144 ;
  wire \u2_Display/n6145 ;
  wire \u2_Display/n6146 ;
  wire \u2_Display/n6147 ;
  wire \u2_Display/n6148 ;
  wire \u2_Display/n6149 ;
  wire \u2_Display/n615 ;
  wire \u2_Display/n6150 ;
  wire \u2_Display/n6151 ;
  wire \u2_Display/n6152 ;
  wire \u2_Display/n6153 ;
  wire \u2_Display/n6154 ;
  wire \u2_Display/n6155 ;
  wire \u2_Display/n6156 ;
  wire \u2_Display/n6157 ;
  wire \u2_Display/n6158 ;
  wire \u2_Display/n6159 ;
  wire \u2_Display/n616 ;
  wire \u2_Display/n6160 ;
  wire \u2_Display/n6161 ;
  wire \u2_Display/n6162 ;
  wire \u2_Display/n6163 ;
  wire \u2_Display/n6164 ;
  wire \u2_Display/n6165 ;
  wire \u2_Display/n6166 ;
  wire \u2_Display/n6167 ;
  wire \u2_Display/n6168 ;
  wire \u2_Display/n6169 ;
  wire \u2_Display/n617 ;
  wire \u2_Display/n6170 ;
  wire \u2_Display/n6171 ;
  wire \u2_Display/n6173 ;
  wire \u2_Display/n6175 ;
  wire \u2_Display/n6176 ;
  wire \u2_Display/n6177 ;
  wire \u2_Display/n6178 ;
  wire \u2_Display/n6179 ;
  wire \u2_Display/n618 ;
  wire \u2_Display/n6180 ;
  wire \u2_Display/n6181 ;
  wire \u2_Display/n6182 ;
  wire \u2_Display/n6183 ;
  wire \u2_Display/n6184 ;
  wire \u2_Display/n6185 ;
  wire \u2_Display/n6186 ;
  wire \u2_Display/n6187 ;
  wire \u2_Display/n6188 ;
  wire \u2_Display/n6189 ;
  wire \u2_Display/n619 ;
  wire \u2_Display/n6190 ;
  wire \u2_Display/n6191 ;
  wire \u2_Display/n6192 ;
  wire \u2_Display/n6193 ;
  wire \u2_Display/n6194 ;
  wire \u2_Display/n6195 ;
  wire \u2_Display/n6196 ;
  wire \u2_Display/n6197 ;
  wire \u2_Display/n6198 ;
  wire \u2_Display/n6199 ;
  wire \u2_Display/n620 ;
  wire \u2_Display/n6200 ;
  wire \u2_Display/n6201 ;
  wire \u2_Display/n6202 ;
  wire \u2_Display/n6203 ;
  wire \u2_Display/n6204 ;
  wire \u2_Display/n6205 ;
  wire \u2_Display/n6206 ;
  wire \u2_Display/n6208 ;
  wire \u2_Display/n621 ;
  wire \u2_Display/n6210 ;
  wire \u2_Display/n6211 ;
  wire \u2_Display/n6212 ;
  wire \u2_Display/n6213 ;
  wire \u2_Display/n6214 ;
  wire \u2_Display/n6215 ;
  wire \u2_Display/n6216 ;
  wire \u2_Display/n6217 ;
  wire \u2_Display/n6218 ;
  wire \u2_Display/n6219 ;
  wire \u2_Display/n622 ;
  wire \u2_Display/n6220 ;
  wire \u2_Display/n6221 ;
  wire \u2_Display/n6222 ;
  wire \u2_Display/n6223 ;
  wire \u2_Display/n6224 ;
  wire \u2_Display/n6225 ;
  wire \u2_Display/n6226 ;
  wire \u2_Display/n6227 ;
  wire \u2_Display/n6228 ;
  wire \u2_Display/n6229 ;
  wire \u2_Display/n623 ;
  wire \u2_Display/n6230 ;
  wire \u2_Display/n6231 ;
  wire \u2_Display/n6232 ;
  wire \u2_Display/n6233 ;
  wire \u2_Display/n6234 ;
  wire \u2_Display/n6235 ;
  wire \u2_Display/n6236 ;
  wire \u2_Display/n6237 ;
  wire \u2_Display/n6238 ;
  wire \u2_Display/n6239 ;
  wire \u2_Display/n624 ;
  wire \u2_Display/n6240 ;
  wire \u2_Display/n6241 ;
  wire \u2_Display/n6243 ;
  wire \u2_Display/n6245 ;
  wire \u2_Display/n6246 ;
  wire \u2_Display/n6247 ;
  wire \u2_Display/n6248 ;
  wire \u2_Display/n6249 ;
  wire \u2_Display/n625 ;
  wire \u2_Display/n6250 ;
  wire \u2_Display/n6251 ;
  wire \u2_Display/n6252 ;
  wire \u2_Display/n6253 ;
  wire \u2_Display/n6254 ;
  wire \u2_Display/n6255 ;
  wire \u2_Display/n6256 ;
  wire \u2_Display/n6257 ;
  wire \u2_Display/n6258 ;
  wire \u2_Display/n6259 ;
  wire \u2_Display/n626 ;
  wire \u2_Display/n6260 ;
  wire \u2_Display/n6261 ;
  wire \u2_Display/n6262 ;
  wire \u2_Display/n6263 ;
  wire \u2_Display/n6264 ;
  wire \u2_Display/n6265 ;
  wire \u2_Display/n6266 ;
  wire \u2_Display/n6267 ;
  wire \u2_Display/n6268 ;
  wire \u2_Display/n6269 ;
  wire \u2_Display/n627 ;
  wire \u2_Display/n6270 ;
  wire \u2_Display/n6271 ;
  wire \u2_Display/n6272 ;
  wire \u2_Display/n6273 ;
  wire \u2_Display/n6274 ;
  wire \u2_Display/n6275 ;
  wire \u2_Display/n6276 ;
  wire \u2_Display/n6278 ;
  wire \u2_Display/n628 ;
  wire \u2_Display/n6280 ;
  wire \u2_Display/n6281 ;
  wire \u2_Display/n6282 ;
  wire \u2_Display/n6283 ;
  wire \u2_Display/n6284 ;
  wire \u2_Display/n6285 ;
  wire \u2_Display/n6286 ;
  wire \u2_Display/n6287 ;
  wire \u2_Display/n6288 ;
  wire \u2_Display/n6289 ;
  wire \u2_Display/n6290 ;
  wire \u2_Display/n6291 ;
  wire \u2_Display/n6292 ;
  wire \u2_Display/n6293 ;
  wire \u2_Display/n6294 ;
  wire \u2_Display/n6295 ;
  wire \u2_Display/n6296 ;
  wire \u2_Display/n6297 ;
  wire \u2_Display/n6298 ;
  wire \u2_Display/n6299 ;
  wire \u2_Display/n630 ;
  wire \u2_Display/n6300 ;
  wire \u2_Display/n6301 ;
  wire \u2_Display/n6302 ;
  wire \u2_Display/n6303 ;
  wire \u2_Display/n6304 ;
  wire \u2_Display/n6305 ;
  wire \u2_Display/n6306 ;
  wire \u2_Display/n6307 ;
  wire \u2_Display/n6308 ;
  wire \u2_Display/n6309 ;
  wire \u2_Display/n631 ;
  wire \u2_Display/n6310 ;
  wire \u2_Display/n6311 ;
  wire \u2_Display/n6313 ;
  wire \u2_Display/n6315 ;
  wire \u2_Display/n6316 ;
  wire \u2_Display/n6317 ;
  wire \u2_Display/n6318 ;
  wire \u2_Display/n6319 ;
  wire \u2_Display/n632 ;
  wire \u2_Display/n6320 ;
  wire \u2_Display/n6321 ;
  wire \u2_Display/n6322 ;
  wire \u2_Display/n6323 ;
  wire \u2_Display/n6324 ;
  wire \u2_Display/n6325 ;
  wire \u2_Display/n6326 ;
  wire \u2_Display/n6327 ;
  wire \u2_Display/n6328 ;
  wire \u2_Display/n6329 ;
  wire \u2_Display/n633 ;
  wire \u2_Display/n6330 ;
  wire \u2_Display/n6331 ;
  wire \u2_Display/n6332 ;
  wire \u2_Display/n6333 ;
  wire \u2_Display/n6334 ;
  wire \u2_Display/n6335 ;
  wire \u2_Display/n6336 ;
  wire \u2_Display/n6337 ;
  wire \u2_Display/n6338 ;
  wire \u2_Display/n6339 ;
  wire \u2_Display/n634 ;
  wire \u2_Display/n6340 ;
  wire \u2_Display/n6341 ;
  wire \u2_Display/n6342 ;
  wire \u2_Display/n6343 ;
  wire \u2_Display/n6344 ;
  wire \u2_Display/n6345 ;
  wire \u2_Display/n6346 ;
  wire \u2_Display/n6348 ;
  wire \u2_Display/n635 ;
  wire \u2_Display/n6350 ;
  wire \u2_Display/n6351 ;
  wire \u2_Display/n6352 ;
  wire \u2_Display/n6353 ;
  wire \u2_Display/n636 ;
  wire \u2_Display/n637 ;
  wire \u2_Display/n638 ;
  wire \u2_Display/n639 ;
  wire \u2_Display/n640 ;
  wire \u2_Display/n641 ;
  wire \u2_Display/n642 ;
  wire \u2_Display/n643 ;
  wire \u2_Display/n644 ;
  wire \u2_Display/n645 ;
  wire \u2_Display/n646 ;
  wire \u2_Display/n647 ;
  wire \u2_Display/n648 ;
  wire \u2_Display/n649 ;
  wire \u2_Display/n650 ;
  wire \u2_Display/n651 ;
  wire \u2_Display/n652 ;
  wire \u2_Display/n653 ;
  wire \u2_Display/n654 ;
  wire \u2_Display/n655 ;
  wire \u2_Display/n656 ;
  wire \u2_Display/n657 ;
  wire \u2_Display/n658 ;
  wire \u2_Display/n659 ;
  wire \u2_Display/n660 ;
  wire \u2_Display/n661 ;
  wire \u2_Display/n662 ;
  wire \u2_Display/n663 ;
  wire \u2_Display/n665 ;
  wire \u2_Display/n666 ;
  wire \u2_Display/n667 ;
  wire \u2_Display/n668 ;
  wire \u2_Display/n669 ;
  wire \u2_Display/n670 ;
  wire \u2_Display/n671 ;
  wire \u2_Display/n672 ;
  wire \u2_Display/n673 ;
  wire \u2_Display/n674 ;
  wire \u2_Display/n675 ;
  wire \u2_Display/n676 ;
  wire \u2_Display/n677 ;
  wire \u2_Display/n678 ;
  wire \u2_Display/n679 ;
  wire \u2_Display/n680 ;
  wire \u2_Display/n681 ;
  wire \u2_Display/n682 ;
  wire \u2_Display/n683 ;
  wire \u2_Display/n684 ;
  wire \u2_Display/n685 ;
  wire \u2_Display/n686 ;
  wire \u2_Display/n687 ;
  wire \u2_Display/n688 ;
  wire \u2_Display/n689 ;
  wire \u2_Display/n690 ;
  wire \u2_Display/n691 ;
  wire \u2_Display/n692 ;
  wire \u2_Display/n693 ;
  wire \u2_Display/n694 ;
  wire \u2_Display/n695 ;
  wire \u2_Display/n696 ;
  wire \u2_Display/n697 ;
  wire \u2_Display/n698 ;
  wire \u2_Display/n700 ;
  wire \u2_Display/n701 ;
  wire \u2_Display/n702 ;
  wire \u2_Display/n703 ;
  wire \u2_Display/n704 ;
  wire \u2_Display/n705 ;
  wire \u2_Display/n706 ;
  wire \u2_Display/n707 ;
  wire \u2_Display/n708 ;
  wire \u2_Display/n709 ;
  wire \u2_Display/n710 ;
  wire \u2_Display/n711 ;
  wire \u2_Display/n712 ;
  wire \u2_Display/n713 ;
  wire \u2_Display/n714 ;
  wire \u2_Display/n715 ;
  wire \u2_Display/n716 ;
  wire \u2_Display/n717 ;
  wire \u2_Display/n718 ;
  wire \u2_Display/n719 ;
  wire \u2_Display/n720 ;
  wire \u2_Display/n721 ;
  wire \u2_Display/n722 ;
  wire \u2_Display/n723 ;
  wire \u2_Display/n724 ;
  wire \u2_Display/n725 ;
  wire \u2_Display/n726 ;
  wire \u2_Display/n727 ;
  wire \u2_Display/n728 ;
  wire \u2_Display/n729 ;
  wire \u2_Display/n730 ;
  wire \u2_Display/n731 ;
  wire \u2_Display/n732 ;
  wire \u2_Display/n733 ;
  wire \u2_Display/n735 ;
  wire \u2_Display/n736 ;
  wire \u2_Display/n737 ;
  wire \u2_Display/n738 ;
  wire \u2_Display/n739 ;
  wire \u2_Display/n740 ;
  wire \u2_Display/n741 ;
  wire \u2_Display/n742 ;
  wire \u2_Display/n743 ;
  wire \u2_Display/n744 ;
  wire \u2_Display/n745 ;
  wire \u2_Display/n746 ;
  wire \u2_Display/n747 ;
  wire \u2_Display/n748 ;
  wire \u2_Display/n749 ;
  wire \u2_Display/n750 ;
  wire \u2_Display/n751 ;
  wire \u2_Display/n752 ;
  wire \u2_Display/n753 ;
  wire \u2_Display/n754 ;
  wire \u2_Display/n755 ;
  wire \u2_Display/n756 ;
  wire \u2_Display/n757 ;
  wire \u2_Display/n758 ;
  wire \u2_Display/n759 ;
  wire \u2_Display/n760 ;
  wire \u2_Display/n761 ;
  wire \u2_Display/n762 ;
  wire \u2_Display/n763 ;
  wire \u2_Display/n764 ;
  wire \u2_Display/n765 ;
  wire \u2_Display/n766 ;
  wire \u2_Display/n767 ;
  wire \u2_Display/n768 ;
  wire \u2_Display/n770 ;
  wire \u2_Display/n771 ;
  wire \u2_Display/n772 ;
  wire \u2_Display/n773 ;
  wire \u2_Display/n774 ;
  wire \u2_Display/n775 ;
  wire \u2_Display/n776 ;
  wire \u2_Display/n777 ;
  wire \u2_Display/n778 ;
  wire \u2_Display/n779 ;
  wire \u2_Display/n780 ;
  wire \u2_Display/n781 ;
  wire \u2_Display/n782 ;
  wire \u2_Display/n783 ;
  wire \u2_Display/n784 ;
  wire \u2_Display/n785 ;
  wire \u2_Display/n786 ;
  wire \u2_Display/n787 ;
  wire \u2_Display/n788 ;
  wire \u2_Display/n789 ;
  wire \u2_Display/n790 ;
  wire \u2_Display/n791 ;
  wire \u2_Display/n792 ;
  wire \u2_Display/n793 ;
  wire \u2_Display/n794 ;
  wire \u2_Display/n795 ;
  wire \u2_Display/n796 ;
  wire \u2_Display/n797 ;
  wire \u2_Display/n798 ;
  wire \u2_Display/n799 ;
  wire \u2_Display/n800 ;
  wire \u2_Display/n801 ;
  wire \u2_Display/n802 ;
  wire \u2_Display/n803 ;
  wire \u2_Display/n805 ;
  wire \u2_Display/n806 ;
  wire \u2_Display/n807 ;
  wire \u2_Display/n808 ;
  wire \u2_Display/n809 ;
  wire \u2_Display/n810 ;
  wire \u2_Display/n811 ;
  wire \u2_Display/n812 ;
  wire \u2_Display/n813 ;
  wire \u2_Display/n814 ;
  wire \u2_Display/n815 ;
  wire \u2_Display/n816 ;
  wire \u2_Display/n817 ;
  wire \u2_Display/n818 ;
  wire \u2_Display/n819 ;
  wire \u2_Display/n820 ;
  wire \u2_Display/n821 ;
  wire \u2_Display/n822 ;
  wire \u2_Display/n823 ;
  wire \u2_Display/n824 ;
  wire \u2_Display/n825 ;
  wire \u2_Display/n826 ;
  wire \u2_Display/n827 ;
  wire \u2_Display/n828 ;
  wire \u2_Display/n829 ;
  wire \u2_Display/n830 ;
  wire \u2_Display/n831 ;
  wire \u2_Display/n832 ;
  wire \u2_Display/n833 ;
  wire \u2_Display/n834 ;
  wire \u2_Display/n835 ;
  wire \u2_Display/n836 ;
  wire \u2_Display/n837 ;
  wire \u2_Display/n838 ;
  wire \u2_Display/n840 ;
  wire \u2_Display/n841 ;
  wire \u2_Display/n842 ;
  wire \u2_Display/n843 ;
  wire \u2_Display/n844 ;
  wire \u2_Display/n845 ;
  wire \u2_Display/n846 ;
  wire \u2_Display/n847 ;
  wire \u2_Display/n848 ;
  wire \u2_Display/n849 ;
  wire \u2_Display/n850 ;
  wire \u2_Display/n851 ;
  wire \u2_Display/n852 ;
  wire \u2_Display/n853 ;
  wire \u2_Display/n854 ;
  wire \u2_Display/n855 ;
  wire \u2_Display/n856 ;
  wire \u2_Display/n857 ;
  wire \u2_Display/n858 ;
  wire \u2_Display/n859 ;
  wire \u2_Display/n860 ;
  wire \u2_Display/n861 ;
  wire \u2_Display/n862 ;
  wire \u2_Display/n863 ;
  wire \u2_Display/n864 ;
  wire \u2_Display/n865 ;
  wire \u2_Display/n866 ;
  wire \u2_Display/n867 ;
  wire \u2_Display/n868 ;
  wire \u2_Display/n869 ;
  wire \u2_Display/n870 ;
  wire \u2_Display/n871 ;
  wire \u2_Display/n872 ;
  wire \u2_Display/n873 ;
  wire \u2_Display/n875 ;
  wire \u2_Display/n876 ;
  wire \u2_Display/n877 ;
  wire \u2_Display/n878 ;
  wire \u2_Display/n879 ;
  wire \u2_Display/n880 ;
  wire \u2_Display/n881 ;
  wire \u2_Display/n882 ;
  wire \u2_Display/n883 ;
  wire \u2_Display/n884 ;
  wire \u2_Display/n885 ;
  wire \u2_Display/n886 ;
  wire \u2_Display/n887 ;
  wire \u2_Display/n888 ;
  wire \u2_Display/n889 ;
  wire \u2_Display/n890 ;
  wire \u2_Display/n891 ;
  wire \u2_Display/n892 ;
  wire \u2_Display/n893 ;
  wire \u2_Display/n894 ;
  wire \u2_Display/n895 ;
  wire \u2_Display/n896 ;
  wire \u2_Display/n897 ;
  wire \u2_Display/n898 ;
  wire \u2_Display/n899 ;
  wire \u2_Display/n900 ;
  wire \u2_Display/n901 ;
  wire \u2_Display/n902 ;
  wire \u2_Display/n903 ;
  wire \u2_Display/n904 ;
  wire \u2_Display/n905 ;
  wire \u2_Display/n906 ;
  wire \u2_Display/n907 ;
  wire \u2_Display/n908 ;
  wire \u2_Display/n910 ;
  wire \u2_Display/n911 ;
  wire \u2_Display/n912 ;
  wire \u2_Display/n913 ;
  wire \u2_Display/n914 ;
  wire \u2_Display/n915 ;
  wire \u2_Display/n916 ;
  wire \u2_Display/n917 ;
  wire \u2_Display/n918 ;
  wire \u2_Display/n919 ;
  wire \u2_Display/n920 ;
  wire \u2_Display/n921 ;
  wire \u2_Display/n922 ;
  wire \u2_Display/n923 ;
  wire \u2_Display/n924 ;
  wire \u2_Display/n925 ;
  wire \u2_Display/n926 ;
  wire \u2_Display/n927 ;
  wire \u2_Display/n928 ;
  wire \u2_Display/n929 ;
  wire \u2_Display/n930 ;
  wire \u2_Display/n931 ;
  wire \u2_Display/n932 ;
  wire \u2_Display/n933 ;
  wire \u2_Display/n934 ;
  wire \u2_Display/n935 ;
  wire \u2_Display/n936 ;
  wire \u2_Display/n937 ;
  wire \u2_Display/n938 ;
  wire \u2_Display/n939 ;
  wire \u2_Display/n940 ;
  wire \u2_Display/n941 ;
  wire \u2_Display/n942 ;
  wire \u2_Display/n943 ;
  wire \u2_Display/n945 ;
  wire \u2_Display/n946 ;
  wire \u2_Display/n947 ;
  wire \u2_Display/n948 ;
  wire \u2_Display/n949 ;
  wire \u2_Display/n95 ;
  wire \u2_Display/n950 ;
  wire \u2_Display/n951 ;
  wire \u2_Display/n952 ;
  wire \u2_Display/n953 ;
  wire \u2_Display/n954 ;
  wire \u2_Display/n955 ;
  wire \u2_Display/n956 ;
  wire \u2_Display/n957 ;
  wire \u2_Display/n958 ;
  wire \u2_Display/n959 ;
  wire \u2_Display/n960 ;
  wire \u2_Display/n961 ;
  wire \u2_Display/n962 ;
  wire \u2_Display/n963 ;
  wire \u2_Display/n964 ;
  wire \u2_Display/n965 ;
  wire \u2_Display/n966 ;
  wire \u2_Display/n967 ;
  wire \u2_Display/n968 ;
  wire \u2_Display/n969 ;
  wire \u2_Display/n97 ;
  wire \u2_Display/n970 ;
  wire \u2_Display/n971 ;
  wire \u2_Display/n972 ;
  wire \u2_Display/n973 ;
  wire \u2_Display/n974 ;
  wire \u2_Display/n975 ;
  wire \u2_Display/n976 ;
  wire \u2_Display/n977 ;
  wire \u2_Display/n978 ;
  wire \u2_Display/n98 ;
  wire \u2_Display/n980 ;
  wire \u2_Display/n981 ;
  wire \u2_Display/n982 ;
  wire \u2_Display/n983 ;
  wire \u2_Display/n984 ;
  wire \u2_Display/n985 ;
  wire \u2_Display/n986 ;
  wire \u2_Display/n987 ;
  wire \u2_Display/n988 ;
  wire \u2_Display/n989 ;
  wire \u2_Display/n990 ;
  wire \u2_Display/n991 ;
  wire \u2_Display/n992 ;
  wire \u2_Display/n993 ;
  wire \u2_Display/n994 ;
  wire \u2_Display/n995 ;
  wire \u2_Display/n996 ;
  wire \u2_Display/n997 ;
  wire \u2_Display/n998 ;
  wire \u2_Display/n999 ;

  assign vga_b[7] = vga_b[0];
  assign vga_b[6] = vga_b[0];
  assign vga_b[5] = vga_b[0];
  assign vga_b[4] = vga_b[0];
  assign vga_b[3] = vga_b[0];
  assign vga_b[2] = vga_b[0];
  assign vga_b[1] = vga_b[0];
  assign vga_g[7] = vga_b[0];
  assign vga_g[6] = vga_b[0];
  assign vga_g[5] = vga_b[0];
  assign vga_g[4] = vga_b[0];
  assign vga_g[3] = vga_b[0];
  assign vga_g[2] = vga_b[0];
  assign vga_g[1] = vga_b[0];
  assign vga_g[0] = vga_b[0];
  assign vga_r[7] = vga_b[0];
  assign vga_r[6] = vga_b[0];
  assign vga_r[5] = vga_b[0];
  assign vga_r[4] = vga_b[0];
  assign vga_r[3] = vga_b[0];
  assign vga_r[2] = vga_b[0];
  assign vga_r[1] = vga_b[0];
  assign vga_r[0] = vga_b[0];
  not \on_off[0]_inv  (\on_off[0]_neg , on_off[0]);
  not \on_off[1]_inv  (\on_off[1]_neg , on_off[1]);
  not \on_off[2]_inv  (\on_off[2]_neg , on_off[2]);
  not \on_off[3]_inv  (\on_off[3]_neg , on_off[3]);
  not \on_off[4]_inv  (\on_off[4]_neg , on_off[4]);
  not \u0_PLL/u0  (\u0_PLL/n0 , rst_n);  // source/rtl/Clk_div.v(15)
  EG_LOGIC_BUFG \u0_PLL/uut/bufg_feedback  (
    .i(\u0_PLL/uut/clk0_buf ),
    .o(clk_vga));  // al_ip/PLL.v(34)
  EG_PHY_PLL #(
    .CLKC0_CPHASE(8),
    .CLKC0_DIV(9),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(1),
    .CLKC1_DIV(1),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_ENABLE("DISABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(1),
    .CLKC2_DIV(1),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("DISABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(1),
    .CLKC3_DIV(1),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("DISABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(9),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("24.000"),
    .FREQ_LOCK_ACCURACY(2),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .REFCLK_DIV(2),
    .REFCLK_SEL("INTERNAL"),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \u0_PLL/uut/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dwe(1'b0),
    .fbclk(clk_vga),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(clk_24m),
    .reset(\u0_PLL/n0 ),
    .stdby(1'b0),
    .clkc({open_n1,open_n2,open_n3,open_n4,\u0_PLL/uut/clk0_buf }));  // al_ip/PLL.v(57)
  add_pu12_pu12_o12 \u1_Driver/add0  (
    .i0(\u1_Driver/hcnt ),
    .i1(12'b000000000001),
    .o(\u1_Driver/n2 ));  // source/rtl/Driver.v(59)
  add_pu12_pu12_o12 \u1_Driver/add1  (
    .i0(\u1_Driver/vcnt ),
    .i1(12'b000000000001),
    .o(\u1_Driver/n7 ));  // source/rtl/Driver.v(77)
  eq_w12 \u1_Driver/eq0  (
    .i0(\u1_Driver/hcnt ),
    .i1(12'b011010010111),
    .o(\u1_Driver/n5 ));  // source/rtl/Driver.v(72)
  eq_w12 \u1_Driver/eq1  (
    .i0(\u1_Driver/vcnt ),
    .i1(12'b010000101001),
    .o(\u1_Driver/n6 ));  // source/rtl/Driver.v(74)
  lt_u12_u12 \u1_Driver/lt0  (
    .ci(1'b0),
    .i0(\u1_Driver/hcnt ),
    .i1(12'b011010010111),
    .o(\u1_Driver/n1 ));  // source/rtl/Driver.v(58)
  lt_u12_u12 \u1_Driver/lt1  (
    .ci(1'b1),
    .i0(\u1_Driver/hcnt ),
    .i1(12'b000001101111),
    .o(\u1_Driver/n4 ));  // source/rtl/Driver.v(65)
  lt_u12_u12 \u1_Driver/lt2  (
    .ci(1'b1),
    .i0(\u1_Driver/vcnt ),
    .i1(12'b000000000010),
    .o(\u1_Driver/n10 ));  // source/rtl/Driver.v(81)
  lt_u12_u12 \u1_Driver/lt3  (
    .ci(1'b1),
    .i0(12'b000101101000),
    .i1(\u1_Driver/hcnt ),
    .o(\u1_Driver/n11 ));  // source/rtl/Driver.v(87)
  lt_u12_u12 \u1_Driver/lt4  (
    .ci(1'b0),
    .i0(\u1_Driver/hcnt ),
    .i1(12'b011001101000),
    .o(\u1_Driver/n12 ));  // source/rtl/Driver.v(87)
  lt_u12_u12 \u1_Driver/lt5  (
    .ci(1'b1),
    .i0(12'b000000101001),
    .i1(\u1_Driver/vcnt ),
    .o(\u1_Driver/n14 ));  // source/rtl/Driver.v(88)
  lt_u12_u12 \u1_Driver/lt6  (
    .ci(1'b0),
    .i0(\u1_Driver/vcnt ),
    .i1(12'b010000101001),
    .o(\u1_Driver/n15 ));  // source/rtl/Driver.v(88)
  lt_u12_u12 \u1_Driver/lt7  (
    .ci(1'b1),
    .i0(12'b000101100111),
    .i1(\u1_Driver/hcnt ),
    .o(\u1_Driver/n17 ));  // source/rtl/Driver.v(94)
  lt_u12_u12 \u1_Driver/lt8  (
    .ci(1'b0),
    .i0(\u1_Driver/hcnt ),
    .i1(12'b011001100111),
    .o(\u1_Driver/n18 ));  // source/rtl/Driver.v(94)
  binary_mux_s1_w1 \u1_Driver/mux0_b0  (
    .i0(1'b0),
    .i1(\u1_Driver/n2 [0]),
    .sel(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [0]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 \u1_Driver/mux0_b1  (
    .i0(1'b0),
    .i1(\u1_Driver/n2 [1]),
    .sel(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [1]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 \u1_Driver/mux0_b10  (
    .i0(1'b0),
    .i1(\u1_Driver/n2 [10]),
    .sel(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [10]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 \u1_Driver/mux0_b11  (
    .i0(1'b0),
    .i1(\u1_Driver/n2 [11]),
    .sel(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [11]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 \u1_Driver/mux0_b2  (
    .i0(1'b0),
    .i1(\u1_Driver/n2 [2]),
    .sel(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [2]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 \u1_Driver/mux0_b3  (
    .i0(1'b0),
    .i1(\u1_Driver/n2 [3]),
    .sel(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [3]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 \u1_Driver/mux0_b4  (
    .i0(1'b0),
    .i1(\u1_Driver/n2 [4]),
    .sel(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [4]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 \u1_Driver/mux0_b5  (
    .i0(1'b0),
    .i1(\u1_Driver/n2 [5]),
    .sel(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [5]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 \u1_Driver/mux0_b6  (
    .i0(1'b0),
    .i1(\u1_Driver/n2 [6]),
    .sel(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [6]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 \u1_Driver/mux0_b7  (
    .i0(1'b0),
    .i1(\u1_Driver/n2 [7]),
    .sel(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [7]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 \u1_Driver/mux0_b8  (
    .i0(1'b0),
    .i1(\u1_Driver/n2 [8]),
    .sel(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [8]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 \u1_Driver/mux0_b9  (
    .i0(1'b0),
    .i1(\u1_Driver/n2 [9]),
    .sel(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [9]));  // source/rtl/Driver.v(61)
  binary_mux_s1_w1 \u1_Driver/mux1_b0  (
    .i0(\u1_Driver/n7 [0]),
    .i1(1'b0),
    .sel(\u1_Driver/n6 ),
    .o(\u1_Driver/n8 [0]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 \u1_Driver/mux1_b1  (
    .i0(\u1_Driver/n7 [1]),
    .i1(1'b0),
    .sel(\u1_Driver/n6 ),
    .o(\u1_Driver/n8 [1]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 \u1_Driver/mux1_b10  (
    .i0(\u1_Driver/n7 [10]),
    .i1(1'b0),
    .sel(\u1_Driver/n6 ),
    .o(\u1_Driver/n8 [10]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 \u1_Driver/mux1_b11  (
    .i0(\u1_Driver/n7 [11]),
    .i1(1'b0),
    .sel(\u1_Driver/n6 ),
    .o(\u1_Driver/n8 [11]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 \u1_Driver/mux1_b2  (
    .i0(\u1_Driver/n7 [2]),
    .i1(1'b0),
    .sel(\u1_Driver/n6 ),
    .o(\u1_Driver/n8 [2]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 \u1_Driver/mux1_b3  (
    .i0(\u1_Driver/n7 [3]),
    .i1(1'b0),
    .sel(\u1_Driver/n6 ),
    .o(\u1_Driver/n8 [3]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 \u1_Driver/mux1_b4  (
    .i0(\u1_Driver/n7 [4]),
    .i1(1'b0),
    .sel(\u1_Driver/n6 ),
    .o(\u1_Driver/n8 [4]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 \u1_Driver/mux1_b5  (
    .i0(\u1_Driver/n7 [5]),
    .i1(1'b0),
    .sel(\u1_Driver/n6 ),
    .o(\u1_Driver/n8 [5]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 \u1_Driver/mux1_b6  (
    .i0(\u1_Driver/n7 [6]),
    .i1(1'b0),
    .sel(\u1_Driver/n6 ),
    .o(\u1_Driver/n8 [6]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 \u1_Driver/mux1_b7  (
    .i0(\u1_Driver/n7 [7]),
    .i1(1'b0),
    .sel(\u1_Driver/n6 ),
    .o(\u1_Driver/n8 [7]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 \u1_Driver/mux1_b8  (
    .i0(\u1_Driver/n7 [8]),
    .i1(1'b0),
    .sel(\u1_Driver/n6 ),
    .o(\u1_Driver/n8 [8]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 \u1_Driver/mux1_b9  (
    .i0(\u1_Driver/n7 [9]),
    .i1(1'b0),
    .sel(\u1_Driver/n6 ),
    .o(\u1_Driver/n8 [9]));  // source/rtl/Driver.v(77)
  binary_mux_s1_w1 \u1_Driver/mux3_b0  (
    .i0(1'b0),
    .i1(lcd_data[23]),
    .sel(vga_de),
    .o(vga_b[0]));  // source/rtl/Driver.v(91)
  binary_mux_s1_w1 \u1_Driver/mux4_b0  (
    .i0(1'b0),
    .i1(\u1_Driver/n20 [0]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_xpos[0]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 \u1_Driver/mux4_b1  (
    .i0(1'b0),
    .i1(\u1_Driver/n20 [1]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_xpos[1]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 \u1_Driver/mux4_b10  (
    .i0(1'b0),
    .i1(\u1_Driver/n20 [10]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_xpos[10]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 \u1_Driver/mux4_b11  (
    .i0(1'b0),
    .i1(\u1_Driver/n20 [11]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_xpos[11]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 \u1_Driver/mux4_b2  (
    .i0(1'b0),
    .i1(\u1_Driver/n20 [2]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_xpos[2]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 \u1_Driver/mux4_b3  (
    .i0(1'b0),
    .i1(\u1_Driver/n20 [3]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_xpos[3]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 \u1_Driver/mux4_b4  (
    .i0(1'b0),
    .i1(\u1_Driver/n20 [4]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_xpos[4]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 \u1_Driver/mux4_b5  (
    .i0(1'b0),
    .i1(\u1_Driver/n20 [5]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_xpos[5]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 \u1_Driver/mux4_b6  (
    .i0(1'b0),
    .i1(\u1_Driver/n20 [6]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_xpos[6]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 \u1_Driver/mux4_b7  (
    .i0(1'b0),
    .i1(\u1_Driver/n20 [7]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_xpos[7]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 \u1_Driver/mux4_b8  (
    .i0(1'b0),
    .i1(\u1_Driver/n20 [8]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_xpos[8]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 \u1_Driver/mux4_b9  (
    .i0(1'b0),
    .i1(\u1_Driver/n20 [9]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_xpos[9]));  // source/rtl/Driver.v(98)
  binary_mux_s1_w1 \u1_Driver/mux5_b0  (
    .i0(1'b0),
    .i1(\u1_Driver/n21 [0]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_ypos[0]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 \u1_Driver/mux5_b1  (
    .i0(1'b0),
    .i1(\u1_Driver/n21 [1]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_ypos[1]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 \u1_Driver/mux5_b10  (
    .i0(1'b0),
    .i1(\u1_Driver/n21 [10]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_ypos[10]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 \u1_Driver/mux5_b11  (
    .i0(1'b0),
    .i1(\u1_Driver/n21 [11]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_ypos[11]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 \u1_Driver/mux5_b2  (
    .i0(1'b0),
    .i1(\u1_Driver/n21 [2]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_ypos[2]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 \u1_Driver/mux5_b3  (
    .i0(1'b0),
    .i1(\u1_Driver/n21 [3]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_ypos[3]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 \u1_Driver/mux5_b4  (
    .i0(1'b0),
    .i1(\u1_Driver/n21 [4]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_ypos[4]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 \u1_Driver/mux5_b5  (
    .i0(1'b0),
    .i1(\u1_Driver/n21 [5]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_ypos[5]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 \u1_Driver/mux5_b6  (
    .i0(1'b0),
    .i1(\u1_Driver/n21 [6]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_ypos[6]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 \u1_Driver/mux5_b7  (
    .i0(1'b0),
    .i1(\u1_Driver/n21 [7]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_ypos[7]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 \u1_Driver/mux5_b8  (
    .i0(1'b0),
    .i1(\u1_Driver/n21 [8]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_ypos[8]));  // source/rtl/Driver.v(99)
  binary_mux_s1_w1 \u1_Driver/mux5_b9  (
    .i0(1'b0),
    .i1(\u1_Driver/n21 [9]),
    .sel(\u1_Driver/lcd_request ),
    .o(lcd_ypos[9]));  // source/rtl/Driver.v(99)
  reg_ar_as_w1 \u1_Driver/reg0_b0  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [0]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/vcnt [0]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b1  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [1]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/vcnt [1]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b10  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [10]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/vcnt [10]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b11  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [11]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/vcnt [11]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b2  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [2]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/vcnt [2]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b3  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [3]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/vcnt [3]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b4  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [4]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/vcnt [4]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b5  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [5]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/vcnt [5]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b6  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [6]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/vcnt [6]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b7  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [7]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/vcnt [7]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b8  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [8]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/vcnt [8]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b9  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [9]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/vcnt [9]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg1_b0  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [0]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/hcnt [0]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b1  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [1]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/hcnt [1]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b10  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [10]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/hcnt [10]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b11  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [11]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/hcnt [11]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b2  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [2]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/hcnt [2]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b3  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [3]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/hcnt [3]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b4  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [4]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/hcnt [4]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b5  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [5]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/hcnt [5]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b6  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [6]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/hcnt [6]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b7  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [7]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/hcnt [7]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b8  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [8]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/hcnt [8]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b9  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [9]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(\u1_Driver/hcnt [9]));  // source/rtl/Driver.v(62)
  add_pu12_mu12_o12 \u1_Driver/sub0  (
    .i0(\u1_Driver/hcnt ),
    .i1(12'b000101100111),
    .o(\u1_Driver/n20 [11:0]));  // source/rtl/Driver.v(98)
  add_pu12_mu12_o12 \u1_Driver/sub1  (
    .i0(\u1_Driver/vcnt ),
    .i1(12'b000000101001),
    .o(\u1_Driver/n21 [11:0]));  // source/rtl/Driver.v(99)
  and \u1_Driver/u10  (\u1_Driver/lcd_request , \u1_Driver/n19 , \u1_Driver/n16 );  // source/rtl/Driver.v(95)
  not \u1_Driver/u3  (vga_hs, \u1_Driver/n4 );  // source/rtl/Driver.v(65)
  not \u1_Driver/u4  (vga_vs, \u1_Driver/n10 );  // source/rtl/Driver.v(81)
  not \u1_Driver/u5  (vga_clk, clk_vga);  // source/rtl/Driver.v(84)
  and \u1_Driver/u6  (\u1_Driver/n13 , \u1_Driver/n11 , \u1_Driver/n12 );  // source/rtl/Driver.v(87)
  and \u1_Driver/u7  (\u1_Driver/n16 , \u1_Driver/n14 , \u1_Driver/n15 );  // source/rtl/Driver.v(88)
  and \u1_Driver/u8  (vga_de, \u1_Driver/n13 , \u1_Driver/n16 );  // source/rtl/Driver.v(88)
  and \u1_Driver/u9  (\u1_Driver/n19 , \u1_Driver/n17 , \u1_Driver/n18 );  // source/rtl/Driver.v(94)
  add_pu31_pu31_o31 \u2_Display/add0  (
    .i0(\u2_Display/n ),
    .i1(31'b0000000000000000000000000000001),
    .o(\u2_Display/n37 ));  // source/rtl/Display.v(60)
  add_pu32_pu32_o32 \u2_Display/add1  (
    .i0(\u2_Display/counta ),
    .i1(32'b00000000000000000000000000000001),
    .o(\u2_Display/n41 ));  // source/rtl/Display.v(155)
  add_pu32_pu32_pu1_o32 \u2_Display/add100  (
    .i0({\u2_Display/n3191 ,\u2_Display/n3192 ,\u2_Display/n3193 ,\u2_Display/n3194 ,\u2_Display/n3195 ,\u2_Display/n3196 ,\u2_Display/n3197 ,\u2_Display/n3198 ,\u2_Display/n3199 ,\u2_Display/n3200 ,\u2_Display/n3201 ,\u2_Display/n3202 ,\u2_Display/n3203 ,\u2_Display/n3204 ,\u2_Display/n3205 ,\u2_Display/n3206 ,\u2_Display/n3207 ,\u2_Display/n3208 ,\u2_Display/n3209 ,\u2_Display/n3210 ,\u2_Display/n3211 ,\u2_Display/n3212 ,\u2_Display/n3213 ,\u2_Display/n3214 ,\u2_Display/n3215 ,\u2_Display/n3216 ,\u2_Display/n3217 ,\u2_Display/n3218 ,\u2_Display/n3219 ,\u2_Display/n3220 ,\u2_Display/n3221 ,\u2_Display/n3222 }),
    .i1(32'b11111111111111110110100111111111),
    .i2(1'b1),
    .o(\u2_Display/n3225 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add101  (
    .i0({\u2_Display/n3226 ,\u2_Display/n3227 ,\u2_Display/n3228 ,\u2_Display/n3229 ,\u2_Display/n3230 ,\u2_Display/n3231 ,\u2_Display/n3232 ,\u2_Display/n3233 ,\u2_Display/n3234 ,\u2_Display/n3235 ,\u2_Display/n3236 ,\u2_Display/n3237 ,\u2_Display/n3238 ,\u2_Display/n3239 ,\u2_Display/n3240 ,\u2_Display/n3241 ,\u2_Display/n3242 ,\u2_Display/n3243 ,\u2_Display/n3244 ,\u2_Display/n3245 ,\u2_Display/n3246 ,\u2_Display/n3247 ,\u2_Display/n3248 ,\u2_Display/n3249 ,\u2_Display/n3250 ,\u2_Display/n3251 ,\u2_Display/n3252 ,\u2_Display/n3253 ,\u2_Display/n3254 ,\u2_Display/n3255 ,\u2_Display/n3256 ,\u2_Display/n3257 }),
    .i1(32'b11111111111111111011010011111111),
    .i2(1'b1),
    .o(\u2_Display/n3260 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add102  (
    .i0({\u2_Display/n3261 ,\u2_Display/n3262 ,\u2_Display/n3263 ,\u2_Display/n3264 ,\u2_Display/n3265 ,\u2_Display/n3266 ,\u2_Display/n3267 ,\u2_Display/n3268 ,\u2_Display/n3269 ,\u2_Display/n3270 ,\u2_Display/n3271 ,\u2_Display/n3272 ,\u2_Display/n3273 ,\u2_Display/n3274 ,\u2_Display/n3275 ,\u2_Display/n3276 ,\u2_Display/n3277 ,\u2_Display/n3278 ,\u2_Display/n3279 ,\u2_Display/n3280 ,\u2_Display/n3281 ,\u2_Display/n3282 ,\u2_Display/n3283 ,\u2_Display/n3284 ,\u2_Display/n3285 ,\u2_Display/n3286 ,\u2_Display/n3287 ,\u2_Display/n3288 ,\u2_Display/n3289 ,\u2_Display/n3290 ,\u2_Display/n3291 ,\u2_Display/n3292 }),
    .i1(32'b11111111111111111101101001111111),
    .i2(1'b1),
    .o(\u2_Display/n3295 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add103  (
    .i0({\u2_Display/n3296 ,\u2_Display/n3297 ,\u2_Display/n3298 ,\u2_Display/n3299 ,\u2_Display/n3300 ,\u2_Display/n3301 ,\u2_Display/n3302 ,\u2_Display/n3303 ,\u2_Display/n3304 ,\u2_Display/n3305 ,\u2_Display/n3306 ,\u2_Display/n3307 ,\u2_Display/n3308 ,\u2_Display/n3309 ,\u2_Display/n3310 ,\u2_Display/n3311 ,\u2_Display/n3312 ,\u2_Display/n3313 ,\u2_Display/n3314 ,\u2_Display/n3315 ,\u2_Display/n3316 ,\u2_Display/n3317 ,\u2_Display/n3318 ,\u2_Display/n3319 ,\u2_Display/n3320 ,\u2_Display/n3321 ,\u2_Display/n3322 ,\u2_Display/n3323 ,\u2_Display/n3324 ,\u2_Display/n3325 ,\u2_Display/n3326 ,\u2_Display/n3327 }),
    .i1(32'b11111111111111111110110100111111),
    .i2(1'b1),
    .o(\u2_Display/n3330 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add104  (
    .i0({\u2_Display/n3331 ,\u2_Display/n3332 ,\u2_Display/n3333 ,\u2_Display/n3334 ,\u2_Display/n3335 ,\u2_Display/n3336 ,\u2_Display/n3337 ,\u2_Display/n3338 ,\u2_Display/n3339 ,\u2_Display/n3340 ,\u2_Display/n3341 ,\u2_Display/n3342 ,\u2_Display/n3343 ,\u2_Display/n3344 ,\u2_Display/n3345 ,\u2_Display/n3346 ,\u2_Display/n3347 ,\u2_Display/n3348 ,\u2_Display/n3349 ,\u2_Display/n3350 ,\u2_Display/n3351 ,\u2_Display/n3352 ,\u2_Display/n3353 ,\u2_Display/n3354 ,\u2_Display/n3355 ,\u2_Display/n3356 ,\u2_Display/n3357 ,\u2_Display/n3358 ,\u2_Display/n3359 ,\u2_Display/n3360 ,\u2_Display/n3361 ,\u2_Display/n3362 }),
    .i1(32'b11111111111111111111011010011111),
    .i2(1'b1),
    .o(\u2_Display/n3365 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add105  (
    .i0({\u2_Display/n3366 ,\u2_Display/n3367 ,\u2_Display/n3368 ,\u2_Display/n3369 ,\u2_Display/n3370 ,\u2_Display/n3371 ,\u2_Display/n3372 ,\u2_Display/n3373 ,\u2_Display/n3374 ,\u2_Display/n3375 ,\u2_Display/n3376 ,\u2_Display/n3377 ,\u2_Display/n3378 ,\u2_Display/n3379 ,\u2_Display/n3380 ,\u2_Display/n3381 ,\u2_Display/n3382 ,\u2_Display/n3383 ,\u2_Display/n3384 ,\u2_Display/n3385 ,\u2_Display/n3386 ,\u2_Display/n3387 ,\u2_Display/n3388 ,\u2_Display/n3389 ,\u2_Display/n3390 ,\u2_Display/n3391 ,\u2_Display/n3392 ,\u2_Display/n3393 ,\u2_Display/n3394 ,\u2_Display/n3395 ,\u2_Display/n3396 ,\u2_Display/n3397 }),
    .i1(32'b11111111111111111111101101001111),
    .i2(1'b1),
    .o(\u2_Display/n3400 ));  // source/rtl/Display.v(196)
  add_pu10_pu10_pu1_o10 \u2_Display/add106  (
    .i0({\u2_Display/n3423 ,\u2_Display/n3424 ,\u2_Display/n3425 ,\u2_Display/n3426 ,\u2_Display/n3427 ,\u2_Display/n3428 ,\u2_Display/n3429 ,\u2_Display/n3430 ,\u2_Display/n3431 ,\u2_Display/n3432 }),
    .i1(10'b0110100111),
    .i2(1'b1),
    .o(\u2_Display/n3435 [9:0]));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add117  (
    .i0(\u2_Display/counta ),
    .i1(32'b00110111111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n3788 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add118  (
    .i0({\u2_Display/n3789 ,\u2_Display/n3790 ,\u2_Display/n3791 ,\u2_Display/n3792 ,\u2_Display/n3793 ,\u2_Display/n3794 ,\u2_Display/n3795 ,\u2_Display/n3796 ,\u2_Display/n3797 ,\u2_Display/n3798 ,\u2_Display/n3799 ,\u2_Display/n3800 ,\u2_Display/n3801 ,\u2_Display/n3802 ,\u2_Display/n3803 ,\u2_Display/n3804 ,\u2_Display/n3805 ,\u2_Display/n3806 ,\u2_Display/n3807 ,\u2_Display/n3808 ,\u2_Display/n3809 ,\u2_Display/n3810 ,\u2_Display/n3811 ,\u2_Display/n3812 ,\u2_Display/n3813 ,\u2_Display/n3814 ,\u2_Display/n3815 ,\u2_Display/n3816 ,\u2_Display/n3817 ,\u2_Display/n3818 ,\u2_Display/n3819 ,\u2_Display/n3820 }),
    .i1(32'b10011011111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n3823 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add119  (
    .i0({\u2_Display/n3824 ,\u2_Display/n3825 ,\u2_Display/n3826 ,\u2_Display/n3827 ,\u2_Display/n3828 ,\u2_Display/n3829 ,\u2_Display/n3830 ,\u2_Display/n3831 ,\u2_Display/n3832 ,\u2_Display/n3833 ,\u2_Display/n3834 ,\u2_Display/n3835 ,\u2_Display/n3836 ,\u2_Display/n3837 ,\u2_Display/n3838 ,\u2_Display/n3839 ,\u2_Display/n3840 ,\u2_Display/n3841 ,\u2_Display/n3842 ,\u2_Display/n3843 ,\u2_Display/n3844 ,\u2_Display/n3845 ,\u2_Display/n3846 ,\u2_Display/n3847 ,\u2_Display/n3848 ,\u2_Display/n3849 ,\u2_Display/n3850 ,\u2_Display/n3851 ,\u2_Display/n3852 ,\u2_Display/n3853 ,\u2_Display/n3854 ,\u2_Display/n3855 }),
    .i1(32'b11001101111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n3858 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add120  (
    .i0({\u2_Display/n3859 ,\u2_Display/n3860 ,\u2_Display/n3861 ,\u2_Display/n3862 ,\u2_Display/n3863 ,\u2_Display/n3864 ,\u2_Display/n3865 ,\u2_Display/n3866 ,\u2_Display/n3867 ,\u2_Display/n3868 ,\u2_Display/n3869 ,\u2_Display/n3870 ,\u2_Display/n3871 ,\u2_Display/n3872 ,\u2_Display/n3873 ,\u2_Display/n3874 ,\u2_Display/n3875 ,\u2_Display/n3876 ,\u2_Display/n3877 ,\u2_Display/n3878 ,\u2_Display/n3879 ,\u2_Display/n3880 ,\u2_Display/n3881 ,\u2_Display/n3882 ,\u2_Display/n3883 ,\u2_Display/n3884 ,\u2_Display/n3885 ,\u2_Display/n3886 ,\u2_Display/n3887 ,\u2_Display/n3888 ,\u2_Display/n3889 ,\u2_Display/n3890 }),
    .i1(32'b11100110111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n3893 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add121  (
    .i0({\u2_Display/n3894 ,\u2_Display/n3895 ,\u2_Display/n3896 ,\u2_Display/n3897 ,\u2_Display/n3898 ,\u2_Display/n3899 ,\u2_Display/n3900 ,\u2_Display/n3901 ,\u2_Display/n3902 ,\u2_Display/n3903 ,\u2_Display/n3904 ,\u2_Display/n3905 ,\u2_Display/n3906 ,\u2_Display/n3907 ,\u2_Display/n3908 ,\u2_Display/n3909 ,\u2_Display/n3910 ,\u2_Display/n3911 ,\u2_Display/n3912 ,\u2_Display/n3913 ,\u2_Display/n3914 ,\u2_Display/n3915 ,\u2_Display/n3916 ,\u2_Display/n3917 ,\u2_Display/n3918 ,\u2_Display/n3919 ,\u2_Display/n3920 ,\u2_Display/n3921 ,\u2_Display/n3922 ,\u2_Display/n3923 ,\u2_Display/n3924 ,\u2_Display/n3925 }),
    .i1(32'b11110011011111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n3928 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add122  (
    .i0({\u2_Display/n3929 ,\u2_Display/n3930 ,\u2_Display/n3931 ,\u2_Display/n3932 ,\u2_Display/n3933 ,\u2_Display/n3934 ,\u2_Display/n3935 ,\u2_Display/n3936 ,\u2_Display/n3937 ,\u2_Display/n3938 ,\u2_Display/n3939 ,\u2_Display/n3940 ,\u2_Display/n3941 ,\u2_Display/n3942 ,\u2_Display/n3943 ,\u2_Display/n3944 ,\u2_Display/n3945 ,\u2_Display/n3946 ,\u2_Display/n3947 ,\u2_Display/n3948 ,\u2_Display/n3949 ,\u2_Display/n3950 ,\u2_Display/n3951 ,\u2_Display/n3952 ,\u2_Display/n3953 ,\u2_Display/n3954 ,\u2_Display/n3955 ,\u2_Display/n3956 ,\u2_Display/n3957 ,\u2_Display/n3958 ,\u2_Display/n3959 ,\u2_Display/n3960 }),
    .i1(32'b11111001101111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n3963 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add123  (
    .i0({\u2_Display/n3964 ,\u2_Display/n3965 ,\u2_Display/n3966 ,\u2_Display/n3967 ,\u2_Display/n3968 ,\u2_Display/n3969 ,\u2_Display/n3970 ,\u2_Display/n3971 ,\u2_Display/n3972 ,\u2_Display/n3973 ,\u2_Display/n3974 ,\u2_Display/n3975 ,\u2_Display/n3976 ,\u2_Display/n3977 ,\u2_Display/n3978 ,\u2_Display/n3979 ,\u2_Display/n3980 ,\u2_Display/n3981 ,\u2_Display/n3982 ,\u2_Display/n3983 ,\u2_Display/n3984 ,\u2_Display/n3985 ,\u2_Display/n3986 ,\u2_Display/n3987 ,\u2_Display/n3988 ,\u2_Display/n3989 ,\u2_Display/n3990 ,\u2_Display/n3991 ,\u2_Display/n3992 ,\u2_Display/n3993 ,\u2_Display/n3994 ,\u2_Display/n3995 }),
    .i1(32'b11111100110111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n3998 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add124  (
    .i0({\u2_Display/n3999 ,\u2_Display/n4000 ,\u2_Display/n4001 ,\u2_Display/n4002 ,\u2_Display/n4003 ,\u2_Display/n4004 ,\u2_Display/n4005 ,\u2_Display/n4006 ,\u2_Display/n4007 ,\u2_Display/n4008 ,\u2_Display/n4009 ,\u2_Display/n4010 ,\u2_Display/n4011 ,\u2_Display/n4012 ,\u2_Display/n4013 ,\u2_Display/n4014 ,\u2_Display/n4015 ,\u2_Display/n4016 ,\u2_Display/n4017 ,\u2_Display/n4018 ,\u2_Display/n4019 ,\u2_Display/n4020 ,\u2_Display/n4021 ,\u2_Display/n4022 ,\u2_Display/n4023 ,\u2_Display/n4024 ,\u2_Display/n4025 ,\u2_Display/n4026 ,\u2_Display/n4027 ,\u2_Display/n4028 ,\u2_Display/n4029 ,\u2_Display/n4030 }),
    .i1(32'b11111110011011111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n4033 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add125  (
    .i0({\u2_Display/n4034 ,\u2_Display/n4035 ,\u2_Display/n4036 ,\u2_Display/n4037 ,\u2_Display/n4038 ,\u2_Display/n4039 ,\u2_Display/n4040 ,\u2_Display/n4041 ,\u2_Display/n4042 ,\u2_Display/n4043 ,\u2_Display/n4044 ,\u2_Display/n4045 ,\u2_Display/n4046 ,\u2_Display/n4047 ,\u2_Display/n4048 ,\u2_Display/n4049 ,\u2_Display/n4050 ,\u2_Display/n4051 ,\u2_Display/n4052 ,\u2_Display/n4053 ,\u2_Display/n4054 ,\u2_Display/n4055 ,\u2_Display/n4056 ,\u2_Display/n4057 ,\u2_Display/n4058 ,\u2_Display/n4059 ,\u2_Display/n4060 ,\u2_Display/n4061 ,\u2_Display/n4062 ,\u2_Display/n4063 ,\u2_Display/n4064 ,\u2_Display/n4065 }),
    .i1(32'b11111111001101111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n4068 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add126  (
    .i0({\u2_Display/n4069 ,\u2_Display/n4070 ,\u2_Display/n4071 ,\u2_Display/n4072 ,\u2_Display/n4073 ,\u2_Display/n4074 ,\u2_Display/n4075 ,\u2_Display/n4076 ,\u2_Display/n4077 ,\u2_Display/n4078 ,\u2_Display/n4079 ,\u2_Display/n4080 ,\u2_Display/n4081 ,\u2_Display/n4082 ,\u2_Display/n4083 ,\u2_Display/n4084 ,\u2_Display/n4085 ,\u2_Display/n4086 ,\u2_Display/n4087 ,\u2_Display/n4088 ,\u2_Display/n4089 ,\u2_Display/n4090 ,\u2_Display/n4091 ,\u2_Display/n4092 ,\u2_Display/n4093 ,\u2_Display/n4094 ,\u2_Display/n4095 ,\u2_Display/n4096 ,\u2_Display/n4097 ,\u2_Display/n4098 ,\u2_Display/n4099 ,\u2_Display/n4100 }),
    .i1(32'b11111111100110111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n4103 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add127  (
    .i0({\u2_Display/n4104 ,\u2_Display/n4105 ,\u2_Display/n4106 ,\u2_Display/n4107 ,\u2_Display/n4108 ,\u2_Display/n4109 ,\u2_Display/n4110 ,\u2_Display/n4111 ,\u2_Display/n4112 ,\u2_Display/n4113 ,\u2_Display/n4114 ,\u2_Display/n4115 ,\u2_Display/n4116 ,\u2_Display/n4117 ,\u2_Display/n4118 ,\u2_Display/n4119 ,\u2_Display/n4120 ,\u2_Display/n4121 ,\u2_Display/n4122 ,\u2_Display/n4123 ,\u2_Display/n4124 ,\u2_Display/n4125 ,\u2_Display/n4126 ,\u2_Display/n4127 ,\u2_Display/n4128 ,\u2_Display/n4129 ,\u2_Display/n4130 ,\u2_Display/n4131 ,\u2_Display/n4132 ,\u2_Display/n4133 ,\u2_Display/n4134 ,\u2_Display/n4135 }),
    .i1(32'b11111111110011011111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n4138 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add128  (
    .i0({\u2_Display/n4139 ,\u2_Display/n4140 ,\u2_Display/n4141 ,\u2_Display/n4142 ,\u2_Display/n4143 ,\u2_Display/n4144 ,\u2_Display/n4145 ,\u2_Display/n4146 ,\u2_Display/n4147 ,\u2_Display/n4148 ,\u2_Display/n4149 ,\u2_Display/n4150 ,\u2_Display/n4151 ,\u2_Display/n4152 ,\u2_Display/n4153 ,\u2_Display/n4154 ,\u2_Display/n4155 ,\u2_Display/n4156 ,\u2_Display/n4157 ,\u2_Display/n4158 ,\u2_Display/n4159 ,\u2_Display/n4160 ,\u2_Display/n4161 ,\u2_Display/n4162 ,\u2_Display/n4163 ,\u2_Display/n4164 ,\u2_Display/n4165 ,\u2_Display/n4166 ,\u2_Display/n4167 ,\u2_Display/n4168 ,\u2_Display/n4169 ,\u2_Display/n4170 }),
    .i1(32'b11111111111001101111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n4173 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add129  (
    .i0({\u2_Display/n4174 ,\u2_Display/n4175 ,\u2_Display/n4176 ,\u2_Display/n4177 ,\u2_Display/n4178 ,\u2_Display/n4179 ,\u2_Display/n4180 ,\u2_Display/n4181 ,\u2_Display/n4182 ,\u2_Display/n4183 ,\u2_Display/n4184 ,\u2_Display/n4185 ,\u2_Display/n4186 ,\u2_Display/n4187 ,\u2_Display/n4188 ,\u2_Display/n4189 ,\u2_Display/n4190 ,\u2_Display/n4191 ,\u2_Display/n4192 ,\u2_Display/n4193 ,\u2_Display/n4194 ,\u2_Display/n4195 ,\u2_Display/n4196 ,\u2_Display/n4197 ,\u2_Display/n4198 ,\u2_Display/n4199 ,\u2_Display/n4200 ,\u2_Display/n4201 ,\u2_Display/n4202 ,\u2_Display/n4203 ,\u2_Display/n4204 ,\u2_Display/n4205 }),
    .i1(32'b11111111111100110111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n4208 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add130  (
    .i0({\u2_Display/n4209 ,\u2_Display/n4210 ,\u2_Display/n4211 ,\u2_Display/n4212 ,\u2_Display/n4213 ,\u2_Display/n4214 ,\u2_Display/n4215 ,\u2_Display/n4216 ,\u2_Display/n4217 ,\u2_Display/n4218 ,\u2_Display/n4219 ,\u2_Display/n4220 ,\u2_Display/n4221 ,\u2_Display/n4222 ,\u2_Display/n4223 ,\u2_Display/n4224 ,\u2_Display/n4225 ,\u2_Display/n4226 ,\u2_Display/n4227 ,\u2_Display/n4228 ,\u2_Display/n4229 ,\u2_Display/n4230 ,\u2_Display/n4231 ,\u2_Display/n4232 ,\u2_Display/n4233 ,\u2_Display/n4234 ,\u2_Display/n4235 ,\u2_Display/n4236 ,\u2_Display/n4237 ,\u2_Display/n4238 ,\u2_Display/n4239 ,\u2_Display/n4240 }),
    .i1(32'b11111111111110011011111111111111),
    .i2(1'b1),
    .o(\u2_Display/n4243 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add131  (
    .i0({\u2_Display/n4244 ,\u2_Display/n4245 ,\u2_Display/n4246 ,\u2_Display/n4247 ,\u2_Display/n4248 ,\u2_Display/n4249 ,\u2_Display/n4250 ,\u2_Display/n4251 ,\u2_Display/n4252 ,\u2_Display/n4253 ,\u2_Display/n4254 ,\u2_Display/n4255 ,\u2_Display/n4256 ,\u2_Display/n4257 ,\u2_Display/n4258 ,\u2_Display/n4259 ,\u2_Display/n4260 ,\u2_Display/n4261 ,\u2_Display/n4262 ,\u2_Display/n4263 ,\u2_Display/n4264 ,\u2_Display/n4265 ,\u2_Display/n4266 ,\u2_Display/n4267 ,\u2_Display/n4268 ,\u2_Display/n4269 ,\u2_Display/n4270 ,\u2_Display/n4271 ,\u2_Display/n4272 ,\u2_Display/n4273 ,\u2_Display/n4274 ,\u2_Display/n4275 }),
    .i1(32'b11111111111111001101111111111111),
    .i2(1'b1),
    .o(\u2_Display/n4278 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add132  (
    .i0({\u2_Display/n4279 ,\u2_Display/n4280 ,\u2_Display/n4281 ,\u2_Display/n4282 ,\u2_Display/n4283 ,\u2_Display/n4284 ,\u2_Display/n4285 ,\u2_Display/n4286 ,\u2_Display/n4287 ,\u2_Display/n4288 ,\u2_Display/n4289 ,\u2_Display/n4290 ,\u2_Display/n4291 ,\u2_Display/n4292 ,\u2_Display/n4293 ,\u2_Display/n4294 ,\u2_Display/n4295 ,\u2_Display/n4296 ,\u2_Display/n4297 ,\u2_Display/n4298 ,\u2_Display/n4299 ,\u2_Display/n4300 ,\u2_Display/n4301 ,\u2_Display/n4302 ,\u2_Display/n4303 ,\u2_Display/n4304 ,\u2_Display/n4305 ,\u2_Display/n4306 ,\u2_Display/n4307 ,\u2_Display/n4308 ,\u2_Display/n4309 ,\u2_Display/n4310 }),
    .i1(32'b11111111111111100110111111111111),
    .i2(1'b1),
    .o(\u2_Display/n4313 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add133  (
    .i0({\u2_Display/n4314 ,\u2_Display/n4315 ,\u2_Display/n4316 ,\u2_Display/n4317 ,\u2_Display/n4318 ,\u2_Display/n4319 ,\u2_Display/n4320 ,\u2_Display/n4321 ,\u2_Display/n4322 ,\u2_Display/n4323 ,\u2_Display/n4324 ,\u2_Display/n4325 ,\u2_Display/n4326 ,\u2_Display/n4327 ,\u2_Display/n4328 ,\u2_Display/n4329 ,\u2_Display/n4330 ,\u2_Display/n4331 ,\u2_Display/n4332 ,\u2_Display/n4333 ,\u2_Display/n4334 ,\u2_Display/n4335 ,\u2_Display/n4336 ,\u2_Display/n4337 ,\u2_Display/n4338 ,\u2_Display/n4339 ,\u2_Display/n4340 ,\u2_Display/n4341 ,\u2_Display/n4342 ,\u2_Display/n4343 ,\u2_Display/n4344 ,\u2_Display/n4345 }),
    .i1(32'b11111111111111110011011111111111),
    .i2(1'b1),
    .o(\u2_Display/n4348 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add134  (
    .i0({\u2_Display/n4349 ,\u2_Display/n4350 ,\u2_Display/n4351 ,\u2_Display/n4352 ,\u2_Display/n4353 ,\u2_Display/n4354 ,\u2_Display/n4355 ,\u2_Display/n4356 ,\u2_Display/n4357 ,\u2_Display/n4358 ,\u2_Display/n4359 ,\u2_Display/n4360 ,\u2_Display/n4361 ,\u2_Display/n4362 ,\u2_Display/n4363 ,\u2_Display/n4364 ,\u2_Display/n4365 ,\u2_Display/n4366 ,\u2_Display/n4367 ,\u2_Display/n4368 ,\u2_Display/n4369 ,\u2_Display/n4370 ,\u2_Display/n4371 ,\u2_Display/n4372 ,\u2_Display/n4373 ,\u2_Display/n4374 ,\u2_Display/n4375 ,\u2_Display/n4376 ,\u2_Display/n4377 ,\u2_Display/n4378 ,\u2_Display/n4379 ,\u2_Display/n4380 }),
    .i1(32'b11111111111111111001101111111111),
    .i2(1'b1),
    .o(\u2_Display/n4383 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add135  (
    .i0({\u2_Display/n4384 ,\u2_Display/n4385 ,\u2_Display/n4386 ,\u2_Display/n4387 ,\u2_Display/n4388 ,\u2_Display/n4389 ,\u2_Display/n4390 ,\u2_Display/n4391 ,\u2_Display/n4392 ,\u2_Display/n4393 ,\u2_Display/n4394 ,\u2_Display/n4395 ,\u2_Display/n4396 ,\u2_Display/n4397 ,\u2_Display/n4398 ,\u2_Display/n4399 ,\u2_Display/n4400 ,\u2_Display/n4401 ,\u2_Display/n4402 ,\u2_Display/n4403 ,\u2_Display/n4404 ,\u2_Display/n4405 ,\u2_Display/n4406 ,\u2_Display/n4407 ,\u2_Display/n4408 ,\u2_Display/n4409 ,\u2_Display/n4410 ,\u2_Display/n4411 ,\u2_Display/n4412 ,\u2_Display/n4413 ,\u2_Display/n4414 ,\u2_Display/n4415 }),
    .i1(32'b11111111111111111100110111111111),
    .i2(1'b1),
    .o(\u2_Display/n4418 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add136  (
    .i0({\u2_Display/n4419 ,\u2_Display/n4420 ,\u2_Display/n4421 ,\u2_Display/n4422 ,\u2_Display/n4423 ,\u2_Display/n4424 ,\u2_Display/n4425 ,\u2_Display/n4426 ,\u2_Display/n4427 ,\u2_Display/n4428 ,\u2_Display/n4429 ,\u2_Display/n4430 ,\u2_Display/n4431 ,\u2_Display/n4432 ,\u2_Display/n4433 ,\u2_Display/n4434 ,\u2_Display/n4435 ,\u2_Display/n4436 ,\u2_Display/n4437 ,\u2_Display/n4438 ,\u2_Display/n4439 ,\u2_Display/n4440 ,\u2_Display/n4441 ,\u2_Display/n4442 ,\u2_Display/n4443 ,\u2_Display/n4444 ,\u2_Display/n4445 ,\u2_Display/n4446 ,\u2_Display/n4447 ,\u2_Display/n4448 ,\u2_Display/n4449 ,\u2_Display/n4450 }),
    .i1(32'b11111111111111111110011011111111),
    .i2(1'b1),
    .o(\u2_Display/n4453 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add137  (
    .i0({\u2_Display/n4454 ,\u2_Display/n4455 ,\u2_Display/n4456 ,\u2_Display/n4457 ,\u2_Display/n4458 ,\u2_Display/n4459 ,\u2_Display/n4460 ,\u2_Display/n4461 ,\u2_Display/n4462 ,\u2_Display/n4463 ,\u2_Display/n4464 ,\u2_Display/n4465 ,\u2_Display/n4466 ,\u2_Display/n4467 ,\u2_Display/n4468 ,\u2_Display/n4469 ,\u2_Display/n4470 ,\u2_Display/n4471 ,\u2_Display/n4472 ,\u2_Display/n4473 ,\u2_Display/n4474 ,\u2_Display/n4475 ,\u2_Display/n4476 ,\u2_Display/n4477 ,\u2_Display/n4478 ,\u2_Display/n4479 ,\u2_Display/n4480 ,\u2_Display/n4481 ,\u2_Display/n4482 ,\u2_Display/n4483 ,\u2_Display/n4484 ,\u2_Display/n4485 }),
    .i1(32'b11111111111111111111001101111111),
    .i2(1'b1),
    .o(\u2_Display/n4488 ));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add138  (
    .i0({\u2_Display/n4489 ,\u2_Display/n4490 ,\u2_Display/n4491 ,\u2_Display/n4492 ,\u2_Display/n4493 ,\u2_Display/n4494 ,\u2_Display/n4495 ,\u2_Display/n4496 ,\u2_Display/n4497 ,\u2_Display/n4498 ,\u2_Display/n4499 ,\u2_Display/n4500 ,\u2_Display/n4501 ,\u2_Display/n4502 ,\u2_Display/n4503 ,\u2_Display/n4504 ,\u2_Display/n4505 ,\u2_Display/n4506 ,\u2_Display/n4507 ,\u2_Display/n4508 ,\u2_Display/n4509 ,\u2_Display/n4510 ,\u2_Display/n4511 ,\u2_Display/n4512 ,\u2_Display/n4513 ,\u2_Display/n4514 ,\u2_Display/n4515 ,\u2_Display/n4516 ,\u2_Display/n4517 ,\u2_Display/n4518 ,\u2_Display/n4519 ,\u2_Display/n4520 }),
    .i1(32'b11111111111111111111100110111111),
    .i2(1'b1),
    .o(\u2_Display/n4523 ));  // source/rtl/Display.v(195)
  add_pu10_pu10_pu1_o10 \u2_Display/add139  (
    .i0({\u2_Display/n4546 ,\u2_Display/n4547 ,\u2_Display/n4548 ,\u2_Display/n4549 ,\u2_Display/n4550 ,\u2_Display/n4551 ,\u2_Display/n4552 ,\u2_Display/n4553 ,\u2_Display/n4554 ,\u2_Display/n4555 }),
    .i1(10'b0011011111),
    .i2(1'b1),
    .o(\u2_Display/n4558 [9:0]));  // source/rtl/Display.v(195)
  add_pu32_pu32_pu1_o32 \u2_Display/add14  (
    .i0(\u2_Display/counta ),
    .i1(32'b01011111111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n4911 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add151  (
    .i0({\u2_Display/n6070 ,\u2_Display/n6071 ,\u2_Display/n6072 ,\u2_Display/n6073 ,\u2_Display/n6074 ,\u2_Display/n6075 ,\u2_Display/n6076 ,\u2_Display/n6077 ,\u2_Display/n6078 ,\u2_Display/n6079 ,\u2_Display/n6080 ,\u2_Display/n6081 ,\u2_Display/n6082 ,\u2_Display/n6083 ,\u2_Display/n6084 ,\u2_Display/n6085 ,\u2_Display/n6086 ,\u2_Display/n6087 ,\u2_Display/n6088 ,\u2_Display/n6089 ,\u2_Display/n6090 ,\u2_Display/n6091 ,\u2_Display/n6092 ,\u2_Display/n6093 ,\u2_Display/n6094 ,\u2_Display/n6095 ,\u2_Display/n6096 ,\u2_Display/n6097 ,\u2_Display/n6098 ,\u2_Display/n6099 ,\u2_Display/n6100 ,\u2_Display/n6101 }),
    .i1(32'b10101111111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n4946 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add152  (
    .i0({\u2_Display/n6105 ,\u2_Display/n6106 ,\u2_Display/n6107 ,\u2_Display/n6108 ,\u2_Display/n6109 ,\u2_Display/n6110 ,\u2_Display/n6111 ,\u2_Display/n6112 ,\u2_Display/n6113 ,\u2_Display/n6114 ,\u2_Display/n6115 ,\u2_Display/n6116 ,\u2_Display/n6117 ,\u2_Display/n6118 ,\u2_Display/n6119 ,\u2_Display/n6120 ,\u2_Display/n6121 ,\u2_Display/n6122 ,\u2_Display/n6123 ,\u2_Display/n6124 ,\u2_Display/n6125 ,\u2_Display/n6126 ,\u2_Display/n6127 ,\u2_Display/n6128 ,\u2_Display/n6129 ,\u2_Display/n6130 ,\u2_Display/n6131 ,\u2_Display/n6132 ,\u2_Display/n6133 ,\u2_Display/n6134 ,\u2_Display/n6135 ,\u2_Display/n6136 }),
    .i1(32'b11010111111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n4981 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add153  (
    .i0({\u2_Display/n6140 ,\u2_Display/n6141 ,\u2_Display/n6142 ,\u2_Display/n6143 ,\u2_Display/n6144 ,\u2_Display/n6145 ,\u2_Display/n6146 ,\u2_Display/n6147 ,\u2_Display/n6148 ,\u2_Display/n6149 ,\u2_Display/n6150 ,\u2_Display/n6151 ,\u2_Display/n6152 ,\u2_Display/n6153 ,\u2_Display/n6154 ,\u2_Display/n6155 ,\u2_Display/n6156 ,\u2_Display/n6157 ,\u2_Display/n6158 ,\u2_Display/n6159 ,\u2_Display/n6160 ,\u2_Display/n6161 ,\u2_Display/n6162 ,\u2_Display/n6163 ,\u2_Display/n6164 ,\u2_Display/n6165 ,\u2_Display/n6166 ,\u2_Display/n6167 ,\u2_Display/n6168 ,\u2_Display/n6169 ,\u2_Display/n6170 ,\u2_Display/n6171 }),
    .i1(32'b11101011111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5016 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add154  (
    .i0({\u2_Display/n6175 ,\u2_Display/n6176 ,\u2_Display/n6177 ,\u2_Display/n6178 ,\u2_Display/n6179 ,\u2_Display/n6180 ,\u2_Display/n6181 ,\u2_Display/n6182 ,\u2_Display/n6183 ,\u2_Display/n6184 ,\u2_Display/n6185 ,\u2_Display/n6186 ,\u2_Display/n6187 ,\u2_Display/n6188 ,\u2_Display/n6189 ,\u2_Display/n6190 ,\u2_Display/n6191 ,\u2_Display/n6192 ,\u2_Display/n6193 ,\u2_Display/n6194 ,\u2_Display/n6195 ,\u2_Display/n6196 ,\u2_Display/n6197 ,\u2_Display/n6198 ,\u2_Display/n6199 ,\u2_Display/n6200 ,\u2_Display/n6201 ,\u2_Display/n6202 ,\u2_Display/n6203 ,\u2_Display/n6204 ,\u2_Display/n6205 ,\u2_Display/n6206 }),
    .i1(32'b11110101111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5051 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add155  (
    .i0({\u2_Display/n6210 ,\u2_Display/n6211 ,\u2_Display/n6212 ,\u2_Display/n6213 ,\u2_Display/n6214 ,\u2_Display/n6215 ,\u2_Display/n6216 ,\u2_Display/n6217 ,\u2_Display/n6218 ,\u2_Display/n6219 ,\u2_Display/n6220 ,\u2_Display/n6221 ,\u2_Display/n6222 ,\u2_Display/n6223 ,\u2_Display/n6224 ,\u2_Display/n6225 ,\u2_Display/n6226 ,\u2_Display/n6227 ,\u2_Display/n6228 ,\u2_Display/n6229 ,\u2_Display/n6230 ,\u2_Display/n6231 ,\u2_Display/n6232 ,\u2_Display/n6233 ,\u2_Display/n6234 ,\u2_Display/n6235 ,\u2_Display/n6236 ,\u2_Display/n6237 ,\u2_Display/n6238 ,\u2_Display/n6239 ,\u2_Display/n6240 ,\u2_Display/n6241 }),
    .i1(32'b11111010111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5086 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add156  (
    .i0({\u2_Display/n6245 ,\u2_Display/n6246 ,\u2_Display/n6247 ,\u2_Display/n6248 ,\u2_Display/n6249 ,\u2_Display/n6250 ,\u2_Display/n6251 ,\u2_Display/n6252 ,\u2_Display/n6253 ,\u2_Display/n6254 ,\u2_Display/n6255 ,\u2_Display/n6256 ,\u2_Display/n6257 ,\u2_Display/n6258 ,\u2_Display/n6259 ,\u2_Display/n6260 ,\u2_Display/n6261 ,\u2_Display/n6262 ,\u2_Display/n6263 ,\u2_Display/n6264 ,\u2_Display/n6265 ,\u2_Display/n6266 ,\u2_Display/n6267 ,\u2_Display/n6268 ,\u2_Display/n6269 ,\u2_Display/n6270 ,\u2_Display/n6271 ,\u2_Display/n6272 ,\u2_Display/n6273 ,\u2_Display/n6274 ,\u2_Display/n6275 ,\u2_Display/n6276 }),
    .i1(32'b11111101011111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5121 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add157  (
    .i0({\u2_Display/n6280 ,\u2_Display/n6281 ,\u2_Display/n6282 ,\u2_Display/n6283 ,\u2_Display/n6284 ,\u2_Display/n6285 ,\u2_Display/n6286 ,\u2_Display/n6287 ,\u2_Display/n6288 ,\u2_Display/n6289 ,\u2_Display/n6290 ,\u2_Display/n6291 ,\u2_Display/n6292 ,\u2_Display/n6293 ,\u2_Display/n6294 ,\u2_Display/n6295 ,\u2_Display/n6296 ,\u2_Display/n6297 ,\u2_Display/n6298 ,\u2_Display/n6299 ,\u2_Display/n6300 ,\u2_Display/n6301 ,\u2_Display/n6302 ,\u2_Display/n6303 ,\u2_Display/n6304 ,\u2_Display/n6305 ,\u2_Display/n6306 ,\u2_Display/n6307 ,\u2_Display/n6308 ,\u2_Display/n6309 ,\u2_Display/n6310 ,\u2_Display/n6311 }),
    .i1(32'b11111110101111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5156 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add158  (
    .i0({\u2_Display/n6315 ,\u2_Display/n6316 ,\u2_Display/n6317 ,\u2_Display/n6318 ,\u2_Display/n6319 ,\u2_Display/n6320 ,\u2_Display/n6321 ,\u2_Display/n6322 ,\u2_Display/n6323 ,\u2_Display/n6324 ,\u2_Display/n6325 ,\u2_Display/n6326 ,\u2_Display/n6327 ,\u2_Display/n6328 ,\u2_Display/n6329 ,\u2_Display/n6330 ,\u2_Display/n6331 ,\u2_Display/n6332 ,\u2_Display/n6333 ,\u2_Display/n6334 ,\u2_Display/n6335 ,\u2_Display/n6336 ,\u2_Display/n6337 ,\u2_Display/n6338 ,\u2_Display/n6339 ,\u2_Display/n6340 ,\u2_Display/n6341 ,\u2_Display/n6342 ,\u2_Display/n6343 ,\u2_Display/n6344 ,\u2_Display/n6345 ,\u2_Display/n6346 }),
    .i1(32'b11111111010111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5191 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add159  (
    .i0({\u2_Display/n6350 ,\u2_Display/n6351 ,\u2_Display/n6352 ,\u2_Display/n6353 ,\u2_Display/n5196 ,\u2_Display/n5197 ,\u2_Display/n5198 ,\u2_Display/n5199 ,\u2_Display/n5200 ,\u2_Display/n5201 ,\u2_Display/n5202 ,\u2_Display/n5203 ,\u2_Display/n5204 ,\u2_Display/n5205 ,\u2_Display/n5206 ,\u2_Display/n5207 ,\u2_Display/n5208 ,\u2_Display/n5209 ,\u2_Display/n5210 ,\u2_Display/n5211 ,\u2_Display/n5212 ,\u2_Display/n5213 ,\u2_Display/n5214 ,\u2_Display/n5215 ,\u2_Display/n5216 ,\u2_Display/n5217 ,\u2_Display/n5218 ,\u2_Display/n5219 ,\u2_Display/n5220 ,\u2_Display/n5221 ,\u2_Display/n5222 ,\u2_Display/n5223 }),
    .i1(32'b11111111101011111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5226 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add160  (
    .i0({\u2_Display/n5227 ,\u2_Display/n5228 ,\u2_Display/n5229 ,\u2_Display/n5230 ,\u2_Display/n5231 ,\u2_Display/n5232 ,\u2_Display/n5233 ,\u2_Display/n5234 ,\u2_Display/n5235 ,\u2_Display/n5236 ,\u2_Display/n5237 ,\u2_Display/n5238 ,\u2_Display/n5239 ,\u2_Display/n5240 ,\u2_Display/n5241 ,\u2_Display/n5242 ,\u2_Display/n5243 ,\u2_Display/n5244 ,\u2_Display/n5245 ,\u2_Display/n5246 ,\u2_Display/n5247 ,\u2_Display/n5248 ,\u2_Display/n5249 ,\u2_Display/n5250 ,\u2_Display/n5251 ,\u2_Display/n5252 ,\u2_Display/n5253 ,\u2_Display/n5254 ,\u2_Display/n5255 ,\u2_Display/n5256 ,\u2_Display/n5257 ,\u2_Display/n5258 }),
    .i1(32'b11111111110101111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5261 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add161  (
    .i0({\u2_Display/n5262 ,\u2_Display/n5263 ,\u2_Display/n5264 ,\u2_Display/n5265 ,\u2_Display/n5266 ,\u2_Display/n5267 ,\u2_Display/n5268 ,\u2_Display/n5269 ,\u2_Display/n5270 ,\u2_Display/n5271 ,\u2_Display/n5272 ,\u2_Display/n5273 ,\u2_Display/n5274 ,\u2_Display/n5275 ,\u2_Display/n5276 ,\u2_Display/n5277 ,\u2_Display/n5278 ,\u2_Display/n5279 ,\u2_Display/n5280 ,\u2_Display/n5281 ,\u2_Display/n5282 ,\u2_Display/n5283 ,\u2_Display/n5284 ,\u2_Display/n5285 ,\u2_Display/n5286 ,\u2_Display/n5287 ,\u2_Display/n5288 ,\u2_Display/n5289 ,\u2_Display/n5290 ,\u2_Display/n5291 ,\u2_Display/n5292 ,\u2_Display/n5293 }),
    .i1(32'b11111111111010111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5296 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add162  (
    .i0({\u2_Display/n5297 ,\u2_Display/n5298 ,\u2_Display/n5299 ,\u2_Display/n5300 ,\u2_Display/n5301 ,\u2_Display/n5302 ,\u2_Display/n5303 ,\u2_Display/n5304 ,\u2_Display/n5305 ,\u2_Display/n5306 ,\u2_Display/n5307 ,\u2_Display/n5308 ,\u2_Display/n5309 ,\u2_Display/n5310 ,\u2_Display/n5311 ,\u2_Display/n5312 ,\u2_Display/n5313 ,\u2_Display/n5314 ,\u2_Display/n5315 ,\u2_Display/n5316 ,\u2_Display/n5317 ,\u2_Display/n5318 ,\u2_Display/n5319 ,\u2_Display/n5320 ,\u2_Display/n5321 ,\u2_Display/n5322 ,\u2_Display/n5323 ,\u2_Display/n5324 ,\u2_Display/n5325 ,\u2_Display/n5326 ,\u2_Display/n5327 ,\u2_Display/n5328 }),
    .i1(32'b11111111111101011111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5331 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add163  (
    .i0({\u2_Display/n5332 ,\u2_Display/n5333 ,\u2_Display/n5334 ,\u2_Display/n5335 ,\u2_Display/n5336 ,\u2_Display/n5337 ,\u2_Display/n5338 ,\u2_Display/n5339 ,\u2_Display/n5340 ,\u2_Display/n5341 ,\u2_Display/n5342 ,\u2_Display/n5343 ,\u2_Display/n5344 ,\u2_Display/n5345 ,\u2_Display/n5346 ,\u2_Display/n5347 ,\u2_Display/n5348 ,\u2_Display/n5349 ,\u2_Display/n5350 ,\u2_Display/n5351 ,\u2_Display/n5352 ,\u2_Display/n5353 ,\u2_Display/n5354 ,\u2_Display/n5355 ,\u2_Display/n5356 ,\u2_Display/n5357 ,\u2_Display/n5358 ,\u2_Display/n5359 ,\u2_Display/n5360 ,\u2_Display/n5361 ,\u2_Display/n5362 ,\u2_Display/n5363 }),
    .i1(32'b11111111111110101111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5366 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add164  (
    .i0({\u2_Display/n5367 ,\u2_Display/n5368 ,\u2_Display/n5369 ,\u2_Display/n5370 ,\u2_Display/n5371 ,\u2_Display/n5372 ,\u2_Display/n5373 ,\u2_Display/n5374 ,\u2_Display/n5375 ,\u2_Display/n5376 ,\u2_Display/n5377 ,\u2_Display/n5378 ,\u2_Display/n5379 ,\u2_Display/n5380 ,\u2_Display/n5381 ,\u2_Display/n5382 ,\u2_Display/n5383 ,\u2_Display/n5384 ,\u2_Display/n5385 ,\u2_Display/n5386 ,\u2_Display/n5387 ,\u2_Display/n5388 ,\u2_Display/n5389 ,\u2_Display/n5390 ,\u2_Display/n5391 ,\u2_Display/n5392 ,\u2_Display/n5393 ,\u2_Display/n5394 ,\u2_Display/n5395 ,\u2_Display/n5396 ,\u2_Display/n5397 ,\u2_Display/n5398 }),
    .i1(32'b11111111111111010111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5401 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add165  (
    .i0({\u2_Display/n5402 ,\u2_Display/n5403 ,\u2_Display/n5404 ,\u2_Display/n5405 ,\u2_Display/n5406 ,\u2_Display/n5407 ,\u2_Display/n5408 ,\u2_Display/n5409 ,\u2_Display/n5410 ,\u2_Display/n5411 ,\u2_Display/n5412 ,\u2_Display/n5413 ,\u2_Display/n5414 ,\u2_Display/n5415 ,\u2_Display/n5416 ,\u2_Display/n5417 ,\u2_Display/n5418 ,\u2_Display/n5419 ,\u2_Display/n5420 ,\u2_Display/n5421 ,\u2_Display/n5422 ,\u2_Display/n5423 ,\u2_Display/n5424 ,\u2_Display/n5425 ,\u2_Display/n5426 ,\u2_Display/n5427 ,\u2_Display/n5428 ,\u2_Display/n5429 ,\u2_Display/n5430 ,\u2_Display/n5431 ,\u2_Display/n5432 ,\u2_Display/n5433 }),
    .i1(32'b11111111111111101011111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5436 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add166  (
    .i0({\u2_Display/n5437 ,\u2_Display/n5438 ,\u2_Display/n5439 ,\u2_Display/n5440 ,\u2_Display/n5441 ,\u2_Display/n5442 ,\u2_Display/n5443 ,\u2_Display/n5444 ,\u2_Display/n5445 ,\u2_Display/n5446 ,\u2_Display/n5447 ,\u2_Display/n5448 ,\u2_Display/n5449 ,\u2_Display/n5450 ,\u2_Display/n5451 ,\u2_Display/n5452 ,\u2_Display/n5453 ,\u2_Display/n5454 ,\u2_Display/n5455 ,\u2_Display/n5456 ,\u2_Display/n5457 ,\u2_Display/n5458 ,\u2_Display/n5459 ,\u2_Display/n5460 ,\u2_Display/n5461 ,\u2_Display/n5462 ,\u2_Display/n5463 ,\u2_Display/n5464 ,\u2_Display/n5465 ,\u2_Display/n5466 ,\u2_Display/n5467 ,\u2_Display/n5468 }),
    .i1(32'b11111111111111110101111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5471 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add167  (
    .i0({\u2_Display/n5472 ,\u2_Display/n5473 ,\u2_Display/n5474 ,\u2_Display/n5475 ,\u2_Display/n5476 ,\u2_Display/n5477 ,\u2_Display/n5478 ,\u2_Display/n5479 ,\u2_Display/n5480 ,\u2_Display/n5481 ,\u2_Display/n5482 ,\u2_Display/n5483 ,\u2_Display/n5484 ,\u2_Display/n5485 ,\u2_Display/n5486 ,\u2_Display/n5487 ,\u2_Display/n5488 ,\u2_Display/n5489 ,\u2_Display/n5490 ,\u2_Display/n5491 ,\u2_Display/n5492 ,\u2_Display/n5493 ,\u2_Display/n5494 ,\u2_Display/n5495 ,\u2_Display/n5496 ,\u2_Display/n5497 ,\u2_Display/n5498 ,\u2_Display/n5499 ,\u2_Display/n5500 ,\u2_Display/n5501 ,\u2_Display/n5502 ,\u2_Display/n5503 }),
    .i1(32'b11111111111111111010111111111111),
    .i2(1'b1),
    .o(\u2_Display/n5506 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add168  (
    .i0({\u2_Display/n5507 ,\u2_Display/n5508 ,\u2_Display/n5509 ,\u2_Display/n5510 ,\u2_Display/n5511 ,\u2_Display/n5512 ,\u2_Display/n5513 ,\u2_Display/n5514 ,\u2_Display/n5515 ,\u2_Display/n5516 ,\u2_Display/n5517 ,\u2_Display/n5518 ,\u2_Display/n5519 ,\u2_Display/n5520 ,\u2_Display/n5521 ,\u2_Display/n5522 ,\u2_Display/n5523 ,\u2_Display/n5524 ,\u2_Display/n5525 ,\u2_Display/n5526 ,\u2_Display/n5527 ,\u2_Display/n5528 ,\u2_Display/n5529 ,\u2_Display/n5530 ,\u2_Display/n5531 ,\u2_Display/n5532 ,\u2_Display/n5533 ,\u2_Display/n5534 ,\u2_Display/n5535 ,\u2_Display/n5536 ,\u2_Display/n5537 ,\u2_Display/n5538 }),
    .i1(32'b11111111111111111101011111111111),
    .i2(1'b1),
    .o(\u2_Display/n5541 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add169  (
    .i0({\u2_Display/n5542 ,\u2_Display/n5543 ,\u2_Display/n5544 ,\u2_Display/n5545 ,\u2_Display/n5546 ,\u2_Display/n5547 ,\u2_Display/n5548 ,\u2_Display/n5549 ,\u2_Display/n5550 ,\u2_Display/n5551 ,\u2_Display/n5552 ,\u2_Display/n5553 ,\u2_Display/n5554 ,\u2_Display/n5555 ,\u2_Display/n5556 ,\u2_Display/n5557 ,\u2_Display/n5558 ,\u2_Display/n5559 ,\u2_Display/n5560 ,\u2_Display/n5561 ,\u2_Display/n5562 ,\u2_Display/n5563 ,\u2_Display/n5564 ,\u2_Display/n5565 ,\u2_Display/n5566 ,\u2_Display/n5567 ,\u2_Display/n5568 ,\u2_Display/n5569 ,\u2_Display/n5570 ,\u2_Display/n5571 ,\u2_Display/n5572 ,\u2_Display/n5573 }),
    .i1(32'b11111111111111111110101111111111),
    .i2(1'b1),
    .o(\u2_Display/n5576 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add170  (
    .i0({\u2_Display/n5577 ,\u2_Display/n5578 ,\u2_Display/n5579 ,\u2_Display/n5580 ,\u2_Display/n5581 ,\u2_Display/n5582 ,\u2_Display/n5583 ,\u2_Display/n5584 ,\u2_Display/n5585 ,\u2_Display/n5586 ,\u2_Display/n5587 ,\u2_Display/n5588 ,\u2_Display/n5589 ,\u2_Display/n5590 ,\u2_Display/n5591 ,\u2_Display/n5592 ,\u2_Display/n5593 ,\u2_Display/n5594 ,\u2_Display/n5595 ,\u2_Display/n5596 ,\u2_Display/n5597 ,\u2_Display/n5598 ,\u2_Display/n5599 ,\u2_Display/n5600 ,\u2_Display/n5601 ,\u2_Display/n5602 ,\u2_Display/n5603 ,\u2_Display/n5604 ,\u2_Display/n5605 ,\u2_Display/n5606 ,\u2_Display/n5607 ,\u2_Display/n5608 }),
    .i1(32'b11111111111111111111010111111111),
    .i2(1'b1),
    .o(\u2_Display/n5611 ));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add171  (
    .i0({\u2_Display/n5612 ,\u2_Display/n5613 ,\u2_Display/n5614 ,\u2_Display/n5615 ,\u2_Display/n5616 ,\u2_Display/n5617 ,\u2_Display/n5618 ,\u2_Display/n5619 ,\u2_Display/n5620 ,\u2_Display/n5621 ,\u2_Display/n5622 ,\u2_Display/n5623 ,\u2_Display/n5624 ,\u2_Display/n5625 ,\u2_Display/n5626 ,\u2_Display/n5627 ,\u2_Display/n5628 ,\u2_Display/n5629 ,\u2_Display/n5630 ,\u2_Display/n5631 ,\u2_Display/n5632 ,\u2_Display/n5633 ,\u2_Display/n5634 ,\u2_Display/n5635 ,\u2_Display/n5636 ,\u2_Display/n5637 ,\u2_Display/n5638 ,\u2_Display/n5639 ,\u2_Display/n5640 ,\u2_Display/n5641 ,\u2_Display/n5642 ,\u2_Display/n5643 }),
    .i1(32'b11111111111111111111101011111111),
    .i2(1'b1),
    .o(\u2_Display/n5646 ));  // source/rtl/Display.v(179)
  add_pu10_pu10_pu1_o10 \u2_Display/add172  (
    .i0({\u2_Display/n5669 ,\u2_Display/n5670 ,\u2_Display/n5671 ,\u2_Display/n5672 ,\u2_Display/n5673 ,\u2_Display/n5674 ,\u2_Display/n5675 ,\u2_Display/n5676 ,\u2_Display/n5677 ,\u2_Display/n5678 }),
    .i1(10'b0101111111),
    .i2(1'b1),
    .o(\u2_Display/n5681 [9:0]));  // source/rtl/Display.v(179)
  add_pu32_pu32_pu1_o32 \u2_Display/add18  (
    .i0(\u2_Display/counta ),
    .i1(32'b00000101111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n419 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add19  (
    .i0({\u2_Display/n420 ,\u2_Display/n421 ,\u2_Display/n422 ,\u2_Display/n423 ,\u2_Display/n424 ,\u2_Display/n425 ,\u2_Display/n426 ,\u2_Display/n427 ,\u2_Display/n428 ,\u2_Display/n429 ,\u2_Display/n430 ,\u2_Display/n431 ,\u2_Display/n432 ,\u2_Display/n433 ,\u2_Display/n434 ,\u2_Display/n435 ,\u2_Display/n436 ,\u2_Display/n437 ,\u2_Display/n438 ,\u2_Display/n439 ,\u2_Display/n440 ,\u2_Display/n441 ,\u2_Display/n442 ,\u2_Display/n443 ,\u2_Display/n444 ,\u2_Display/n445 ,\u2_Display/n446 ,\u2_Display/n447 ,\u2_Display/n448 ,\u2_Display/n449 ,\u2_Display/n450 ,\u2_Display/n451 }),
    .i1(32'b10000010111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n454 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add20  (
    .i0({\u2_Display/n455 ,\u2_Display/n456 ,\u2_Display/n457 ,\u2_Display/n458 ,\u2_Display/n459 ,\u2_Display/n460 ,\u2_Display/n461 ,\u2_Display/n462 ,\u2_Display/n463 ,\u2_Display/n464 ,\u2_Display/n465 ,\u2_Display/n466 ,\u2_Display/n467 ,\u2_Display/n468 ,\u2_Display/n469 ,\u2_Display/n470 ,\u2_Display/n471 ,\u2_Display/n472 ,\u2_Display/n473 ,\u2_Display/n474 ,\u2_Display/n475 ,\u2_Display/n476 ,\u2_Display/n477 ,\u2_Display/n478 ,\u2_Display/n479 ,\u2_Display/n480 ,\u2_Display/n481 ,\u2_Display/n482 ,\u2_Display/n483 ,\u2_Display/n484 ,\u2_Display/n485 ,\u2_Display/n486 }),
    .i1(32'b11000001011111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n489 ));  // source/rtl/Display.v(230)
  add_pu11_pu11_pu1_o11 \u2_Display/add205  (
    .i0({\u2_Display/n5633 ,\u2_Display/n5634 ,\u2_Display/n5635 ,\u2_Display/n5636 ,\u2_Display/n5637 ,\u2_Display/n5638 ,\u2_Display/n5639 ,\u2_Display/n5640 ,\u2_Display/n5641 ,\u2_Display/n5642 ,\u2_Display/n5643 }),
    .i1(11'b01011111111),
    .i2(1'b1),
    .o(\u2_Display/n6804 [10:0]));  // source/rtl/Display.v(163)
  add_pu32_pu32_pu1_o32 \u2_Display/add21  (
    .i0({\u2_Display/n490 ,\u2_Display/n491 ,\u2_Display/n492 ,\u2_Display/n493 ,\u2_Display/n494 ,\u2_Display/n495 ,\u2_Display/n496 ,\u2_Display/n497 ,\u2_Display/n498 ,\u2_Display/n499 ,\u2_Display/n500 ,\u2_Display/n501 ,\u2_Display/n502 ,\u2_Display/n503 ,\u2_Display/n504 ,\u2_Display/n505 ,\u2_Display/n506 ,\u2_Display/n507 ,\u2_Display/n508 ,\u2_Display/n509 ,\u2_Display/n510 ,\u2_Display/n511 ,\u2_Display/n512 ,\u2_Display/n513 ,\u2_Display/n514 ,\u2_Display/n515 ,\u2_Display/n516 ,\u2_Display/n517 ,\u2_Display/n518 ,\u2_Display/n519 ,\u2_Display/n520 ,\u2_Display/n521 }),
    .i1(32'b11100000101111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n524 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add22  (
    .i0({\u2_Display/n525 ,\u2_Display/n526 ,\u2_Display/n527 ,\u2_Display/n528 ,\u2_Display/n529 ,\u2_Display/n530 ,\u2_Display/n531 ,\u2_Display/n532 ,\u2_Display/n533 ,\u2_Display/n534 ,\u2_Display/n535 ,\u2_Display/n536 ,\u2_Display/n537 ,\u2_Display/n538 ,\u2_Display/n539 ,\u2_Display/n540 ,\u2_Display/n541 ,\u2_Display/n542 ,\u2_Display/n543 ,\u2_Display/n544 ,\u2_Display/n545 ,\u2_Display/n546 ,\u2_Display/n547 ,\u2_Display/n548 ,\u2_Display/n549 ,\u2_Display/n550 ,\u2_Display/n551 ,\u2_Display/n552 ,\u2_Display/n553 ,\u2_Display/n554 ,\u2_Display/n555 ,\u2_Display/n556 }),
    .i1(32'b11110000010111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n559 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add23  (
    .i0({\u2_Display/n560 ,\u2_Display/n561 ,\u2_Display/n562 ,\u2_Display/n563 ,\u2_Display/n564 ,\u2_Display/n565 ,\u2_Display/n566 ,\u2_Display/n567 ,\u2_Display/n568 ,\u2_Display/n569 ,\u2_Display/n570 ,\u2_Display/n571 ,\u2_Display/n572 ,\u2_Display/n573 ,\u2_Display/n574 ,\u2_Display/n575 ,\u2_Display/n576 ,\u2_Display/n577 ,\u2_Display/n578 ,\u2_Display/n579 ,\u2_Display/n580 ,\u2_Display/n581 ,\u2_Display/n582 ,\u2_Display/n583 ,\u2_Display/n584 ,\u2_Display/n585 ,\u2_Display/n586 ,\u2_Display/n587 ,\u2_Display/n588 ,\u2_Display/n589 ,\u2_Display/n590 ,\u2_Display/n591 }),
    .i1(32'b11111000001011111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n594 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add24  (
    .i0({\u2_Display/n595 ,\u2_Display/n596 ,\u2_Display/n597 ,\u2_Display/n598 ,\u2_Display/n599 ,\u2_Display/n600 ,\u2_Display/n601 ,\u2_Display/n602 ,\u2_Display/n603 ,\u2_Display/n604 ,\u2_Display/n605 ,\u2_Display/n606 ,\u2_Display/n607 ,\u2_Display/n608 ,\u2_Display/n609 ,\u2_Display/n610 ,\u2_Display/n611 ,\u2_Display/n612 ,\u2_Display/n613 ,\u2_Display/n614 ,\u2_Display/n615 ,\u2_Display/n616 ,\u2_Display/n617 ,\u2_Display/n618 ,\u2_Display/n619 ,\u2_Display/n620 ,\u2_Display/n621 ,\u2_Display/n622 ,\u2_Display/n623 ,\u2_Display/n624 ,\u2_Display/n625 ,\u2_Display/n626 }),
    .i1(32'b11111100000101111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n629 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add25  (
    .i0({\u2_Display/n630 ,\u2_Display/n631 ,\u2_Display/n632 ,\u2_Display/n633 ,\u2_Display/n634 ,\u2_Display/n635 ,\u2_Display/n636 ,\u2_Display/n637 ,\u2_Display/n638 ,\u2_Display/n639 ,\u2_Display/n640 ,\u2_Display/n641 ,\u2_Display/n642 ,\u2_Display/n643 ,\u2_Display/n644 ,\u2_Display/n645 ,\u2_Display/n646 ,\u2_Display/n647 ,\u2_Display/n648 ,\u2_Display/n649 ,\u2_Display/n650 ,\u2_Display/n651 ,\u2_Display/n652 ,\u2_Display/n653 ,\u2_Display/n654 ,\u2_Display/n655 ,\u2_Display/n656 ,\u2_Display/n657 ,\u2_Display/n658 ,\u2_Display/n659 ,\u2_Display/n660 ,\u2_Display/n661 }),
    .i1(32'b11111110000010111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n664 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add26  (
    .i0({\u2_Display/n665 ,\u2_Display/n666 ,\u2_Display/n667 ,\u2_Display/n668 ,\u2_Display/n669 ,\u2_Display/n670 ,\u2_Display/n671 ,\u2_Display/n672 ,\u2_Display/n673 ,\u2_Display/n674 ,\u2_Display/n675 ,\u2_Display/n676 ,\u2_Display/n677 ,\u2_Display/n678 ,\u2_Display/n679 ,\u2_Display/n680 ,\u2_Display/n681 ,\u2_Display/n682 ,\u2_Display/n683 ,\u2_Display/n684 ,\u2_Display/n685 ,\u2_Display/n686 ,\u2_Display/n687 ,\u2_Display/n688 ,\u2_Display/n689 ,\u2_Display/n690 ,\u2_Display/n691 ,\u2_Display/n692 ,\u2_Display/n693 ,\u2_Display/n694 ,\u2_Display/n695 ,\u2_Display/n696 }),
    .i1(32'b11111111000001011111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n699 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add27  (
    .i0({\u2_Display/n700 ,\u2_Display/n701 ,\u2_Display/n702 ,\u2_Display/n703 ,\u2_Display/n704 ,\u2_Display/n705 ,\u2_Display/n706 ,\u2_Display/n707 ,\u2_Display/n708 ,\u2_Display/n709 ,\u2_Display/n710 ,\u2_Display/n711 ,\u2_Display/n712 ,\u2_Display/n713 ,\u2_Display/n714 ,\u2_Display/n715 ,\u2_Display/n716 ,\u2_Display/n717 ,\u2_Display/n718 ,\u2_Display/n719 ,\u2_Display/n720 ,\u2_Display/n721 ,\u2_Display/n722 ,\u2_Display/n723 ,\u2_Display/n724 ,\u2_Display/n725 ,\u2_Display/n726 ,\u2_Display/n727 ,\u2_Display/n728 ,\u2_Display/n729 ,\u2_Display/n730 ,\u2_Display/n731 }),
    .i1(32'b11111111100000101111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n734 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add28  (
    .i0({\u2_Display/n735 ,\u2_Display/n736 ,\u2_Display/n737 ,\u2_Display/n738 ,\u2_Display/n739 ,\u2_Display/n740 ,\u2_Display/n741 ,\u2_Display/n742 ,\u2_Display/n743 ,\u2_Display/n744 ,\u2_Display/n745 ,\u2_Display/n746 ,\u2_Display/n747 ,\u2_Display/n748 ,\u2_Display/n749 ,\u2_Display/n750 ,\u2_Display/n751 ,\u2_Display/n752 ,\u2_Display/n753 ,\u2_Display/n754 ,\u2_Display/n755 ,\u2_Display/n756 ,\u2_Display/n757 ,\u2_Display/n758 ,\u2_Display/n759 ,\u2_Display/n760 ,\u2_Display/n761 ,\u2_Display/n762 ,\u2_Display/n763 ,\u2_Display/n764 ,\u2_Display/n765 ,\u2_Display/n766 }),
    .i1(32'b11111111110000010111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n769 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add29  (
    .i0({\u2_Display/n770 ,\u2_Display/n771 ,\u2_Display/n772 ,\u2_Display/n773 ,\u2_Display/n774 ,\u2_Display/n775 ,\u2_Display/n776 ,\u2_Display/n777 ,\u2_Display/n778 ,\u2_Display/n779 ,\u2_Display/n780 ,\u2_Display/n781 ,\u2_Display/n782 ,\u2_Display/n783 ,\u2_Display/n784 ,\u2_Display/n785 ,\u2_Display/n786 ,\u2_Display/n787 ,\u2_Display/n788 ,\u2_Display/n789 ,\u2_Display/n790 ,\u2_Display/n791 ,\u2_Display/n792 ,\u2_Display/n793 ,\u2_Display/n794 ,\u2_Display/n795 ,\u2_Display/n796 ,\u2_Display/n797 ,\u2_Display/n798 ,\u2_Display/n799 ,\u2_Display/n800 ,\u2_Display/n801 }),
    .i1(32'b11111111111000001011111111111111),
    .i2(1'b1),
    .o(\u2_Display/n804 ));  // source/rtl/Display.v(230)
  add_pu3_pu3_o4 \u2_Display/add2_2  (
    .i0(3'b101),
    .i1(\u2_Display/i [10:8]),
    .o({\u2_Display/add2_2_co ,\u2_Display/n43 [2:0]}));  // source/rtl/Display.v(165)
  add_pu32_pu32_pu1_o32 \u2_Display/add30  (
    .i0({\u2_Display/n805 ,\u2_Display/n806 ,\u2_Display/n807 ,\u2_Display/n808 ,\u2_Display/n809 ,\u2_Display/n810 ,\u2_Display/n811 ,\u2_Display/n812 ,\u2_Display/n813 ,\u2_Display/n814 ,\u2_Display/n815 ,\u2_Display/n816 ,\u2_Display/n817 ,\u2_Display/n818 ,\u2_Display/n819 ,\u2_Display/n820 ,\u2_Display/n821 ,\u2_Display/n822 ,\u2_Display/n823 ,\u2_Display/n824 ,\u2_Display/n825 ,\u2_Display/n826 ,\u2_Display/n827 ,\u2_Display/n828 ,\u2_Display/n829 ,\u2_Display/n830 ,\u2_Display/n831 ,\u2_Display/n832 ,\u2_Display/n833 ,\u2_Display/n834 ,\u2_Display/n835 ,\u2_Display/n836 }),
    .i1(32'b11111111111100000101111111111111),
    .i2(1'b1),
    .o(\u2_Display/n839 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add31  (
    .i0({\u2_Display/n840 ,\u2_Display/n841 ,\u2_Display/n842 ,\u2_Display/n843 ,\u2_Display/n844 ,\u2_Display/n845 ,\u2_Display/n846 ,\u2_Display/n847 ,\u2_Display/n848 ,\u2_Display/n849 ,\u2_Display/n850 ,\u2_Display/n851 ,\u2_Display/n852 ,\u2_Display/n853 ,\u2_Display/n854 ,\u2_Display/n855 ,\u2_Display/n856 ,\u2_Display/n857 ,\u2_Display/n858 ,\u2_Display/n859 ,\u2_Display/n860 ,\u2_Display/n861 ,\u2_Display/n862 ,\u2_Display/n863 ,\u2_Display/n864 ,\u2_Display/n865 ,\u2_Display/n866 ,\u2_Display/n867 ,\u2_Display/n868 ,\u2_Display/n869 ,\u2_Display/n870 ,\u2_Display/n871 }),
    .i1(32'b11111111111110000010111111111111),
    .i2(1'b1),
    .o(\u2_Display/n874 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add32  (
    .i0({\u2_Display/n875 ,\u2_Display/n876 ,\u2_Display/n877 ,\u2_Display/n878 ,\u2_Display/n879 ,\u2_Display/n880 ,\u2_Display/n881 ,\u2_Display/n882 ,\u2_Display/n883 ,\u2_Display/n884 ,\u2_Display/n885 ,\u2_Display/n886 ,\u2_Display/n887 ,\u2_Display/n888 ,\u2_Display/n889 ,\u2_Display/n890 ,\u2_Display/n891 ,\u2_Display/n892 ,\u2_Display/n893 ,\u2_Display/n894 ,\u2_Display/n895 ,\u2_Display/n896 ,\u2_Display/n897 ,\u2_Display/n898 ,\u2_Display/n899 ,\u2_Display/n900 ,\u2_Display/n901 ,\u2_Display/n902 ,\u2_Display/n903 ,\u2_Display/n904 ,\u2_Display/n905 ,\u2_Display/n906 }),
    .i1(32'b11111111111111000001011111111111),
    .i2(1'b1),
    .o(\u2_Display/n909 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add33  (
    .i0({\u2_Display/n910 ,\u2_Display/n911 ,\u2_Display/n912 ,\u2_Display/n913 ,\u2_Display/n914 ,\u2_Display/n915 ,\u2_Display/n916 ,\u2_Display/n917 ,\u2_Display/n918 ,\u2_Display/n919 ,\u2_Display/n920 ,\u2_Display/n921 ,\u2_Display/n922 ,\u2_Display/n923 ,\u2_Display/n924 ,\u2_Display/n925 ,\u2_Display/n926 ,\u2_Display/n927 ,\u2_Display/n928 ,\u2_Display/n929 ,\u2_Display/n930 ,\u2_Display/n931 ,\u2_Display/n932 ,\u2_Display/n933 ,\u2_Display/n934 ,\u2_Display/n935 ,\u2_Display/n936 ,\u2_Display/n937 ,\u2_Display/n938 ,\u2_Display/n939 ,\u2_Display/n940 ,\u2_Display/n941 }),
    .i1(32'b11111111111111100000101111111111),
    .i2(1'b1),
    .o(\u2_Display/n944 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add34  (
    .i0({\u2_Display/n945 ,\u2_Display/n946 ,\u2_Display/n947 ,\u2_Display/n948 ,\u2_Display/n949 ,\u2_Display/n950 ,\u2_Display/n951 ,\u2_Display/n952 ,\u2_Display/n953 ,\u2_Display/n954 ,\u2_Display/n955 ,\u2_Display/n956 ,\u2_Display/n957 ,\u2_Display/n958 ,\u2_Display/n959 ,\u2_Display/n960 ,\u2_Display/n961 ,\u2_Display/n962 ,\u2_Display/n963 ,\u2_Display/n964 ,\u2_Display/n965 ,\u2_Display/n966 ,\u2_Display/n967 ,\u2_Display/n968 ,\u2_Display/n969 ,\u2_Display/n970 ,\u2_Display/n971 ,\u2_Display/n972 ,\u2_Display/n973 ,\u2_Display/n974 ,\u2_Display/n975 ,\u2_Display/n976 }),
    .i1(32'b11111111111111110000010111111111),
    .i2(1'b1),
    .o(\u2_Display/n979 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add35  (
    .i0({\u2_Display/n980 ,\u2_Display/n981 ,\u2_Display/n982 ,\u2_Display/n983 ,\u2_Display/n984 ,\u2_Display/n985 ,\u2_Display/n986 ,\u2_Display/n987 ,\u2_Display/n988 ,\u2_Display/n989 ,\u2_Display/n990 ,\u2_Display/n991 ,\u2_Display/n992 ,\u2_Display/n993 ,\u2_Display/n994 ,\u2_Display/n995 ,\u2_Display/n996 ,\u2_Display/n997 ,\u2_Display/n998 ,\u2_Display/n999 ,\u2_Display/n1000 ,\u2_Display/n1001 ,\u2_Display/n1002 ,\u2_Display/n1003 ,\u2_Display/n1004 ,\u2_Display/n1005 ,\u2_Display/n1006 ,\u2_Display/n1007 ,\u2_Display/n1008 ,\u2_Display/n1009 ,\u2_Display/n1010 ,\u2_Display/n1011 }),
    .i1(32'b11111111111111111000001011111111),
    .i2(1'b1),
    .o(\u2_Display/n1014 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add36  (
    .i0({\u2_Display/n1015 ,\u2_Display/n1016 ,\u2_Display/n1017 ,\u2_Display/n1018 ,\u2_Display/n1019 ,\u2_Display/n1020 ,\u2_Display/n1021 ,\u2_Display/n1022 ,\u2_Display/n1023 ,\u2_Display/n1024 ,\u2_Display/n1025 ,\u2_Display/n1026 ,\u2_Display/n1027 ,\u2_Display/n1028 ,\u2_Display/n1029 ,\u2_Display/n1030 ,\u2_Display/n1031 ,\u2_Display/n1032 ,\u2_Display/n1033 ,\u2_Display/n1034 ,\u2_Display/n1035 ,\u2_Display/n1036 ,\u2_Display/n1037 ,\u2_Display/n1038 ,\u2_Display/n1039 ,\u2_Display/n1040 ,\u2_Display/n1041 ,\u2_Display/n1042 ,\u2_Display/n1043 ,\u2_Display/n1044 ,\u2_Display/n1045 ,\u2_Display/n1046 }),
    .i1(32'b11111111111111111100000101111111),
    .i2(1'b1),
    .o(\u2_Display/n1049 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add37  (
    .i0({\u2_Display/n1050 ,\u2_Display/n1051 ,\u2_Display/n1052 ,\u2_Display/n1053 ,\u2_Display/n1054 ,\u2_Display/n1055 ,\u2_Display/n1056 ,\u2_Display/n1057 ,\u2_Display/n1058 ,\u2_Display/n1059 ,\u2_Display/n1060 ,\u2_Display/n1061 ,\u2_Display/n1062 ,\u2_Display/n1063 ,\u2_Display/n1064 ,\u2_Display/n1065 ,\u2_Display/n1066 ,\u2_Display/n1067 ,\u2_Display/n1068 ,\u2_Display/n1069 ,\u2_Display/n1070 ,\u2_Display/n1071 ,\u2_Display/n1072 ,\u2_Display/n1073 ,\u2_Display/n1074 ,\u2_Display/n1075 ,\u2_Display/n1076 ,\u2_Display/n1077 ,\u2_Display/n1078 ,\u2_Display/n1079 ,\u2_Display/n1080 ,\u2_Display/n1081 }),
    .i1(32'b11111111111111111110000010111111),
    .i2(1'b1),
    .o(\u2_Display/n1084 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add38  (
    .i0({\u2_Display/n1085 ,\u2_Display/n1086 ,\u2_Display/n1087 ,\u2_Display/n1088 ,\u2_Display/n1089 ,\u2_Display/n1090 ,\u2_Display/n1091 ,\u2_Display/n1092 ,\u2_Display/n1093 ,\u2_Display/n1094 ,\u2_Display/n1095 ,\u2_Display/n1096 ,\u2_Display/n1097 ,\u2_Display/n1098 ,\u2_Display/n1099 ,\u2_Display/n1100 ,\u2_Display/n1101 ,\u2_Display/n1102 ,\u2_Display/n1103 ,\u2_Display/n1104 ,\u2_Display/n1105 ,\u2_Display/n1106 ,\u2_Display/n1107 ,\u2_Display/n1108 ,\u2_Display/n1109 ,\u2_Display/n1110 ,\u2_Display/n1111 ,\u2_Display/n1112 ,\u2_Display/n1113 ,\u2_Display/n1114 ,\u2_Display/n1115 ,\u2_Display/n1116 }),
    .i1(32'b11111111111111111111000001011111),
    .i2(1'b1),
    .o(\u2_Display/n1119 ));  // source/rtl/Display.v(230)
  add_pu32_pu32_pu1_o32 \u2_Display/add39  (
    .i0({\u2_Display/n1120 ,\u2_Display/n1121 ,\u2_Display/n1122 ,\u2_Display/n1123 ,\u2_Display/n1124 ,\u2_Display/n1125 ,\u2_Display/n1126 ,\u2_Display/n1127 ,\u2_Display/n1128 ,\u2_Display/n1129 ,\u2_Display/n1130 ,\u2_Display/n1131 ,\u2_Display/n1132 ,\u2_Display/n1133 ,\u2_Display/n1134 ,\u2_Display/n1135 ,\u2_Display/n1136 ,\u2_Display/n1137 ,\u2_Display/n1138 ,\u2_Display/n1139 ,\u2_Display/n1140 ,\u2_Display/n1141 ,\u2_Display/n1142 ,\u2_Display/n1143 ,\u2_Display/n1144 ,\u2_Display/n1145 ,\u2_Display/n1146 ,\u2_Display/n1147 ,\u2_Display/n1148 ,\u2_Display/n1149 ,\u2_Display/n1150 ,\u2_Display/n1151 }),
    .i1(32'b11111111111111111111100000101111),
    .i2(1'b1),
    .o(\u2_Display/n1154 ));  // source/rtl/Display.v(230)
  add_pu10_pu10_pu1_o10 \u2_Display/add40  (
    .i0({\u2_Display/n1177 ,\u2_Display/n1178 ,\u2_Display/n1179 ,\u2_Display/n1180 ,\u2_Display/n1181 ,\u2_Display/n1182 ,\u2_Display/n1183 ,\u2_Display/n1184 ,\u2_Display/n1185 ,\u2_Display/n1186 }),
    .i1(10'b0000010111),
    .i2(1'b1),
    .o(\u2_Display/n1189 [9:0]));  // source/rtl/Display.v(230)
  add_pu4_pu4_o5 \u2_Display/add4_2  (
    .i0(4'b0101),
    .i1(\u2_Display/i [10:7]),
    .o({\u2_Display/add4_2_co ,\u2_Display/n94 [3:0]}));  // source/rtl/Display.v(181)
  add_pu32_pu32_pu1_o32 \u2_Display/add51  (
    .i0(\u2_Display/counta ),
    .i1(32'b00011110111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n1542 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add52  (
    .i0({\u2_Display/n1543 ,\u2_Display/n1544 ,\u2_Display/n1545 ,\u2_Display/n1546 ,\u2_Display/n1547 ,\u2_Display/n1548 ,\u2_Display/n1549 ,\u2_Display/n1550 ,\u2_Display/n1551 ,\u2_Display/n1552 ,\u2_Display/n1553 ,\u2_Display/n1554 ,\u2_Display/n1555 ,\u2_Display/n1556 ,\u2_Display/n1557 ,\u2_Display/n1558 ,\u2_Display/n1559 ,\u2_Display/n1560 ,\u2_Display/n1561 ,\u2_Display/n1562 ,\u2_Display/n1563 ,\u2_Display/n1564 ,\u2_Display/n1565 ,\u2_Display/n1566 ,\u2_Display/n1567 ,\u2_Display/n1568 ,\u2_Display/n1569 ,\u2_Display/n1570 ,\u2_Display/n1571 ,\u2_Display/n1572 ,\u2_Display/n1573 ,\u2_Display/n1574 }),
    .i1(32'b10001111011111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n1577 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add53  (
    .i0({\u2_Display/n1578 ,\u2_Display/n1579 ,\u2_Display/n1580 ,\u2_Display/n1581 ,\u2_Display/n1582 ,\u2_Display/n1583 ,\u2_Display/n1584 ,\u2_Display/n1585 ,\u2_Display/n1586 ,\u2_Display/n1587 ,\u2_Display/n1588 ,\u2_Display/n1589 ,\u2_Display/n1590 ,\u2_Display/n1591 ,\u2_Display/n1592 ,\u2_Display/n1593 ,\u2_Display/n1594 ,\u2_Display/n1595 ,\u2_Display/n1596 ,\u2_Display/n1597 ,\u2_Display/n1598 ,\u2_Display/n1599 ,\u2_Display/n1600 ,\u2_Display/n1601 ,\u2_Display/n1602 ,\u2_Display/n1603 ,\u2_Display/n1604 ,\u2_Display/n1605 ,\u2_Display/n1606 ,\u2_Display/n1607 ,\u2_Display/n1608 ,\u2_Display/n1609 }),
    .i1(32'b11000111101111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n1612 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add54  (
    .i0({\u2_Display/n1613 ,\u2_Display/n1614 ,\u2_Display/n1615 ,\u2_Display/n1616 ,\u2_Display/n1617 ,\u2_Display/n1618 ,\u2_Display/n1619 ,\u2_Display/n1620 ,\u2_Display/n1621 ,\u2_Display/n1622 ,\u2_Display/n1623 ,\u2_Display/n1624 ,\u2_Display/n1625 ,\u2_Display/n1626 ,\u2_Display/n1627 ,\u2_Display/n1628 ,\u2_Display/n1629 ,\u2_Display/n1630 ,\u2_Display/n1631 ,\u2_Display/n1632 ,\u2_Display/n1633 ,\u2_Display/n1634 ,\u2_Display/n1635 ,\u2_Display/n1636 ,\u2_Display/n1637 ,\u2_Display/n1638 ,\u2_Display/n1639 ,\u2_Display/n1640 ,\u2_Display/n1641 ,\u2_Display/n1642 ,\u2_Display/n1643 ,\u2_Display/n1644 }),
    .i1(32'b11100011110111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n1647 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add55  (
    .i0({\u2_Display/n1648 ,\u2_Display/n1649 ,\u2_Display/n1650 ,\u2_Display/n1651 ,\u2_Display/n1652 ,\u2_Display/n1653 ,\u2_Display/n1654 ,\u2_Display/n1655 ,\u2_Display/n1656 ,\u2_Display/n1657 ,\u2_Display/n1658 ,\u2_Display/n1659 ,\u2_Display/n1660 ,\u2_Display/n1661 ,\u2_Display/n1662 ,\u2_Display/n1663 ,\u2_Display/n1664 ,\u2_Display/n1665 ,\u2_Display/n1666 ,\u2_Display/n1667 ,\u2_Display/n1668 ,\u2_Display/n1669 ,\u2_Display/n1670 ,\u2_Display/n1671 ,\u2_Display/n1672 ,\u2_Display/n1673 ,\u2_Display/n1674 ,\u2_Display/n1675 ,\u2_Display/n1676 ,\u2_Display/n1677 ,\u2_Display/n1678 ,\u2_Display/n1679 }),
    .i1(32'b11110001111011111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n1682 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add56  (
    .i0({\u2_Display/n1683 ,\u2_Display/n1684 ,\u2_Display/n1685 ,\u2_Display/n1686 ,\u2_Display/n1687 ,\u2_Display/n1688 ,\u2_Display/n1689 ,\u2_Display/n1690 ,\u2_Display/n1691 ,\u2_Display/n1692 ,\u2_Display/n1693 ,\u2_Display/n1694 ,\u2_Display/n1695 ,\u2_Display/n1696 ,\u2_Display/n1697 ,\u2_Display/n1698 ,\u2_Display/n1699 ,\u2_Display/n1700 ,\u2_Display/n1701 ,\u2_Display/n1702 ,\u2_Display/n1703 ,\u2_Display/n1704 ,\u2_Display/n1705 ,\u2_Display/n1706 ,\u2_Display/n1707 ,\u2_Display/n1708 ,\u2_Display/n1709 ,\u2_Display/n1710 ,\u2_Display/n1711 ,\u2_Display/n1712 ,\u2_Display/n1713 ,\u2_Display/n1714 }),
    .i1(32'b11111000111101111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n1717 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add57  (
    .i0({\u2_Display/n1718 ,\u2_Display/n1719 ,\u2_Display/n1720 ,\u2_Display/n1721 ,\u2_Display/n1722 ,\u2_Display/n1723 ,\u2_Display/n1724 ,\u2_Display/n1725 ,\u2_Display/n1726 ,\u2_Display/n1727 ,\u2_Display/n1728 ,\u2_Display/n1729 ,\u2_Display/n1730 ,\u2_Display/n1731 ,\u2_Display/n1732 ,\u2_Display/n1733 ,\u2_Display/n1734 ,\u2_Display/n1735 ,\u2_Display/n1736 ,\u2_Display/n1737 ,\u2_Display/n1738 ,\u2_Display/n1739 ,\u2_Display/n1740 ,\u2_Display/n1741 ,\u2_Display/n1742 ,\u2_Display/n1743 ,\u2_Display/n1744 ,\u2_Display/n1745 ,\u2_Display/n1746 ,\u2_Display/n1747 ,\u2_Display/n1748 ,\u2_Display/n1749 }),
    .i1(32'b11111100011110111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n1752 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add58  (
    .i0({\u2_Display/n1753 ,\u2_Display/n1754 ,\u2_Display/n1755 ,\u2_Display/n1756 ,\u2_Display/n1757 ,\u2_Display/n1758 ,\u2_Display/n1759 ,\u2_Display/n1760 ,\u2_Display/n1761 ,\u2_Display/n1762 ,\u2_Display/n1763 ,\u2_Display/n1764 ,\u2_Display/n1765 ,\u2_Display/n1766 ,\u2_Display/n1767 ,\u2_Display/n1768 ,\u2_Display/n1769 ,\u2_Display/n1770 ,\u2_Display/n1771 ,\u2_Display/n1772 ,\u2_Display/n1773 ,\u2_Display/n1774 ,\u2_Display/n1775 ,\u2_Display/n1776 ,\u2_Display/n1777 ,\u2_Display/n1778 ,\u2_Display/n1779 ,\u2_Display/n1780 ,\u2_Display/n1781 ,\u2_Display/n1782 ,\u2_Display/n1783 ,\u2_Display/n1784 }),
    .i1(32'b11111110001111011111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n1787 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add59  (
    .i0({\u2_Display/n1788 ,\u2_Display/n1789 ,\u2_Display/n1790 ,\u2_Display/n1791 ,\u2_Display/n1792 ,\u2_Display/n1793 ,\u2_Display/n1794 ,\u2_Display/n1795 ,\u2_Display/n1796 ,\u2_Display/n1797 ,\u2_Display/n1798 ,\u2_Display/n1799 ,\u2_Display/n1800 ,\u2_Display/n1801 ,\u2_Display/n1802 ,\u2_Display/n1803 ,\u2_Display/n1804 ,\u2_Display/n1805 ,\u2_Display/n1806 ,\u2_Display/n1807 ,\u2_Display/n1808 ,\u2_Display/n1809 ,\u2_Display/n1810 ,\u2_Display/n1811 ,\u2_Display/n1812 ,\u2_Display/n1813 ,\u2_Display/n1814 ,\u2_Display/n1815 ,\u2_Display/n1816 ,\u2_Display/n1817 ,\u2_Display/n1818 ,\u2_Display/n1819 }),
    .i1(32'b11111111000111101111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n1822 ));  // source/rtl/Display.v(213)
  add_pu1_pu1_o2 \u2_Display/add5_2  (
    .i0(1'b1),
    .i1(\u2_Display/j [9]),
    .o({\u2_Display/add5_2_co ,\u2_Display/n99 [0]}));  // source/rtl/Display.v(181)
  add_pu32_pu32_pu1_o32 \u2_Display/add60  (
    .i0({\u2_Display/n1823 ,\u2_Display/n1824 ,\u2_Display/n1825 ,\u2_Display/n1826 ,\u2_Display/n1827 ,\u2_Display/n1828 ,\u2_Display/n1829 ,\u2_Display/n1830 ,\u2_Display/n1831 ,\u2_Display/n1832 ,\u2_Display/n1833 ,\u2_Display/n1834 ,\u2_Display/n1835 ,\u2_Display/n1836 ,\u2_Display/n1837 ,\u2_Display/n1838 ,\u2_Display/n1839 ,\u2_Display/n1840 ,\u2_Display/n1841 ,\u2_Display/n1842 ,\u2_Display/n1843 ,\u2_Display/n1844 ,\u2_Display/n1845 ,\u2_Display/n1846 ,\u2_Display/n1847 ,\u2_Display/n1848 ,\u2_Display/n1849 ,\u2_Display/n1850 ,\u2_Display/n1851 ,\u2_Display/n1852 ,\u2_Display/n1853 ,\u2_Display/n1854 }),
    .i1(32'b11111111100011110111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n1857 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add61  (
    .i0({\u2_Display/n1858 ,\u2_Display/n1859 ,\u2_Display/n1860 ,\u2_Display/n1861 ,\u2_Display/n1862 ,\u2_Display/n1863 ,\u2_Display/n1864 ,\u2_Display/n1865 ,\u2_Display/n1866 ,\u2_Display/n1867 ,\u2_Display/n1868 ,\u2_Display/n1869 ,\u2_Display/n1870 ,\u2_Display/n1871 ,\u2_Display/n1872 ,\u2_Display/n1873 ,\u2_Display/n1874 ,\u2_Display/n1875 ,\u2_Display/n1876 ,\u2_Display/n1877 ,\u2_Display/n1878 ,\u2_Display/n1879 ,\u2_Display/n1880 ,\u2_Display/n1881 ,\u2_Display/n1882 ,\u2_Display/n1883 ,\u2_Display/n1884 ,\u2_Display/n1885 ,\u2_Display/n1886 ,\u2_Display/n1887 ,\u2_Display/n1888 ,\u2_Display/n1889 }),
    .i1(32'b11111111110001111011111111111111),
    .i2(1'b1),
    .o(\u2_Display/n1892 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add62  (
    .i0({\u2_Display/n1893 ,\u2_Display/n1894 ,\u2_Display/n1895 ,\u2_Display/n1896 ,\u2_Display/n1897 ,\u2_Display/n1898 ,\u2_Display/n1899 ,\u2_Display/n1900 ,\u2_Display/n1901 ,\u2_Display/n1902 ,\u2_Display/n1903 ,\u2_Display/n1904 ,\u2_Display/n1905 ,\u2_Display/n1906 ,\u2_Display/n1907 ,\u2_Display/n1908 ,\u2_Display/n1909 ,\u2_Display/n1910 ,\u2_Display/n1911 ,\u2_Display/n1912 ,\u2_Display/n1913 ,\u2_Display/n1914 ,\u2_Display/n1915 ,\u2_Display/n1916 ,\u2_Display/n1917 ,\u2_Display/n1918 ,\u2_Display/n1919 ,\u2_Display/n1920 ,\u2_Display/n1921 ,\u2_Display/n1922 ,\u2_Display/n1923 ,\u2_Display/n1924 }),
    .i1(32'b11111111111000111101111111111111),
    .i2(1'b1),
    .o(\u2_Display/n1927 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add63  (
    .i0({\u2_Display/n1928 ,\u2_Display/n1929 ,\u2_Display/n1930 ,\u2_Display/n1931 ,\u2_Display/n1932 ,\u2_Display/n1933 ,\u2_Display/n1934 ,\u2_Display/n1935 ,\u2_Display/n1936 ,\u2_Display/n1937 ,\u2_Display/n1938 ,\u2_Display/n1939 ,\u2_Display/n1940 ,\u2_Display/n1941 ,\u2_Display/n1942 ,\u2_Display/n1943 ,\u2_Display/n1944 ,\u2_Display/n1945 ,\u2_Display/n1946 ,\u2_Display/n1947 ,\u2_Display/n1948 ,\u2_Display/n1949 ,\u2_Display/n1950 ,\u2_Display/n1951 ,\u2_Display/n1952 ,\u2_Display/n1953 ,\u2_Display/n1954 ,\u2_Display/n1955 ,\u2_Display/n1956 ,\u2_Display/n1957 ,\u2_Display/n1958 ,\u2_Display/n1959 }),
    .i1(32'b11111111111100011110111111111111),
    .i2(1'b1),
    .o(\u2_Display/n1962 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add64  (
    .i0({\u2_Display/n1963 ,\u2_Display/n1964 ,\u2_Display/n1965 ,\u2_Display/n1966 ,\u2_Display/n1967 ,\u2_Display/n1968 ,\u2_Display/n1969 ,\u2_Display/n1970 ,\u2_Display/n1971 ,\u2_Display/n1972 ,\u2_Display/n1973 ,\u2_Display/n1974 ,\u2_Display/n1975 ,\u2_Display/n1976 ,\u2_Display/n1977 ,\u2_Display/n1978 ,\u2_Display/n1979 ,\u2_Display/n1980 ,\u2_Display/n1981 ,\u2_Display/n1982 ,\u2_Display/n1983 ,\u2_Display/n1984 ,\u2_Display/n1985 ,\u2_Display/n1986 ,\u2_Display/n1987 ,\u2_Display/n1988 ,\u2_Display/n1989 ,\u2_Display/n1990 ,\u2_Display/n1991 ,\u2_Display/n1992 ,\u2_Display/n1993 ,\u2_Display/n1994 }),
    .i1(32'b11111111111110001111011111111111),
    .i2(1'b1),
    .o(\u2_Display/n1997 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add65  (
    .i0({\u2_Display/n1998 ,\u2_Display/n1999 ,\u2_Display/n2000 ,\u2_Display/n2001 ,\u2_Display/n2002 ,\u2_Display/n2003 ,\u2_Display/n2004 ,\u2_Display/n2005 ,\u2_Display/n2006 ,\u2_Display/n2007 ,\u2_Display/n2008 ,\u2_Display/n2009 ,\u2_Display/n2010 ,\u2_Display/n2011 ,\u2_Display/n2012 ,\u2_Display/n2013 ,\u2_Display/n2014 ,\u2_Display/n2015 ,\u2_Display/n2016 ,\u2_Display/n2017 ,\u2_Display/n2018 ,\u2_Display/n2019 ,\u2_Display/n2020 ,\u2_Display/n2021 ,\u2_Display/n2022 ,\u2_Display/n2023 ,\u2_Display/n2024 ,\u2_Display/n2025 ,\u2_Display/n2026 ,\u2_Display/n2027 ,\u2_Display/n2028 ,\u2_Display/n2029 }),
    .i1(32'b11111111111111000111101111111111),
    .i2(1'b1),
    .o(\u2_Display/n2032 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add66  (
    .i0({\u2_Display/n2033 ,\u2_Display/n2034 ,\u2_Display/n2035 ,\u2_Display/n2036 ,\u2_Display/n2037 ,\u2_Display/n2038 ,\u2_Display/n2039 ,\u2_Display/n2040 ,\u2_Display/n2041 ,\u2_Display/n2042 ,\u2_Display/n2043 ,\u2_Display/n2044 ,\u2_Display/n2045 ,\u2_Display/n2046 ,\u2_Display/n2047 ,\u2_Display/n2048 ,\u2_Display/n2049 ,\u2_Display/n2050 ,\u2_Display/n2051 ,\u2_Display/n2052 ,\u2_Display/n2053 ,\u2_Display/n2054 ,\u2_Display/n2055 ,\u2_Display/n2056 ,\u2_Display/n2057 ,\u2_Display/n2058 ,\u2_Display/n2059 ,\u2_Display/n2060 ,\u2_Display/n2061 ,\u2_Display/n2062 ,\u2_Display/n2063 ,\u2_Display/n2064 }),
    .i1(32'b11111111111111100011110111111111),
    .i2(1'b1),
    .o(\u2_Display/n2067 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add67  (
    .i0({\u2_Display/n2068 ,\u2_Display/n2069 ,\u2_Display/n2070 ,\u2_Display/n2071 ,\u2_Display/n2072 ,\u2_Display/n2073 ,\u2_Display/n2074 ,\u2_Display/n2075 ,\u2_Display/n2076 ,\u2_Display/n2077 ,\u2_Display/n2078 ,\u2_Display/n2079 ,\u2_Display/n2080 ,\u2_Display/n2081 ,\u2_Display/n2082 ,\u2_Display/n2083 ,\u2_Display/n2084 ,\u2_Display/n2085 ,\u2_Display/n2086 ,\u2_Display/n2087 ,\u2_Display/n2088 ,\u2_Display/n2089 ,\u2_Display/n2090 ,\u2_Display/n2091 ,\u2_Display/n2092 ,\u2_Display/n2093 ,\u2_Display/n2094 ,\u2_Display/n2095 ,\u2_Display/n2096 ,\u2_Display/n2097 ,\u2_Display/n2098 ,\u2_Display/n2099 }),
    .i1(32'b11111111111111110001111011111111),
    .i2(1'b1),
    .o(\u2_Display/n2102 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add68  (
    .i0({\u2_Display/n2103 ,\u2_Display/n2104 ,\u2_Display/n2105 ,\u2_Display/n2106 ,\u2_Display/n2107 ,\u2_Display/n2108 ,\u2_Display/n2109 ,\u2_Display/n2110 ,\u2_Display/n2111 ,\u2_Display/n2112 ,\u2_Display/n2113 ,\u2_Display/n2114 ,\u2_Display/n2115 ,\u2_Display/n2116 ,\u2_Display/n2117 ,\u2_Display/n2118 ,\u2_Display/n2119 ,\u2_Display/n2120 ,\u2_Display/n2121 ,\u2_Display/n2122 ,\u2_Display/n2123 ,\u2_Display/n2124 ,\u2_Display/n2125 ,\u2_Display/n2126 ,\u2_Display/n2127 ,\u2_Display/n2128 ,\u2_Display/n2129 ,\u2_Display/n2130 ,\u2_Display/n2131 ,\u2_Display/n2132 ,\u2_Display/n2133 ,\u2_Display/n2134 }),
    .i1(32'b11111111111111111000111101111111),
    .i2(1'b1),
    .o(\u2_Display/n2137 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add69  (
    .i0({\u2_Display/n2138 ,\u2_Display/n2139 ,\u2_Display/n2140 ,\u2_Display/n2141 ,\u2_Display/n2142 ,\u2_Display/n2143 ,\u2_Display/n2144 ,\u2_Display/n2145 ,\u2_Display/n2146 ,\u2_Display/n2147 ,\u2_Display/n2148 ,\u2_Display/n2149 ,\u2_Display/n2150 ,\u2_Display/n2151 ,\u2_Display/n2152 ,\u2_Display/n2153 ,\u2_Display/n2154 ,\u2_Display/n2155 ,\u2_Display/n2156 ,\u2_Display/n2157 ,\u2_Display/n2158 ,\u2_Display/n2159 ,\u2_Display/n2160 ,\u2_Display/n2161 ,\u2_Display/n2162 ,\u2_Display/n2163 ,\u2_Display/n2164 ,\u2_Display/n2165 ,\u2_Display/n2166 ,\u2_Display/n2167 ,\u2_Display/n2168 ,\u2_Display/n2169 }),
    .i1(32'b11111111111111111100011110111111),
    .i2(1'b1),
    .o(\u2_Display/n2172 ));  // source/rtl/Display.v(213)
  add_pu3_pu3_o4 \u2_Display/add6_2  (
    .i0(3'b101),
    .i1(\u2_Display/j [9:7]),
    .o({\u2_Display/add6_2_co ,\u2_Display/n135 [2:0]}));  // source/rtl/Display.v(197)
  add_pu32_pu32_pu1_o32 \u2_Display/add70  (
    .i0({\u2_Display/n2173 ,\u2_Display/n2174 ,\u2_Display/n2175 ,\u2_Display/n2176 ,\u2_Display/n2177 ,\u2_Display/n2178 ,\u2_Display/n2179 ,\u2_Display/n2180 ,\u2_Display/n2181 ,\u2_Display/n2182 ,\u2_Display/n2183 ,\u2_Display/n2184 ,\u2_Display/n2185 ,\u2_Display/n2186 ,\u2_Display/n2187 ,\u2_Display/n2188 ,\u2_Display/n2189 ,\u2_Display/n2190 ,\u2_Display/n2191 ,\u2_Display/n2192 ,\u2_Display/n2193 ,\u2_Display/n2194 ,\u2_Display/n2195 ,\u2_Display/n2196 ,\u2_Display/n2197 ,\u2_Display/n2198 ,\u2_Display/n2199 ,\u2_Display/n2200 ,\u2_Display/n2201 ,\u2_Display/n2202 ,\u2_Display/n2203 ,\u2_Display/n2204 }),
    .i1(32'b11111111111111111110001111011111),
    .i2(1'b1),
    .o(\u2_Display/n2207 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add71  (
    .i0({\u2_Display/n2208 ,\u2_Display/n2209 ,\u2_Display/n2210 ,\u2_Display/n2211 ,\u2_Display/n2212 ,\u2_Display/n2213 ,\u2_Display/n2214 ,\u2_Display/n2215 ,\u2_Display/n2216 ,\u2_Display/n2217 ,\u2_Display/n2218 ,\u2_Display/n2219 ,\u2_Display/n2220 ,\u2_Display/n2221 ,\u2_Display/n2222 ,\u2_Display/n2223 ,\u2_Display/n2224 ,\u2_Display/n2225 ,\u2_Display/n2226 ,\u2_Display/n2227 ,\u2_Display/n2228 ,\u2_Display/n2229 ,\u2_Display/n2230 ,\u2_Display/n2231 ,\u2_Display/n2232 ,\u2_Display/n2233 ,\u2_Display/n2234 ,\u2_Display/n2235 ,\u2_Display/n2236 ,\u2_Display/n2237 ,\u2_Display/n2238 ,\u2_Display/n2239 }),
    .i1(32'b11111111111111111111000111101111),
    .i2(1'b1),
    .o(\u2_Display/n2242 ));  // source/rtl/Display.v(213)
  add_pu32_pu32_pu1_o32 \u2_Display/add72  (
    .i0({\u2_Display/n2243 ,\u2_Display/n2244 ,\u2_Display/n2245 ,\u2_Display/n2246 ,\u2_Display/n2247 ,\u2_Display/n2248 ,\u2_Display/n2249 ,\u2_Display/n2250 ,\u2_Display/n2251 ,\u2_Display/n2252 ,\u2_Display/n2253 ,\u2_Display/n2254 ,\u2_Display/n2255 ,\u2_Display/n2256 ,\u2_Display/n2257 ,\u2_Display/n2258 ,\u2_Display/n2259 ,\u2_Display/n2260 ,\u2_Display/n2261 ,\u2_Display/n2262 ,\u2_Display/n2263 ,\u2_Display/n2264 ,\u2_Display/n2265 ,\u2_Display/n2266 ,\u2_Display/n2267 ,\u2_Display/n2268 ,\u2_Display/n2269 ,\u2_Display/n2270 ,\u2_Display/n2271 ,\u2_Display/n2272 ,\u2_Display/n2273 ,\u2_Display/n2274 }),
    .i1(32'b11111111111111111111100011110111),
    .i2(1'b1),
    .o(\u2_Display/n2277 ));  // source/rtl/Display.v(213)
  add_pu10_pu10_pu1_o10 \u2_Display/add73  (
    .i0({\u2_Display/n2300 ,\u2_Display/n2301 ,\u2_Display/n2302 ,\u2_Display/n2303 ,\u2_Display/n2304 ,\u2_Display/n2305 ,\u2_Display/n2306 ,\u2_Display/n2307 ,\u2_Display/n2308 ,\u2_Display/n2309 }),
    .i1(10'b0001111011),
    .i2(1'b1),
    .o(\u2_Display/n2312 [9:0]));  // source/rtl/Display.v(213)
  add_pu2_pu2_o3 \u2_Display/add7_2  (
    .i0(2'b01),
    .i1(\u2_Display/i [10:9]),
    .o({\u2_Display/add7_2_co ,\u2_Display/n140 [1:0]}));  // source/rtl/Display.v(197)
  add_pu32_pu32_pu1_o32 \u2_Display/add84  (
    .i0(\u2_Display/counta ),
    .i1(32'b01101001111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n2665 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add85  (
    .i0({\u2_Display/n2666 ,\u2_Display/n2667 ,\u2_Display/n2668 ,\u2_Display/n2669 ,\u2_Display/n2670 ,\u2_Display/n2671 ,\u2_Display/n2672 ,\u2_Display/n2673 ,\u2_Display/n2674 ,\u2_Display/n2675 ,\u2_Display/n2676 ,\u2_Display/n2677 ,\u2_Display/n2678 ,\u2_Display/n2679 ,\u2_Display/n2680 ,\u2_Display/n2681 ,\u2_Display/n2682 ,\u2_Display/n2683 ,\u2_Display/n2684 ,\u2_Display/n2685 ,\u2_Display/n2686 ,\u2_Display/n2687 ,\u2_Display/n2688 ,\u2_Display/n2689 ,\u2_Display/n2690 ,\u2_Display/n2691 ,\u2_Display/n2692 ,\u2_Display/n2693 ,\u2_Display/n2694 ,\u2_Display/n2695 ,\u2_Display/n2696 ,\u2_Display/n2697 }),
    .i1(32'b10110100111111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n2700 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add86  (
    .i0({\u2_Display/n2701 ,\u2_Display/n2702 ,\u2_Display/n2703 ,\u2_Display/n2704 ,\u2_Display/n2705 ,\u2_Display/n2706 ,\u2_Display/n2707 ,\u2_Display/n2708 ,\u2_Display/n2709 ,\u2_Display/n2710 ,\u2_Display/n2711 ,\u2_Display/n2712 ,\u2_Display/n2713 ,\u2_Display/n2714 ,\u2_Display/n2715 ,\u2_Display/n2716 ,\u2_Display/n2717 ,\u2_Display/n2718 ,\u2_Display/n2719 ,\u2_Display/n2720 ,\u2_Display/n2721 ,\u2_Display/n2722 ,\u2_Display/n2723 ,\u2_Display/n2724 ,\u2_Display/n2725 ,\u2_Display/n2726 ,\u2_Display/n2727 ,\u2_Display/n2728 ,\u2_Display/n2729 ,\u2_Display/n2730 ,\u2_Display/n2731 ,\u2_Display/n2732 }),
    .i1(32'b11011010011111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n2735 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add87  (
    .i0({\u2_Display/n2736 ,\u2_Display/n2737 ,\u2_Display/n2738 ,\u2_Display/n2739 ,\u2_Display/n2740 ,\u2_Display/n2741 ,\u2_Display/n2742 ,\u2_Display/n2743 ,\u2_Display/n2744 ,\u2_Display/n2745 ,\u2_Display/n2746 ,\u2_Display/n2747 ,\u2_Display/n2748 ,\u2_Display/n2749 ,\u2_Display/n2750 ,\u2_Display/n2751 ,\u2_Display/n2752 ,\u2_Display/n2753 ,\u2_Display/n2754 ,\u2_Display/n2755 ,\u2_Display/n2756 ,\u2_Display/n2757 ,\u2_Display/n2758 ,\u2_Display/n2759 ,\u2_Display/n2760 ,\u2_Display/n2761 ,\u2_Display/n2762 ,\u2_Display/n2763 ,\u2_Display/n2764 ,\u2_Display/n2765 ,\u2_Display/n2766 ,\u2_Display/n2767 }),
    .i1(32'b11101101001111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n2770 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add88  (
    .i0({\u2_Display/n2771 ,\u2_Display/n2772 ,\u2_Display/n2773 ,\u2_Display/n2774 ,\u2_Display/n2775 ,\u2_Display/n2776 ,\u2_Display/n2777 ,\u2_Display/n2778 ,\u2_Display/n2779 ,\u2_Display/n2780 ,\u2_Display/n2781 ,\u2_Display/n2782 ,\u2_Display/n2783 ,\u2_Display/n2784 ,\u2_Display/n2785 ,\u2_Display/n2786 ,\u2_Display/n2787 ,\u2_Display/n2788 ,\u2_Display/n2789 ,\u2_Display/n2790 ,\u2_Display/n2791 ,\u2_Display/n2792 ,\u2_Display/n2793 ,\u2_Display/n2794 ,\u2_Display/n2795 ,\u2_Display/n2796 ,\u2_Display/n2797 ,\u2_Display/n2798 ,\u2_Display/n2799 ,\u2_Display/n2800 ,\u2_Display/n2801 ,\u2_Display/n2802 }),
    .i1(32'b11110110100111111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n2805 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add89  (
    .i0({\u2_Display/n2806 ,\u2_Display/n2807 ,\u2_Display/n2808 ,\u2_Display/n2809 ,\u2_Display/n2810 ,\u2_Display/n2811 ,\u2_Display/n2812 ,\u2_Display/n2813 ,\u2_Display/n2814 ,\u2_Display/n2815 ,\u2_Display/n2816 ,\u2_Display/n2817 ,\u2_Display/n2818 ,\u2_Display/n2819 ,\u2_Display/n2820 ,\u2_Display/n2821 ,\u2_Display/n2822 ,\u2_Display/n2823 ,\u2_Display/n2824 ,\u2_Display/n2825 ,\u2_Display/n2826 ,\u2_Display/n2827 ,\u2_Display/n2828 ,\u2_Display/n2829 ,\u2_Display/n2830 ,\u2_Display/n2831 ,\u2_Display/n2832 ,\u2_Display/n2833 ,\u2_Display/n2834 ,\u2_Display/n2835 ,\u2_Display/n2836 ,\u2_Display/n2837 }),
    .i1(32'b11111011010011111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n2840 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add90  (
    .i0({\u2_Display/n2841 ,\u2_Display/n2842 ,\u2_Display/n2843 ,\u2_Display/n2844 ,\u2_Display/n2845 ,\u2_Display/n2846 ,\u2_Display/n2847 ,\u2_Display/n2848 ,\u2_Display/n2849 ,\u2_Display/n2850 ,\u2_Display/n2851 ,\u2_Display/n2852 ,\u2_Display/n2853 ,\u2_Display/n2854 ,\u2_Display/n2855 ,\u2_Display/n2856 ,\u2_Display/n2857 ,\u2_Display/n2858 ,\u2_Display/n2859 ,\u2_Display/n2860 ,\u2_Display/n2861 ,\u2_Display/n2862 ,\u2_Display/n2863 ,\u2_Display/n2864 ,\u2_Display/n2865 ,\u2_Display/n2866 ,\u2_Display/n2867 ,\u2_Display/n2868 ,\u2_Display/n2869 ,\u2_Display/n2870 ,\u2_Display/n2871 ,\u2_Display/n2872 }),
    .i1(32'b11111101101001111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n2875 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add91  (
    .i0({\u2_Display/n2876 ,\u2_Display/n2877 ,\u2_Display/n2878 ,\u2_Display/n2879 ,\u2_Display/n2880 ,\u2_Display/n2881 ,\u2_Display/n2882 ,\u2_Display/n2883 ,\u2_Display/n2884 ,\u2_Display/n2885 ,\u2_Display/n2886 ,\u2_Display/n2887 ,\u2_Display/n2888 ,\u2_Display/n2889 ,\u2_Display/n2890 ,\u2_Display/n2891 ,\u2_Display/n2892 ,\u2_Display/n2893 ,\u2_Display/n2894 ,\u2_Display/n2895 ,\u2_Display/n2896 ,\u2_Display/n2897 ,\u2_Display/n2898 ,\u2_Display/n2899 ,\u2_Display/n2900 ,\u2_Display/n2901 ,\u2_Display/n2902 ,\u2_Display/n2903 ,\u2_Display/n2904 ,\u2_Display/n2905 ,\u2_Display/n2906 ,\u2_Display/n2907 }),
    .i1(32'b11111110110100111111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n2910 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add92  (
    .i0({\u2_Display/n2911 ,\u2_Display/n2912 ,\u2_Display/n2913 ,\u2_Display/n2914 ,\u2_Display/n2915 ,\u2_Display/n2916 ,\u2_Display/n2917 ,\u2_Display/n2918 ,\u2_Display/n2919 ,\u2_Display/n2920 ,\u2_Display/n2921 ,\u2_Display/n2922 ,\u2_Display/n2923 ,\u2_Display/n2924 ,\u2_Display/n2925 ,\u2_Display/n2926 ,\u2_Display/n2927 ,\u2_Display/n2928 ,\u2_Display/n2929 ,\u2_Display/n2930 ,\u2_Display/n2931 ,\u2_Display/n2932 ,\u2_Display/n2933 ,\u2_Display/n2934 ,\u2_Display/n2935 ,\u2_Display/n2936 ,\u2_Display/n2937 ,\u2_Display/n2938 ,\u2_Display/n2939 ,\u2_Display/n2940 ,\u2_Display/n2941 ,\u2_Display/n2942 }),
    .i1(32'b11111111011010011111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n2945 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add93  (
    .i0({\u2_Display/n2946 ,\u2_Display/n2947 ,\u2_Display/n2948 ,\u2_Display/n2949 ,\u2_Display/n2950 ,\u2_Display/n2951 ,\u2_Display/n2952 ,\u2_Display/n2953 ,\u2_Display/n2954 ,\u2_Display/n2955 ,\u2_Display/n2956 ,\u2_Display/n2957 ,\u2_Display/n2958 ,\u2_Display/n2959 ,\u2_Display/n2960 ,\u2_Display/n2961 ,\u2_Display/n2962 ,\u2_Display/n2963 ,\u2_Display/n2964 ,\u2_Display/n2965 ,\u2_Display/n2966 ,\u2_Display/n2967 ,\u2_Display/n2968 ,\u2_Display/n2969 ,\u2_Display/n2970 ,\u2_Display/n2971 ,\u2_Display/n2972 ,\u2_Display/n2973 ,\u2_Display/n2974 ,\u2_Display/n2975 ,\u2_Display/n2976 ,\u2_Display/n2977 }),
    .i1(32'b11111111101101001111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n2980 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add94  (
    .i0({\u2_Display/n2981 ,\u2_Display/n2982 ,\u2_Display/n2983 ,\u2_Display/n2984 ,\u2_Display/n2985 ,\u2_Display/n2986 ,\u2_Display/n2987 ,\u2_Display/n2988 ,\u2_Display/n2989 ,\u2_Display/n2990 ,\u2_Display/n2991 ,\u2_Display/n2992 ,\u2_Display/n2993 ,\u2_Display/n2994 ,\u2_Display/n2995 ,\u2_Display/n2996 ,\u2_Display/n2997 ,\u2_Display/n2998 ,\u2_Display/n2999 ,\u2_Display/n3000 ,\u2_Display/n3001 ,\u2_Display/n3002 ,\u2_Display/n3003 ,\u2_Display/n3004 ,\u2_Display/n3005 ,\u2_Display/n3006 ,\u2_Display/n3007 ,\u2_Display/n3008 ,\u2_Display/n3009 ,\u2_Display/n3010 ,\u2_Display/n3011 ,\u2_Display/n3012 }),
    .i1(32'b11111111110110100111111111111111),
    .i2(1'b1),
    .o(\u2_Display/n3015 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add95  (
    .i0({\u2_Display/n3016 ,\u2_Display/n3017 ,\u2_Display/n3018 ,\u2_Display/n3019 ,\u2_Display/n3020 ,\u2_Display/n3021 ,\u2_Display/n3022 ,\u2_Display/n3023 ,\u2_Display/n3024 ,\u2_Display/n3025 ,\u2_Display/n3026 ,\u2_Display/n3027 ,\u2_Display/n3028 ,\u2_Display/n3029 ,\u2_Display/n3030 ,\u2_Display/n3031 ,\u2_Display/n3032 ,\u2_Display/n3033 ,\u2_Display/n3034 ,\u2_Display/n3035 ,\u2_Display/n3036 ,\u2_Display/n3037 ,\u2_Display/n3038 ,\u2_Display/n3039 ,\u2_Display/n3040 ,\u2_Display/n3041 ,\u2_Display/n3042 ,\u2_Display/n3043 ,\u2_Display/n3044 ,\u2_Display/n3045 ,\u2_Display/n3046 ,\u2_Display/n3047 }),
    .i1(32'b11111111111011010011111111111111),
    .i2(1'b1),
    .o(\u2_Display/n3050 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add96  (
    .i0({\u2_Display/n3051 ,\u2_Display/n3052 ,\u2_Display/n3053 ,\u2_Display/n3054 ,\u2_Display/n3055 ,\u2_Display/n3056 ,\u2_Display/n3057 ,\u2_Display/n3058 ,\u2_Display/n3059 ,\u2_Display/n3060 ,\u2_Display/n3061 ,\u2_Display/n3062 ,\u2_Display/n3063 ,\u2_Display/n3064 ,\u2_Display/n3065 ,\u2_Display/n3066 ,\u2_Display/n3067 ,\u2_Display/n3068 ,\u2_Display/n3069 ,\u2_Display/n3070 ,\u2_Display/n3071 ,\u2_Display/n3072 ,\u2_Display/n3073 ,\u2_Display/n3074 ,\u2_Display/n3075 ,\u2_Display/n3076 ,\u2_Display/n3077 ,\u2_Display/n3078 ,\u2_Display/n3079 ,\u2_Display/n3080 ,\u2_Display/n3081 ,\u2_Display/n3082 }),
    .i1(32'b11111111111101101001111111111111),
    .i2(1'b1),
    .o(\u2_Display/n3085 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add97  (
    .i0({\u2_Display/n3086 ,\u2_Display/n3087 ,\u2_Display/n3088 ,\u2_Display/n3089 ,\u2_Display/n3090 ,\u2_Display/n3091 ,\u2_Display/n3092 ,\u2_Display/n3093 ,\u2_Display/n3094 ,\u2_Display/n3095 ,\u2_Display/n3096 ,\u2_Display/n3097 ,\u2_Display/n3098 ,\u2_Display/n3099 ,\u2_Display/n3100 ,\u2_Display/n3101 ,\u2_Display/n3102 ,\u2_Display/n3103 ,\u2_Display/n3104 ,\u2_Display/n3105 ,\u2_Display/n3106 ,\u2_Display/n3107 ,\u2_Display/n3108 ,\u2_Display/n3109 ,\u2_Display/n3110 ,\u2_Display/n3111 ,\u2_Display/n3112 ,\u2_Display/n3113 ,\u2_Display/n3114 ,\u2_Display/n3115 ,\u2_Display/n3116 ,\u2_Display/n3117 }),
    .i1(32'b11111111111110110100111111111111),
    .i2(1'b1),
    .o(\u2_Display/n3120 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add98  (
    .i0({\u2_Display/n3121 ,\u2_Display/n3122 ,\u2_Display/n3123 ,\u2_Display/n3124 ,\u2_Display/n3125 ,\u2_Display/n3126 ,\u2_Display/n3127 ,\u2_Display/n3128 ,\u2_Display/n3129 ,\u2_Display/n3130 ,\u2_Display/n3131 ,\u2_Display/n3132 ,\u2_Display/n3133 ,\u2_Display/n3134 ,\u2_Display/n3135 ,\u2_Display/n3136 ,\u2_Display/n3137 ,\u2_Display/n3138 ,\u2_Display/n3139 ,\u2_Display/n3140 ,\u2_Display/n3141 ,\u2_Display/n3142 ,\u2_Display/n3143 ,\u2_Display/n3144 ,\u2_Display/n3145 ,\u2_Display/n3146 ,\u2_Display/n3147 ,\u2_Display/n3148 ,\u2_Display/n3149 ,\u2_Display/n3150 ,\u2_Display/n3151 ,\u2_Display/n3152 }),
    .i1(32'b11111111111111011010011111111111),
    .i2(1'b1),
    .o(\u2_Display/n3155 ));  // source/rtl/Display.v(196)
  add_pu32_pu32_pu1_o32 \u2_Display/add99  (
    .i0({\u2_Display/n3156 ,\u2_Display/n3157 ,\u2_Display/n3158 ,\u2_Display/n3159 ,\u2_Display/n3160 ,\u2_Display/n3161 ,\u2_Display/n3162 ,\u2_Display/n3163 ,\u2_Display/n3164 ,\u2_Display/n3165 ,\u2_Display/n3166 ,\u2_Display/n3167 ,\u2_Display/n3168 ,\u2_Display/n3169 ,\u2_Display/n3170 ,\u2_Display/n3171 ,\u2_Display/n3172 ,\u2_Display/n3173 ,\u2_Display/n3174 ,\u2_Display/n3175 ,\u2_Display/n3176 ,\u2_Display/n3177 ,\u2_Display/n3178 ,\u2_Display/n3179 ,\u2_Display/n3180 ,\u2_Display/n3181 ,\u2_Display/n3182 ,\u2_Display/n3183 ,\u2_Display/n3184 ,\u2_Display/n3185 ,\u2_Display/n3186 ,\u2_Display/n3187 }),
    .i1(32'b11111111111111101101001111111111),
    .i2(1'b1),
    .o(\u2_Display/n3190 ));  // source/rtl/Display.v(196)
  reg_ar_as_w1 \u2_Display/clk1s_reg  (
    .clk(clk_vga),
    .d(\u2_Display/n36 ),
    .en(\u2_Display/n35 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/clk1s ));  // source/rtl/Display.v(61)
  eq_w31 \u2_Display/eq0  (
    .i0(\u2_Display/n ),
    .i1(31'b0000000000000000010011100010000),
    .o(\u2_Display/n35 ));  // source/rtl/Display.v(52)
  lt_u12_u12 \u2_Display/lt0_2  (
    .ci(1'b0),
    .i0(lcd_xpos),
    .i1({\u2_Display/add2_2_co ,\u2_Display/n43 [2:0],\u2_Display/i [7:0]}),
    .o(\u2_Display/n44 ));  // source/rtl/Display.v(165)
  lt_u12_u12 \u2_Display/lt1  (
    .ci(1'b0),
    .i0({1'b0,\u2_Display/i [10:0]}),
    .i1(lcd_xpos),
    .o(\u2_Display/n45 ));  // source/rtl/Display.v(165)
  lt_u32_u32 \u2_Display/lt100  (
    .ci(1'b0),
    .i0({\u2_Display/n3051 ,\u2_Display/n3052 ,\u2_Display/n3053 ,\u2_Display/n3054 ,\u2_Display/n3055 ,\u2_Display/n3056 ,\u2_Display/n3057 ,\u2_Display/n3058 ,\u2_Display/n3059 ,\u2_Display/n3060 ,\u2_Display/n3061 ,\u2_Display/n3062 ,\u2_Display/n3063 ,\u2_Display/n3064 ,\u2_Display/n3065 ,\u2_Display/n3066 ,\u2_Display/n3067 ,\u2_Display/n3068 ,\u2_Display/n3069 ,\u2_Display/n3070 ,\u2_Display/n3071 ,\u2_Display/n3072 ,\u2_Display/n3073 ,\u2_Display/n3074 ,\u2_Display/n3075 ,\u2_Display/n3076 ,\u2_Display/n3077 ,\u2_Display/n3078 ,\u2_Display/n3079 ,\u2_Display/n3080 ,\u2_Display/n3081 ,\u2_Display/n3082 }),
    .i1(32'b00000000000010010110000000000000),
    .o(\u2_Display/n3083 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt101  (
    .ci(1'b0),
    .i0({\u2_Display/n3086 ,\u2_Display/n3087 ,\u2_Display/n3088 ,\u2_Display/n3089 ,\u2_Display/n3090 ,\u2_Display/n3091 ,\u2_Display/n3092 ,\u2_Display/n3093 ,\u2_Display/n3094 ,\u2_Display/n3095 ,\u2_Display/n3096 ,\u2_Display/n3097 ,\u2_Display/n3098 ,\u2_Display/n3099 ,\u2_Display/n3100 ,\u2_Display/n3101 ,\u2_Display/n3102 ,\u2_Display/n3103 ,\u2_Display/n3104 ,\u2_Display/n3105 ,\u2_Display/n3106 ,\u2_Display/n3107 ,\u2_Display/n3108 ,\u2_Display/n3109 ,\u2_Display/n3110 ,\u2_Display/n3111 ,\u2_Display/n3112 ,\u2_Display/n3113 ,\u2_Display/n3114 ,\u2_Display/n3115 ,\u2_Display/n3116 ,\u2_Display/n3117 }),
    .i1(32'b00000000000001001011000000000000),
    .o(\u2_Display/n3118 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt102  (
    .ci(1'b0),
    .i0({\u2_Display/n3121 ,\u2_Display/n3122 ,\u2_Display/n3123 ,\u2_Display/n3124 ,\u2_Display/n3125 ,\u2_Display/n3126 ,\u2_Display/n3127 ,\u2_Display/n3128 ,\u2_Display/n3129 ,\u2_Display/n3130 ,\u2_Display/n3131 ,\u2_Display/n3132 ,\u2_Display/n3133 ,\u2_Display/n3134 ,\u2_Display/n3135 ,\u2_Display/n3136 ,\u2_Display/n3137 ,\u2_Display/n3138 ,\u2_Display/n3139 ,\u2_Display/n3140 ,\u2_Display/n3141 ,\u2_Display/n3142 ,\u2_Display/n3143 ,\u2_Display/n3144 ,\u2_Display/n3145 ,\u2_Display/n3146 ,\u2_Display/n3147 ,\u2_Display/n3148 ,\u2_Display/n3149 ,\u2_Display/n3150 ,\u2_Display/n3151 ,\u2_Display/n3152 }),
    .i1(32'b00000000000000100101100000000000),
    .o(\u2_Display/n3153 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt103  (
    .ci(1'b0),
    .i0({\u2_Display/n3156 ,\u2_Display/n3157 ,\u2_Display/n3158 ,\u2_Display/n3159 ,\u2_Display/n3160 ,\u2_Display/n3161 ,\u2_Display/n3162 ,\u2_Display/n3163 ,\u2_Display/n3164 ,\u2_Display/n3165 ,\u2_Display/n3166 ,\u2_Display/n3167 ,\u2_Display/n3168 ,\u2_Display/n3169 ,\u2_Display/n3170 ,\u2_Display/n3171 ,\u2_Display/n3172 ,\u2_Display/n3173 ,\u2_Display/n3174 ,\u2_Display/n3175 ,\u2_Display/n3176 ,\u2_Display/n3177 ,\u2_Display/n3178 ,\u2_Display/n3179 ,\u2_Display/n3180 ,\u2_Display/n3181 ,\u2_Display/n3182 ,\u2_Display/n3183 ,\u2_Display/n3184 ,\u2_Display/n3185 ,\u2_Display/n3186 ,\u2_Display/n3187 }),
    .i1(32'b00000000000000010010110000000000),
    .o(\u2_Display/n3188 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt104  (
    .ci(1'b0),
    .i0({\u2_Display/n3191 ,\u2_Display/n3192 ,\u2_Display/n3193 ,\u2_Display/n3194 ,\u2_Display/n3195 ,\u2_Display/n3196 ,\u2_Display/n3197 ,\u2_Display/n3198 ,\u2_Display/n3199 ,\u2_Display/n3200 ,\u2_Display/n3201 ,\u2_Display/n3202 ,\u2_Display/n3203 ,\u2_Display/n3204 ,\u2_Display/n3205 ,\u2_Display/n3206 ,\u2_Display/n3207 ,\u2_Display/n3208 ,\u2_Display/n3209 ,\u2_Display/n3210 ,\u2_Display/n3211 ,\u2_Display/n3212 ,\u2_Display/n3213 ,\u2_Display/n3214 ,\u2_Display/n3215 ,\u2_Display/n3216 ,\u2_Display/n3217 ,\u2_Display/n3218 ,\u2_Display/n3219 ,\u2_Display/n3220 ,\u2_Display/n3221 ,\u2_Display/n3222 }),
    .i1(32'b00000000000000001001011000000000),
    .o(\u2_Display/n3223 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt105  (
    .ci(1'b0),
    .i0({\u2_Display/n3226 ,\u2_Display/n3227 ,\u2_Display/n3228 ,\u2_Display/n3229 ,\u2_Display/n3230 ,\u2_Display/n3231 ,\u2_Display/n3232 ,\u2_Display/n3233 ,\u2_Display/n3234 ,\u2_Display/n3235 ,\u2_Display/n3236 ,\u2_Display/n3237 ,\u2_Display/n3238 ,\u2_Display/n3239 ,\u2_Display/n3240 ,\u2_Display/n3241 ,\u2_Display/n3242 ,\u2_Display/n3243 ,\u2_Display/n3244 ,\u2_Display/n3245 ,\u2_Display/n3246 ,\u2_Display/n3247 ,\u2_Display/n3248 ,\u2_Display/n3249 ,\u2_Display/n3250 ,\u2_Display/n3251 ,\u2_Display/n3252 ,\u2_Display/n3253 ,\u2_Display/n3254 ,\u2_Display/n3255 ,\u2_Display/n3256 ,\u2_Display/n3257 }),
    .i1(32'b00000000000000000100101100000000),
    .o(\u2_Display/n3258 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt106  (
    .ci(1'b0),
    .i0({\u2_Display/n3261 ,\u2_Display/n3262 ,\u2_Display/n3263 ,\u2_Display/n3264 ,\u2_Display/n3265 ,\u2_Display/n3266 ,\u2_Display/n3267 ,\u2_Display/n3268 ,\u2_Display/n3269 ,\u2_Display/n3270 ,\u2_Display/n3271 ,\u2_Display/n3272 ,\u2_Display/n3273 ,\u2_Display/n3274 ,\u2_Display/n3275 ,\u2_Display/n3276 ,\u2_Display/n3277 ,\u2_Display/n3278 ,\u2_Display/n3279 ,\u2_Display/n3280 ,\u2_Display/n3281 ,\u2_Display/n3282 ,\u2_Display/n3283 ,\u2_Display/n3284 ,\u2_Display/n3285 ,\u2_Display/n3286 ,\u2_Display/n3287 ,\u2_Display/n3288 ,\u2_Display/n3289 ,\u2_Display/n3290 ,\u2_Display/n3291 ,\u2_Display/n3292 }),
    .i1(32'b00000000000000000010010110000000),
    .o(\u2_Display/n3293 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt107  (
    .ci(1'b0),
    .i0({\u2_Display/n3296 ,\u2_Display/n3297 ,\u2_Display/n3298 ,\u2_Display/n3299 ,\u2_Display/n3300 ,\u2_Display/n3301 ,\u2_Display/n3302 ,\u2_Display/n3303 ,\u2_Display/n3304 ,\u2_Display/n3305 ,\u2_Display/n3306 ,\u2_Display/n3307 ,\u2_Display/n3308 ,\u2_Display/n3309 ,\u2_Display/n3310 ,\u2_Display/n3311 ,\u2_Display/n3312 ,\u2_Display/n3313 ,\u2_Display/n3314 ,\u2_Display/n3315 ,\u2_Display/n3316 ,\u2_Display/n3317 ,\u2_Display/n3318 ,\u2_Display/n3319 ,\u2_Display/n3320 ,\u2_Display/n3321 ,\u2_Display/n3322 ,\u2_Display/n3323 ,\u2_Display/n3324 ,\u2_Display/n3325 ,\u2_Display/n3326 ,\u2_Display/n3327 }),
    .i1(32'b00000000000000000001001011000000),
    .o(\u2_Display/n3328 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt108  (
    .ci(1'b0),
    .i0({\u2_Display/n3331 ,\u2_Display/n3332 ,\u2_Display/n3333 ,\u2_Display/n3334 ,\u2_Display/n3335 ,\u2_Display/n3336 ,\u2_Display/n3337 ,\u2_Display/n3338 ,\u2_Display/n3339 ,\u2_Display/n3340 ,\u2_Display/n3341 ,\u2_Display/n3342 ,\u2_Display/n3343 ,\u2_Display/n3344 ,\u2_Display/n3345 ,\u2_Display/n3346 ,\u2_Display/n3347 ,\u2_Display/n3348 ,\u2_Display/n3349 ,\u2_Display/n3350 ,\u2_Display/n3351 ,\u2_Display/n3352 ,\u2_Display/n3353 ,\u2_Display/n3354 ,\u2_Display/n3355 ,\u2_Display/n3356 ,\u2_Display/n3357 ,\u2_Display/n3358 ,\u2_Display/n3359 ,\u2_Display/n3360 ,\u2_Display/n3361 ,\u2_Display/n3362 }),
    .i1(32'b00000000000000000000100101100000),
    .o(\u2_Display/n3363 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt109  (
    .ci(1'b0),
    .i0({\u2_Display/n3366 ,\u2_Display/n3367 ,\u2_Display/n3368 ,\u2_Display/n3369 ,\u2_Display/n3370 ,\u2_Display/n3371 ,\u2_Display/n3372 ,\u2_Display/n3373 ,\u2_Display/n3374 ,\u2_Display/n3375 ,\u2_Display/n3376 ,\u2_Display/n3377 ,\u2_Display/n3378 ,\u2_Display/n3379 ,\u2_Display/n3380 ,\u2_Display/n3381 ,\u2_Display/n3382 ,\u2_Display/n3383 ,\u2_Display/n3384 ,\u2_Display/n3385 ,\u2_Display/n3386 ,\u2_Display/n3387 ,\u2_Display/n3388 ,\u2_Display/n3389 ,\u2_Display/n3390 ,\u2_Display/n3391 ,\u2_Display/n3392 ,\u2_Display/n3393 ,\u2_Display/n3394 ,\u2_Display/n3395 ,\u2_Display/n3396 ,\u2_Display/n3397 }),
    .i1(32'b00000000000000000000010010110000),
    .o(\u2_Display/n3398 ));  // source/rtl/Display.v(196)
  lt_u12_u12 \u2_Display/lt10_2  (
    .ci(1'b0),
    .i0(lcd_ypos),
    .i1({\u2_Display/add7_2_co ,\u2_Display/n140 [1:0],\u2_Display/i [8:0]}),
    .o(\u2_Display/n141 ));  // source/rtl/Display.v(197)
  lt_u32_u32 \u2_Display/lt110  (
    .ci(1'b0),
    .i0({\u2_Display/n3401 ,\u2_Display/n3402 ,\u2_Display/n3403 ,\u2_Display/n3404 ,\u2_Display/n3405 ,\u2_Display/n3406 ,\u2_Display/n3407 ,\u2_Display/n3408 ,\u2_Display/n3409 ,\u2_Display/n3410 ,\u2_Display/n3411 ,\u2_Display/n3412 ,\u2_Display/n3413 ,\u2_Display/n3414 ,\u2_Display/n3415 ,\u2_Display/n3416 ,\u2_Display/n3417 ,\u2_Display/n3418 ,\u2_Display/n3419 ,\u2_Display/n3420 ,\u2_Display/n3421 ,\u2_Display/n3422 ,\u2_Display/n3423 ,\u2_Display/n3424 ,\u2_Display/n3425 ,\u2_Display/n3426 ,\u2_Display/n3427 ,\u2_Display/n3428 ,\u2_Display/n3429 ,\u2_Display/n3430 ,\u2_Display/n3431 ,\u2_Display/n3432 }),
    .i1(32'b00000000000000000000001001011000),
    .o(\u2_Display/n3433 ));  // source/rtl/Display.v(196)
  lt_u13_u13 \u2_Display/lt11_2  (
    .ci(1'b0),
    .i0({\u2_Display/n143 [31],\u2_Display/n143 [31],\u2_Display/n143 [10:0]}),
    .i1({1'b0,lcd_ypos}),
    .o(\u2_Display/n144 ));  // source/rtl/Display.v(197)
  lt_u32_u32 \u2_Display/lt121  (
    .ci(1'b0),
    .i0(\u2_Display/counta ),
    .i1(32'b11001000000000000000000000000000),
    .o(\u2_Display/n3786 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt122  (
    .ci(1'b0),
    .i0({\u2_Display/n3789 ,\u2_Display/n3790 ,\u2_Display/n3791 ,\u2_Display/n3792 ,\u2_Display/n3793 ,\u2_Display/n3794 ,\u2_Display/n3795 ,\u2_Display/n3796 ,\u2_Display/n3797 ,\u2_Display/n3798 ,\u2_Display/n3799 ,\u2_Display/n3800 ,\u2_Display/n3801 ,\u2_Display/n3802 ,\u2_Display/n3803 ,\u2_Display/n3804 ,\u2_Display/n3805 ,\u2_Display/n3806 ,\u2_Display/n3807 ,\u2_Display/n3808 ,\u2_Display/n3809 ,\u2_Display/n3810 ,\u2_Display/n3811 ,\u2_Display/n3812 ,\u2_Display/n3813 ,\u2_Display/n3814 ,\u2_Display/n3815 ,\u2_Display/n3816 ,\u2_Display/n3817 ,\u2_Display/n3818 ,\u2_Display/n3819 ,\u2_Display/n3820 }),
    .i1(32'b01100100000000000000000000000000),
    .o(\u2_Display/n3821 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt123  (
    .ci(1'b0),
    .i0({\u2_Display/n3824 ,\u2_Display/n3825 ,\u2_Display/n3826 ,\u2_Display/n3827 ,\u2_Display/n3828 ,\u2_Display/n3829 ,\u2_Display/n3830 ,\u2_Display/n3831 ,\u2_Display/n3832 ,\u2_Display/n3833 ,\u2_Display/n3834 ,\u2_Display/n3835 ,\u2_Display/n3836 ,\u2_Display/n3837 ,\u2_Display/n3838 ,\u2_Display/n3839 ,\u2_Display/n3840 ,\u2_Display/n3841 ,\u2_Display/n3842 ,\u2_Display/n3843 ,\u2_Display/n3844 ,\u2_Display/n3845 ,\u2_Display/n3846 ,\u2_Display/n3847 ,\u2_Display/n3848 ,\u2_Display/n3849 ,\u2_Display/n3850 ,\u2_Display/n3851 ,\u2_Display/n3852 ,\u2_Display/n3853 ,\u2_Display/n3854 ,\u2_Display/n3855 }),
    .i1(32'b00110010000000000000000000000000),
    .o(\u2_Display/n3856 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt124  (
    .ci(1'b0),
    .i0({\u2_Display/n3859 ,\u2_Display/n3860 ,\u2_Display/n3861 ,\u2_Display/n3862 ,\u2_Display/n3863 ,\u2_Display/n3864 ,\u2_Display/n3865 ,\u2_Display/n3866 ,\u2_Display/n3867 ,\u2_Display/n3868 ,\u2_Display/n3869 ,\u2_Display/n3870 ,\u2_Display/n3871 ,\u2_Display/n3872 ,\u2_Display/n3873 ,\u2_Display/n3874 ,\u2_Display/n3875 ,\u2_Display/n3876 ,\u2_Display/n3877 ,\u2_Display/n3878 ,\u2_Display/n3879 ,\u2_Display/n3880 ,\u2_Display/n3881 ,\u2_Display/n3882 ,\u2_Display/n3883 ,\u2_Display/n3884 ,\u2_Display/n3885 ,\u2_Display/n3886 ,\u2_Display/n3887 ,\u2_Display/n3888 ,\u2_Display/n3889 ,\u2_Display/n3890 }),
    .i1(32'b00011001000000000000000000000000),
    .o(\u2_Display/n3891 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt125  (
    .ci(1'b0),
    .i0({\u2_Display/n3894 ,\u2_Display/n3895 ,\u2_Display/n3896 ,\u2_Display/n3897 ,\u2_Display/n3898 ,\u2_Display/n3899 ,\u2_Display/n3900 ,\u2_Display/n3901 ,\u2_Display/n3902 ,\u2_Display/n3903 ,\u2_Display/n3904 ,\u2_Display/n3905 ,\u2_Display/n3906 ,\u2_Display/n3907 ,\u2_Display/n3908 ,\u2_Display/n3909 ,\u2_Display/n3910 ,\u2_Display/n3911 ,\u2_Display/n3912 ,\u2_Display/n3913 ,\u2_Display/n3914 ,\u2_Display/n3915 ,\u2_Display/n3916 ,\u2_Display/n3917 ,\u2_Display/n3918 ,\u2_Display/n3919 ,\u2_Display/n3920 ,\u2_Display/n3921 ,\u2_Display/n3922 ,\u2_Display/n3923 ,\u2_Display/n3924 ,\u2_Display/n3925 }),
    .i1(32'b00001100100000000000000000000000),
    .o(\u2_Display/n3926 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt126  (
    .ci(1'b0),
    .i0({\u2_Display/n3929 ,\u2_Display/n3930 ,\u2_Display/n3931 ,\u2_Display/n3932 ,\u2_Display/n3933 ,\u2_Display/n3934 ,\u2_Display/n3935 ,\u2_Display/n3936 ,\u2_Display/n3937 ,\u2_Display/n3938 ,\u2_Display/n3939 ,\u2_Display/n3940 ,\u2_Display/n3941 ,\u2_Display/n3942 ,\u2_Display/n3943 ,\u2_Display/n3944 ,\u2_Display/n3945 ,\u2_Display/n3946 ,\u2_Display/n3947 ,\u2_Display/n3948 ,\u2_Display/n3949 ,\u2_Display/n3950 ,\u2_Display/n3951 ,\u2_Display/n3952 ,\u2_Display/n3953 ,\u2_Display/n3954 ,\u2_Display/n3955 ,\u2_Display/n3956 ,\u2_Display/n3957 ,\u2_Display/n3958 ,\u2_Display/n3959 ,\u2_Display/n3960 }),
    .i1(32'b00000110010000000000000000000000),
    .o(\u2_Display/n3961 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt127  (
    .ci(1'b0),
    .i0({\u2_Display/n3964 ,\u2_Display/n3965 ,\u2_Display/n3966 ,\u2_Display/n3967 ,\u2_Display/n3968 ,\u2_Display/n3969 ,\u2_Display/n3970 ,\u2_Display/n3971 ,\u2_Display/n3972 ,\u2_Display/n3973 ,\u2_Display/n3974 ,\u2_Display/n3975 ,\u2_Display/n3976 ,\u2_Display/n3977 ,\u2_Display/n3978 ,\u2_Display/n3979 ,\u2_Display/n3980 ,\u2_Display/n3981 ,\u2_Display/n3982 ,\u2_Display/n3983 ,\u2_Display/n3984 ,\u2_Display/n3985 ,\u2_Display/n3986 ,\u2_Display/n3987 ,\u2_Display/n3988 ,\u2_Display/n3989 ,\u2_Display/n3990 ,\u2_Display/n3991 ,\u2_Display/n3992 ,\u2_Display/n3993 ,\u2_Display/n3994 ,\u2_Display/n3995 }),
    .i1(32'b00000011001000000000000000000000),
    .o(\u2_Display/n3996 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt128  (
    .ci(1'b0),
    .i0({\u2_Display/n3999 ,\u2_Display/n4000 ,\u2_Display/n4001 ,\u2_Display/n4002 ,\u2_Display/n4003 ,\u2_Display/n4004 ,\u2_Display/n4005 ,\u2_Display/n4006 ,\u2_Display/n4007 ,\u2_Display/n4008 ,\u2_Display/n4009 ,\u2_Display/n4010 ,\u2_Display/n4011 ,\u2_Display/n4012 ,\u2_Display/n4013 ,\u2_Display/n4014 ,\u2_Display/n4015 ,\u2_Display/n4016 ,\u2_Display/n4017 ,\u2_Display/n4018 ,\u2_Display/n4019 ,\u2_Display/n4020 ,\u2_Display/n4021 ,\u2_Display/n4022 ,\u2_Display/n4023 ,\u2_Display/n4024 ,\u2_Display/n4025 ,\u2_Display/n4026 ,\u2_Display/n4027 ,\u2_Display/n4028 ,\u2_Display/n4029 ,\u2_Display/n4030 }),
    .i1(32'b00000001100100000000000000000000),
    .o(\u2_Display/n4031 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt129  (
    .ci(1'b0),
    .i0({\u2_Display/n4034 ,\u2_Display/n4035 ,\u2_Display/n4036 ,\u2_Display/n4037 ,\u2_Display/n4038 ,\u2_Display/n4039 ,\u2_Display/n4040 ,\u2_Display/n4041 ,\u2_Display/n4042 ,\u2_Display/n4043 ,\u2_Display/n4044 ,\u2_Display/n4045 ,\u2_Display/n4046 ,\u2_Display/n4047 ,\u2_Display/n4048 ,\u2_Display/n4049 ,\u2_Display/n4050 ,\u2_Display/n4051 ,\u2_Display/n4052 ,\u2_Display/n4053 ,\u2_Display/n4054 ,\u2_Display/n4055 ,\u2_Display/n4056 ,\u2_Display/n4057 ,\u2_Display/n4058 ,\u2_Display/n4059 ,\u2_Display/n4060 ,\u2_Display/n4061 ,\u2_Display/n4062 ,\u2_Display/n4063 ,\u2_Display/n4064 ,\u2_Display/n4065 }),
    .i1(32'b00000000110010000000000000000000),
    .o(\u2_Display/n4066 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt130  (
    .ci(1'b0),
    .i0({\u2_Display/n4069 ,\u2_Display/n4070 ,\u2_Display/n4071 ,\u2_Display/n4072 ,\u2_Display/n4073 ,\u2_Display/n4074 ,\u2_Display/n4075 ,\u2_Display/n4076 ,\u2_Display/n4077 ,\u2_Display/n4078 ,\u2_Display/n4079 ,\u2_Display/n4080 ,\u2_Display/n4081 ,\u2_Display/n4082 ,\u2_Display/n4083 ,\u2_Display/n4084 ,\u2_Display/n4085 ,\u2_Display/n4086 ,\u2_Display/n4087 ,\u2_Display/n4088 ,\u2_Display/n4089 ,\u2_Display/n4090 ,\u2_Display/n4091 ,\u2_Display/n4092 ,\u2_Display/n4093 ,\u2_Display/n4094 ,\u2_Display/n4095 ,\u2_Display/n4096 ,\u2_Display/n4097 ,\u2_Display/n4098 ,\u2_Display/n4099 ,\u2_Display/n4100 }),
    .i1(32'b00000000011001000000000000000000),
    .o(\u2_Display/n4101 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt131  (
    .ci(1'b0),
    .i0({\u2_Display/n4104 ,\u2_Display/n4105 ,\u2_Display/n4106 ,\u2_Display/n4107 ,\u2_Display/n4108 ,\u2_Display/n4109 ,\u2_Display/n4110 ,\u2_Display/n4111 ,\u2_Display/n4112 ,\u2_Display/n4113 ,\u2_Display/n4114 ,\u2_Display/n4115 ,\u2_Display/n4116 ,\u2_Display/n4117 ,\u2_Display/n4118 ,\u2_Display/n4119 ,\u2_Display/n4120 ,\u2_Display/n4121 ,\u2_Display/n4122 ,\u2_Display/n4123 ,\u2_Display/n4124 ,\u2_Display/n4125 ,\u2_Display/n4126 ,\u2_Display/n4127 ,\u2_Display/n4128 ,\u2_Display/n4129 ,\u2_Display/n4130 ,\u2_Display/n4131 ,\u2_Display/n4132 ,\u2_Display/n4133 ,\u2_Display/n4134 ,\u2_Display/n4135 }),
    .i1(32'b00000000001100100000000000000000),
    .o(\u2_Display/n4136 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt132  (
    .ci(1'b0),
    .i0({\u2_Display/n4139 ,\u2_Display/n4140 ,\u2_Display/n4141 ,\u2_Display/n4142 ,\u2_Display/n4143 ,\u2_Display/n4144 ,\u2_Display/n4145 ,\u2_Display/n4146 ,\u2_Display/n4147 ,\u2_Display/n4148 ,\u2_Display/n4149 ,\u2_Display/n4150 ,\u2_Display/n4151 ,\u2_Display/n4152 ,\u2_Display/n4153 ,\u2_Display/n4154 ,\u2_Display/n4155 ,\u2_Display/n4156 ,\u2_Display/n4157 ,\u2_Display/n4158 ,\u2_Display/n4159 ,\u2_Display/n4160 ,\u2_Display/n4161 ,\u2_Display/n4162 ,\u2_Display/n4163 ,\u2_Display/n4164 ,\u2_Display/n4165 ,\u2_Display/n4166 ,\u2_Display/n4167 ,\u2_Display/n4168 ,\u2_Display/n4169 ,\u2_Display/n4170 }),
    .i1(32'b00000000000110010000000000000000),
    .o(\u2_Display/n4171 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt133  (
    .ci(1'b0),
    .i0({\u2_Display/n4174 ,\u2_Display/n4175 ,\u2_Display/n4176 ,\u2_Display/n4177 ,\u2_Display/n4178 ,\u2_Display/n4179 ,\u2_Display/n4180 ,\u2_Display/n4181 ,\u2_Display/n4182 ,\u2_Display/n4183 ,\u2_Display/n4184 ,\u2_Display/n4185 ,\u2_Display/n4186 ,\u2_Display/n4187 ,\u2_Display/n4188 ,\u2_Display/n4189 ,\u2_Display/n4190 ,\u2_Display/n4191 ,\u2_Display/n4192 ,\u2_Display/n4193 ,\u2_Display/n4194 ,\u2_Display/n4195 ,\u2_Display/n4196 ,\u2_Display/n4197 ,\u2_Display/n4198 ,\u2_Display/n4199 ,\u2_Display/n4200 ,\u2_Display/n4201 ,\u2_Display/n4202 ,\u2_Display/n4203 ,\u2_Display/n4204 ,\u2_Display/n4205 }),
    .i1(32'b00000000000011001000000000000000),
    .o(\u2_Display/n4206 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt134  (
    .ci(1'b0),
    .i0({\u2_Display/n4209 ,\u2_Display/n4210 ,\u2_Display/n4211 ,\u2_Display/n4212 ,\u2_Display/n4213 ,\u2_Display/n4214 ,\u2_Display/n4215 ,\u2_Display/n4216 ,\u2_Display/n4217 ,\u2_Display/n4218 ,\u2_Display/n4219 ,\u2_Display/n4220 ,\u2_Display/n4221 ,\u2_Display/n4222 ,\u2_Display/n4223 ,\u2_Display/n4224 ,\u2_Display/n4225 ,\u2_Display/n4226 ,\u2_Display/n4227 ,\u2_Display/n4228 ,\u2_Display/n4229 ,\u2_Display/n4230 ,\u2_Display/n4231 ,\u2_Display/n4232 ,\u2_Display/n4233 ,\u2_Display/n4234 ,\u2_Display/n4235 ,\u2_Display/n4236 ,\u2_Display/n4237 ,\u2_Display/n4238 ,\u2_Display/n4239 ,\u2_Display/n4240 }),
    .i1(32'b00000000000001100100000000000000),
    .o(\u2_Display/n4241 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt135  (
    .ci(1'b0),
    .i0({\u2_Display/n4244 ,\u2_Display/n4245 ,\u2_Display/n4246 ,\u2_Display/n4247 ,\u2_Display/n4248 ,\u2_Display/n4249 ,\u2_Display/n4250 ,\u2_Display/n4251 ,\u2_Display/n4252 ,\u2_Display/n4253 ,\u2_Display/n4254 ,\u2_Display/n4255 ,\u2_Display/n4256 ,\u2_Display/n4257 ,\u2_Display/n4258 ,\u2_Display/n4259 ,\u2_Display/n4260 ,\u2_Display/n4261 ,\u2_Display/n4262 ,\u2_Display/n4263 ,\u2_Display/n4264 ,\u2_Display/n4265 ,\u2_Display/n4266 ,\u2_Display/n4267 ,\u2_Display/n4268 ,\u2_Display/n4269 ,\u2_Display/n4270 ,\u2_Display/n4271 ,\u2_Display/n4272 ,\u2_Display/n4273 ,\u2_Display/n4274 ,\u2_Display/n4275 }),
    .i1(32'b00000000000000110010000000000000),
    .o(\u2_Display/n4276 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt136  (
    .ci(1'b0),
    .i0({\u2_Display/n4279 ,\u2_Display/n4280 ,\u2_Display/n4281 ,\u2_Display/n4282 ,\u2_Display/n4283 ,\u2_Display/n4284 ,\u2_Display/n4285 ,\u2_Display/n4286 ,\u2_Display/n4287 ,\u2_Display/n4288 ,\u2_Display/n4289 ,\u2_Display/n4290 ,\u2_Display/n4291 ,\u2_Display/n4292 ,\u2_Display/n4293 ,\u2_Display/n4294 ,\u2_Display/n4295 ,\u2_Display/n4296 ,\u2_Display/n4297 ,\u2_Display/n4298 ,\u2_Display/n4299 ,\u2_Display/n4300 ,\u2_Display/n4301 ,\u2_Display/n4302 ,\u2_Display/n4303 ,\u2_Display/n4304 ,\u2_Display/n4305 ,\u2_Display/n4306 ,\u2_Display/n4307 ,\u2_Display/n4308 ,\u2_Display/n4309 ,\u2_Display/n4310 }),
    .i1(32'b00000000000000011001000000000000),
    .o(\u2_Display/n4311 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt137  (
    .ci(1'b0),
    .i0({\u2_Display/n4314 ,\u2_Display/n4315 ,\u2_Display/n4316 ,\u2_Display/n4317 ,\u2_Display/n4318 ,\u2_Display/n4319 ,\u2_Display/n4320 ,\u2_Display/n4321 ,\u2_Display/n4322 ,\u2_Display/n4323 ,\u2_Display/n4324 ,\u2_Display/n4325 ,\u2_Display/n4326 ,\u2_Display/n4327 ,\u2_Display/n4328 ,\u2_Display/n4329 ,\u2_Display/n4330 ,\u2_Display/n4331 ,\u2_Display/n4332 ,\u2_Display/n4333 ,\u2_Display/n4334 ,\u2_Display/n4335 ,\u2_Display/n4336 ,\u2_Display/n4337 ,\u2_Display/n4338 ,\u2_Display/n4339 ,\u2_Display/n4340 ,\u2_Display/n4341 ,\u2_Display/n4342 ,\u2_Display/n4343 ,\u2_Display/n4344 ,\u2_Display/n4345 }),
    .i1(32'b00000000000000001100100000000000),
    .o(\u2_Display/n4346 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt138  (
    .ci(1'b0),
    .i0({\u2_Display/n4349 ,\u2_Display/n4350 ,\u2_Display/n4351 ,\u2_Display/n4352 ,\u2_Display/n4353 ,\u2_Display/n4354 ,\u2_Display/n4355 ,\u2_Display/n4356 ,\u2_Display/n4357 ,\u2_Display/n4358 ,\u2_Display/n4359 ,\u2_Display/n4360 ,\u2_Display/n4361 ,\u2_Display/n4362 ,\u2_Display/n4363 ,\u2_Display/n4364 ,\u2_Display/n4365 ,\u2_Display/n4366 ,\u2_Display/n4367 ,\u2_Display/n4368 ,\u2_Display/n4369 ,\u2_Display/n4370 ,\u2_Display/n4371 ,\u2_Display/n4372 ,\u2_Display/n4373 ,\u2_Display/n4374 ,\u2_Display/n4375 ,\u2_Display/n4376 ,\u2_Display/n4377 ,\u2_Display/n4378 ,\u2_Display/n4379 ,\u2_Display/n4380 }),
    .i1(32'b00000000000000000110010000000000),
    .o(\u2_Display/n4381 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt139  (
    .ci(1'b0),
    .i0({\u2_Display/n4384 ,\u2_Display/n4385 ,\u2_Display/n4386 ,\u2_Display/n4387 ,\u2_Display/n4388 ,\u2_Display/n4389 ,\u2_Display/n4390 ,\u2_Display/n4391 ,\u2_Display/n4392 ,\u2_Display/n4393 ,\u2_Display/n4394 ,\u2_Display/n4395 ,\u2_Display/n4396 ,\u2_Display/n4397 ,\u2_Display/n4398 ,\u2_Display/n4399 ,\u2_Display/n4400 ,\u2_Display/n4401 ,\u2_Display/n4402 ,\u2_Display/n4403 ,\u2_Display/n4404 ,\u2_Display/n4405 ,\u2_Display/n4406 ,\u2_Display/n4407 ,\u2_Display/n4408 ,\u2_Display/n4409 ,\u2_Display/n4410 ,\u2_Display/n4411 ,\u2_Display/n4412 ,\u2_Display/n4413 ,\u2_Display/n4414 ,\u2_Display/n4415 }),
    .i1(32'b00000000000000000011001000000000),
    .o(\u2_Display/n4416 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt140  (
    .ci(1'b0),
    .i0({\u2_Display/n4419 ,\u2_Display/n4420 ,\u2_Display/n4421 ,\u2_Display/n4422 ,\u2_Display/n4423 ,\u2_Display/n4424 ,\u2_Display/n4425 ,\u2_Display/n4426 ,\u2_Display/n4427 ,\u2_Display/n4428 ,\u2_Display/n4429 ,\u2_Display/n4430 ,\u2_Display/n4431 ,\u2_Display/n4432 ,\u2_Display/n4433 ,\u2_Display/n4434 ,\u2_Display/n4435 ,\u2_Display/n4436 ,\u2_Display/n4437 ,\u2_Display/n4438 ,\u2_Display/n4439 ,\u2_Display/n4440 ,\u2_Display/n4441 ,\u2_Display/n4442 ,\u2_Display/n4443 ,\u2_Display/n4444 ,\u2_Display/n4445 ,\u2_Display/n4446 ,\u2_Display/n4447 ,\u2_Display/n4448 ,\u2_Display/n4449 ,\u2_Display/n4450 }),
    .i1(32'b00000000000000000001100100000000),
    .o(\u2_Display/n4451 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt141  (
    .ci(1'b0),
    .i0({\u2_Display/n4454 ,\u2_Display/n4455 ,\u2_Display/n4456 ,\u2_Display/n4457 ,\u2_Display/n4458 ,\u2_Display/n4459 ,\u2_Display/n4460 ,\u2_Display/n4461 ,\u2_Display/n4462 ,\u2_Display/n4463 ,\u2_Display/n4464 ,\u2_Display/n4465 ,\u2_Display/n4466 ,\u2_Display/n4467 ,\u2_Display/n4468 ,\u2_Display/n4469 ,\u2_Display/n4470 ,\u2_Display/n4471 ,\u2_Display/n4472 ,\u2_Display/n4473 ,\u2_Display/n4474 ,\u2_Display/n4475 ,\u2_Display/n4476 ,\u2_Display/n4477 ,\u2_Display/n4478 ,\u2_Display/n4479 ,\u2_Display/n4480 ,\u2_Display/n4481 ,\u2_Display/n4482 ,\u2_Display/n4483 ,\u2_Display/n4484 ,\u2_Display/n4485 }),
    .i1(32'b00000000000000000000110010000000),
    .o(\u2_Display/n4486 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt142  (
    .ci(1'b0),
    .i0({\u2_Display/n4489 ,\u2_Display/n4490 ,\u2_Display/n4491 ,\u2_Display/n4492 ,\u2_Display/n4493 ,\u2_Display/n4494 ,\u2_Display/n4495 ,\u2_Display/n4496 ,\u2_Display/n4497 ,\u2_Display/n4498 ,\u2_Display/n4499 ,\u2_Display/n4500 ,\u2_Display/n4501 ,\u2_Display/n4502 ,\u2_Display/n4503 ,\u2_Display/n4504 ,\u2_Display/n4505 ,\u2_Display/n4506 ,\u2_Display/n4507 ,\u2_Display/n4508 ,\u2_Display/n4509 ,\u2_Display/n4510 ,\u2_Display/n4511 ,\u2_Display/n4512 ,\u2_Display/n4513 ,\u2_Display/n4514 ,\u2_Display/n4515 ,\u2_Display/n4516 ,\u2_Display/n4517 ,\u2_Display/n4518 ,\u2_Display/n4519 ,\u2_Display/n4520 }),
    .i1(32'b00000000000000000000011001000000),
    .o(\u2_Display/n4521 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt143  (
    .ci(1'b0),
    .i0({\u2_Display/n4524 ,\u2_Display/n4525 ,\u2_Display/n4526 ,\u2_Display/n4527 ,\u2_Display/n4528 ,\u2_Display/n4529 ,\u2_Display/n4530 ,\u2_Display/n4531 ,\u2_Display/n4532 ,\u2_Display/n4533 ,\u2_Display/n4534 ,\u2_Display/n4535 ,\u2_Display/n4536 ,\u2_Display/n4537 ,\u2_Display/n4538 ,\u2_Display/n4539 ,\u2_Display/n4540 ,\u2_Display/n4541 ,\u2_Display/n4542 ,\u2_Display/n4543 ,\u2_Display/n4544 ,\u2_Display/n4545 ,\u2_Display/n4546 ,\u2_Display/n4547 ,\u2_Display/n4548 ,\u2_Display/n4549 ,\u2_Display/n4550 ,\u2_Display/n4551 ,\u2_Display/n4552 ,\u2_Display/n4553 ,\u2_Display/n4554 ,\u2_Display/n4555 }),
    .i1(32'b00000000000000000000001100100000),
    .o(\u2_Display/n4556 ));  // source/rtl/Display.v(195)
  lt_u32_u32 \u2_Display/lt154  (
    .ci(1'b0),
    .i0(\u2_Display/counta ),
    .i1(32'b10100000000000000000000000000000),
    .o(\u2_Display/n4909 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt155  (
    .ci(1'b0),
    .i0({\u2_Display/n6070 ,\u2_Display/n6071 ,\u2_Display/n6072 ,\u2_Display/n6073 ,\u2_Display/n6074 ,\u2_Display/n6075 ,\u2_Display/n6076 ,\u2_Display/n6077 ,\u2_Display/n6078 ,\u2_Display/n6079 ,\u2_Display/n6080 ,\u2_Display/n6081 ,\u2_Display/n6082 ,\u2_Display/n6083 ,\u2_Display/n6084 ,\u2_Display/n6085 ,\u2_Display/n6086 ,\u2_Display/n6087 ,\u2_Display/n6088 ,\u2_Display/n6089 ,\u2_Display/n6090 ,\u2_Display/n6091 ,\u2_Display/n6092 ,\u2_Display/n6093 ,\u2_Display/n6094 ,\u2_Display/n6095 ,\u2_Display/n6096 ,\u2_Display/n6097 ,\u2_Display/n6098 ,\u2_Display/n6099 ,\u2_Display/n6100 ,\u2_Display/n6101 }),
    .i1(32'b01010000000000000000000000000000),
    .o(\u2_Display/n4944 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt156  (
    .ci(1'b0),
    .i0({\u2_Display/n6105 ,\u2_Display/n6106 ,\u2_Display/n6107 ,\u2_Display/n6108 ,\u2_Display/n6109 ,\u2_Display/n6110 ,\u2_Display/n6111 ,\u2_Display/n6112 ,\u2_Display/n6113 ,\u2_Display/n6114 ,\u2_Display/n6115 ,\u2_Display/n6116 ,\u2_Display/n6117 ,\u2_Display/n6118 ,\u2_Display/n6119 ,\u2_Display/n6120 ,\u2_Display/n6121 ,\u2_Display/n6122 ,\u2_Display/n6123 ,\u2_Display/n6124 ,\u2_Display/n6125 ,\u2_Display/n6126 ,\u2_Display/n6127 ,\u2_Display/n6128 ,\u2_Display/n6129 ,\u2_Display/n6130 ,\u2_Display/n6131 ,\u2_Display/n6132 ,\u2_Display/n6133 ,\u2_Display/n6134 ,\u2_Display/n6135 ,\u2_Display/n6136 }),
    .i1(32'b00101000000000000000000000000000),
    .o(\u2_Display/n4979 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt157  (
    .ci(1'b0),
    .i0({\u2_Display/n6140 ,\u2_Display/n6141 ,\u2_Display/n6142 ,\u2_Display/n6143 ,\u2_Display/n6144 ,\u2_Display/n6145 ,\u2_Display/n6146 ,\u2_Display/n6147 ,\u2_Display/n6148 ,\u2_Display/n6149 ,\u2_Display/n6150 ,\u2_Display/n6151 ,\u2_Display/n6152 ,\u2_Display/n6153 ,\u2_Display/n6154 ,\u2_Display/n6155 ,\u2_Display/n6156 ,\u2_Display/n6157 ,\u2_Display/n6158 ,\u2_Display/n6159 ,\u2_Display/n6160 ,\u2_Display/n6161 ,\u2_Display/n6162 ,\u2_Display/n6163 ,\u2_Display/n6164 ,\u2_Display/n6165 ,\u2_Display/n6166 ,\u2_Display/n6167 ,\u2_Display/n6168 ,\u2_Display/n6169 ,\u2_Display/n6170 ,\u2_Display/n6171 }),
    .i1(32'b00010100000000000000000000000000),
    .o(\u2_Display/n5014 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt158  (
    .ci(1'b0),
    .i0({\u2_Display/n6175 ,\u2_Display/n6176 ,\u2_Display/n6177 ,\u2_Display/n6178 ,\u2_Display/n6179 ,\u2_Display/n6180 ,\u2_Display/n6181 ,\u2_Display/n6182 ,\u2_Display/n6183 ,\u2_Display/n6184 ,\u2_Display/n6185 ,\u2_Display/n6186 ,\u2_Display/n6187 ,\u2_Display/n6188 ,\u2_Display/n6189 ,\u2_Display/n6190 ,\u2_Display/n6191 ,\u2_Display/n6192 ,\u2_Display/n6193 ,\u2_Display/n6194 ,\u2_Display/n6195 ,\u2_Display/n6196 ,\u2_Display/n6197 ,\u2_Display/n6198 ,\u2_Display/n6199 ,\u2_Display/n6200 ,\u2_Display/n6201 ,\u2_Display/n6202 ,\u2_Display/n6203 ,\u2_Display/n6204 ,\u2_Display/n6205 ,\u2_Display/n6206 }),
    .i1(32'b00001010000000000000000000000000),
    .o(\u2_Display/n5049 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt159  (
    .ci(1'b0),
    .i0({\u2_Display/n6210 ,\u2_Display/n6211 ,\u2_Display/n6212 ,\u2_Display/n6213 ,\u2_Display/n6214 ,\u2_Display/n6215 ,\u2_Display/n6216 ,\u2_Display/n6217 ,\u2_Display/n6218 ,\u2_Display/n6219 ,\u2_Display/n6220 ,\u2_Display/n6221 ,\u2_Display/n6222 ,\u2_Display/n6223 ,\u2_Display/n6224 ,\u2_Display/n6225 ,\u2_Display/n6226 ,\u2_Display/n6227 ,\u2_Display/n6228 ,\u2_Display/n6229 ,\u2_Display/n6230 ,\u2_Display/n6231 ,\u2_Display/n6232 ,\u2_Display/n6233 ,\u2_Display/n6234 ,\u2_Display/n6235 ,\u2_Display/n6236 ,\u2_Display/n6237 ,\u2_Display/n6238 ,\u2_Display/n6239 ,\u2_Display/n6240 ,\u2_Display/n6241 }),
    .i1(32'b00000101000000000000000000000000),
    .o(\u2_Display/n5084 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt160  (
    .ci(1'b0),
    .i0({\u2_Display/n6245 ,\u2_Display/n6246 ,\u2_Display/n6247 ,\u2_Display/n6248 ,\u2_Display/n6249 ,\u2_Display/n6250 ,\u2_Display/n6251 ,\u2_Display/n6252 ,\u2_Display/n6253 ,\u2_Display/n6254 ,\u2_Display/n6255 ,\u2_Display/n6256 ,\u2_Display/n6257 ,\u2_Display/n6258 ,\u2_Display/n6259 ,\u2_Display/n6260 ,\u2_Display/n6261 ,\u2_Display/n6262 ,\u2_Display/n6263 ,\u2_Display/n6264 ,\u2_Display/n6265 ,\u2_Display/n6266 ,\u2_Display/n6267 ,\u2_Display/n6268 ,\u2_Display/n6269 ,\u2_Display/n6270 ,\u2_Display/n6271 ,\u2_Display/n6272 ,\u2_Display/n6273 ,\u2_Display/n6274 ,\u2_Display/n6275 ,\u2_Display/n6276 }),
    .i1(32'b00000010100000000000000000000000),
    .o(\u2_Display/n5119 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt161  (
    .ci(1'b0),
    .i0({\u2_Display/n6280 ,\u2_Display/n6281 ,\u2_Display/n6282 ,\u2_Display/n6283 ,\u2_Display/n6284 ,\u2_Display/n6285 ,\u2_Display/n6286 ,\u2_Display/n6287 ,\u2_Display/n6288 ,\u2_Display/n6289 ,\u2_Display/n6290 ,\u2_Display/n6291 ,\u2_Display/n6292 ,\u2_Display/n6293 ,\u2_Display/n6294 ,\u2_Display/n6295 ,\u2_Display/n6296 ,\u2_Display/n6297 ,\u2_Display/n6298 ,\u2_Display/n6299 ,\u2_Display/n6300 ,\u2_Display/n6301 ,\u2_Display/n6302 ,\u2_Display/n6303 ,\u2_Display/n6304 ,\u2_Display/n6305 ,\u2_Display/n6306 ,\u2_Display/n6307 ,\u2_Display/n6308 ,\u2_Display/n6309 ,\u2_Display/n6310 ,\u2_Display/n6311 }),
    .i1(32'b00000001010000000000000000000000),
    .o(\u2_Display/n5154 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt162  (
    .ci(1'b0),
    .i0({\u2_Display/n6315 ,\u2_Display/n6316 ,\u2_Display/n6317 ,\u2_Display/n6318 ,\u2_Display/n6319 ,\u2_Display/n6320 ,\u2_Display/n6321 ,\u2_Display/n6322 ,\u2_Display/n6323 ,\u2_Display/n6324 ,\u2_Display/n6325 ,\u2_Display/n6326 ,\u2_Display/n6327 ,\u2_Display/n6328 ,\u2_Display/n6329 ,\u2_Display/n6330 ,\u2_Display/n6331 ,\u2_Display/n6332 ,\u2_Display/n6333 ,\u2_Display/n6334 ,\u2_Display/n6335 ,\u2_Display/n6336 ,\u2_Display/n6337 ,\u2_Display/n6338 ,\u2_Display/n6339 ,\u2_Display/n6340 ,\u2_Display/n6341 ,\u2_Display/n6342 ,\u2_Display/n6343 ,\u2_Display/n6344 ,\u2_Display/n6345 ,\u2_Display/n6346 }),
    .i1(32'b00000000101000000000000000000000),
    .o(\u2_Display/n5189 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt163  (
    .ci(1'b0),
    .i0({\u2_Display/n6350 ,\u2_Display/n6351 ,\u2_Display/n6352 ,\u2_Display/n6353 ,\u2_Display/n5196 ,\u2_Display/n5197 ,\u2_Display/n5198 ,\u2_Display/n5199 ,\u2_Display/n5200 ,\u2_Display/n5201 ,\u2_Display/n5202 ,\u2_Display/n5203 ,\u2_Display/n5204 ,\u2_Display/n5205 ,\u2_Display/n5206 ,\u2_Display/n5207 ,\u2_Display/n5208 ,\u2_Display/n5209 ,\u2_Display/n5210 ,\u2_Display/n5211 ,\u2_Display/n5212 ,\u2_Display/n5213 ,\u2_Display/n5214 ,\u2_Display/n5215 ,\u2_Display/n5216 ,\u2_Display/n5217 ,\u2_Display/n5218 ,\u2_Display/n5219 ,\u2_Display/n5220 ,\u2_Display/n5221 ,\u2_Display/n5222 ,\u2_Display/n5223 }),
    .i1(32'b00000000010100000000000000000000),
    .o(\u2_Display/n5224 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt164  (
    .ci(1'b0),
    .i0({\u2_Display/n5227 ,\u2_Display/n5228 ,\u2_Display/n5229 ,\u2_Display/n5230 ,\u2_Display/n5231 ,\u2_Display/n5232 ,\u2_Display/n5233 ,\u2_Display/n5234 ,\u2_Display/n5235 ,\u2_Display/n5236 ,\u2_Display/n5237 ,\u2_Display/n5238 ,\u2_Display/n5239 ,\u2_Display/n5240 ,\u2_Display/n5241 ,\u2_Display/n5242 ,\u2_Display/n5243 ,\u2_Display/n5244 ,\u2_Display/n5245 ,\u2_Display/n5246 ,\u2_Display/n5247 ,\u2_Display/n5248 ,\u2_Display/n5249 ,\u2_Display/n5250 ,\u2_Display/n5251 ,\u2_Display/n5252 ,\u2_Display/n5253 ,\u2_Display/n5254 ,\u2_Display/n5255 ,\u2_Display/n5256 ,\u2_Display/n5257 ,\u2_Display/n5258 }),
    .i1(32'b00000000001010000000000000000000),
    .o(\u2_Display/n5259 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt165  (
    .ci(1'b0),
    .i0({\u2_Display/n5262 ,\u2_Display/n5263 ,\u2_Display/n5264 ,\u2_Display/n5265 ,\u2_Display/n5266 ,\u2_Display/n5267 ,\u2_Display/n5268 ,\u2_Display/n5269 ,\u2_Display/n5270 ,\u2_Display/n5271 ,\u2_Display/n5272 ,\u2_Display/n5273 ,\u2_Display/n5274 ,\u2_Display/n5275 ,\u2_Display/n5276 ,\u2_Display/n5277 ,\u2_Display/n5278 ,\u2_Display/n5279 ,\u2_Display/n5280 ,\u2_Display/n5281 ,\u2_Display/n5282 ,\u2_Display/n5283 ,\u2_Display/n5284 ,\u2_Display/n5285 ,\u2_Display/n5286 ,\u2_Display/n5287 ,\u2_Display/n5288 ,\u2_Display/n5289 ,\u2_Display/n5290 ,\u2_Display/n5291 ,\u2_Display/n5292 ,\u2_Display/n5293 }),
    .i1(32'b00000000000101000000000000000000),
    .o(\u2_Display/n5294 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt166  (
    .ci(1'b0),
    .i0({\u2_Display/n5297 ,\u2_Display/n5298 ,\u2_Display/n5299 ,\u2_Display/n5300 ,\u2_Display/n5301 ,\u2_Display/n5302 ,\u2_Display/n5303 ,\u2_Display/n5304 ,\u2_Display/n5305 ,\u2_Display/n5306 ,\u2_Display/n5307 ,\u2_Display/n5308 ,\u2_Display/n5309 ,\u2_Display/n5310 ,\u2_Display/n5311 ,\u2_Display/n5312 ,\u2_Display/n5313 ,\u2_Display/n5314 ,\u2_Display/n5315 ,\u2_Display/n5316 ,\u2_Display/n5317 ,\u2_Display/n5318 ,\u2_Display/n5319 ,\u2_Display/n5320 ,\u2_Display/n5321 ,\u2_Display/n5322 ,\u2_Display/n5323 ,\u2_Display/n5324 ,\u2_Display/n5325 ,\u2_Display/n5326 ,\u2_Display/n5327 ,\u2_Display/n5328 }),
    .i1(32'b00000000000010100000000000000000),
    .o(\u2_Display/n5329 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt167  (
    .ci(1'b0),
    .i0({\u2_Display/n5332 ,\u2_Display/n5333 ,\u2_Display/n5334 ,\u2_Display/n5335 ,\u2_Display/n5336 ,\u2_Display/n5337 ,\u2_Display/n5338 ,\u2_Display/n5339 ,\u2_Display/n5340 ,\u2_Display/n5341 ,\u2_Display/n5342 ,\u2_Display/n5343 ,\u2_Display/n5344 ,\u2_Display/n5345 ,\u2_Display/n5346 ,\u2_Display/n5347 ,\u2_Display/n5348 ,\u2_Display/n5349 ,\u2_Display/n5350 ,\u2_Display/n5351 ,\u2_Display/n5352 ,\u2_Display/n5353 ,\u2_Display/n5354 ,\u2_Display/n5355 ,\u2_Display/n5356 ,\u2_Display/n5357 ,\u2_Display/n5358 ,\u2_Display/n5359 ,\u2_Display/n5360 ,\u2_Display/n5361 ,\u2_Display/n5362 ,\u2_Display/n5363 }),
    .i1(32'b00000000000001010000000000000000),
    .o(\u2_Display/n5364 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt168  (
    .ci(1'b0),
    .i0({\u2_Display/n5367 ,\u2_Display/n5368 ,\u2_Display/n5369 ,\u2_Display/n5370 ,\u2_Display/n5371 ,\u2_Display/n5372 ,\u2_Display/n5373 ,\u2_Display/n5374 ,\u2_Display/n5375 ,\u2_Display/n5376 ,\u2_Display/n5377 ,\u2_Display/n5378 ,\u2_Display/n5379 ,\u2_Display/n5380 ,\u2_Display/n5381 ,\u2_Display/n5382 ,\u2_Display/n5383 ,\u2_Display/n5384 ,\u2_Display/n5385 ,\u2_Display/n5386 ,\u2_Display/n5387 ,\u2_Display/n5388 ,\u2_Display/n5389 ,\u2_Display/n5390 ,\u2_Display/n5391 ,\u2_Display/n5392 ,\u2_Display/n5393 ,\u2_Display/n5394 ,\u2_Display/n5395 ,\u2_Display/n5396 ,\u2_Display/n5397 ,\u2_Display/n5398 }),
    .i1(32'b00000000000000101000000000000000),
    .o(\u2_Display/n5399 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt169  (
    .ci(1'b0),
    .i0({\u2_Display/n5402 ,\u2_Display/n5403 ,\u2_Display/n5404 ,\u2_Display/n5405 ,\u2_Display/n5406 ,\u2_Display/n5407 ,\u2_Display/n5408 ,\u2_Display/n5409 ,\u2_Display/n5410 ,\u2_Display/n5411 ,\u2_Display/n5412 ,\u2_Display/n5413 ,\u2_Display/n5414 ,\u2_Display/n5415 ,\u2_Display/n5416 ,\u2_Display/n5417 ,\u2_Display/n5418 ,\u2_Display/n5419 ,\u2_Display/n5420 ,\u2_Display/n5421 ,\u2_Display/n5422 ,\u2_Display/n5423 ,\u2_Display/n5424 ,\u2_Display/n5425 ,\u2_Display/n5426 ,\u2_Display/n5427 ,\u2_Display/n5428 ,\u2_Display/n5429 ,\u2_Display/n5430 ,\u2_Display/n5431 ,\u2_Display/n5432 ,\u2_Display/n5433 }),
    .i1(32'b00000000000000010100000000000000),
    .o(\u2_Display/n5434 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt170  (
    .ci(1'b0),
    .i0({\u2_Display/n5437 ,\u2_Display/n5438 ,\u2_Display/n5439 ,\u2_Display/n5440 ,\u2_Display/n5441 ,\u2_Display/n5442 ,\u2_Display/n5443 ,\u2_Display/n5444 ,\u2_Display/n5445 ,\u2_Display/n5446 ,\u2_Display/n5447 ,\u2_Display/n5448 ,\u2_Display/n5449 ,\u2_Display/n5450 ,\u2_Display/n5451 ,\u2_Display/n5452 ,\u2_Display/n5453 ,\u2_Display/n5454 ,\u2_Display/n5455 ,\u2_Display/n5456 ,\u2_Display/n5457 ,\u2_Display/n5458 ,\u2_Display/n5459 ,\u2_Display/n5460 ,\u2_Display/n5461 ,\u2_Display/n5462 ,\u2_Display/n5463 ,\u2_Display/n5464 ,\u2_Display/n5465 ,\u2_Display/n5466 ,\u2_Display/n5467 ,\u2_Display/n5468 }),
    .i1(32'b00000000000000001010000000000000),
    .o(\u2_Display/n5469 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt171  (
    .ci(1'b0),
    .i0({\u2_Display/n5472 ,\u2_Display/n5473 ,\u2_Display/n5474 ,\u2_Display/n5475 ,\u2_Display/n5476 ,\u2_Display/n5477 ,\u2_Display/n5478 ,\u2_Display/n5479 ,\u2_Display/n5480 ,\u2_Display/n5481 ,\u2_Display/n5482 ,\u2_Display/n5483 ,\u2_Display/n5484 ,\u2_Display/n5485 ,\u2_Display/n5486 ,\u2_Display/n5487 ,\u2_Display/n5488 ,\u2_Display/n5489 ,\u2_Display/n5490 ,\u2_Display/n5491 ,\u2_Display/n5492 ,\u2_Display/n5493 ,\u2_Display/n5494 ,\u2_Display/n5495 ,\u2_Display/n5496 ,\u2_Display/n5497 ,\u2_Display/n5498 ,\u2_Display/n5499 ,\u2_Display/n5500 ,\u2_Display/n5501 ,\u2_Display/n5502 ,\u2_Display/n5503 }),
    .i1(32'b00000000000000000101000000000000),
    .o(\u2_Display/n5504 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt172  (
    .ci(1'b0),
    .i0({\u2_Display/n5507 ,\u2_Display/n5508 ,\u2_Display/n5509 ,\u2_Display/n5510 ,\u2_Display/n5511 ,\u2_Display/n5512 ,\u2_Display/n5513 ,\u2_Display/n5514 ,\u2_Display/n5515 ,\u2_Display/n5516 ,\u2_Display/n5517 ,\u2_Display/n5518 ,\u2_Display/n5519 ,\u2_Display/n5520 ,\u2_Display/n5521 ,\u2_Display/n5522 ,\u2_Display/n5523 ,\u2_Display/n5524 ,\u2_Display/n5525 ,\u2_Display/n5526 ,\u2_Display/n5527 ,\u2_Display/n5528 ,\u2_Display/n5529 ,\u2_Display/n5530 ,\u2_Display/n5531 ,\u2_Display/n5532 ,\u2_Display/n5533 ,\u2_Display/n5534 ,\u2_Display/n5535 ,\u2_Display/n5536 ,\u2_Display/n5537 ,\u2_Display/n5538 }),
    .i1(32'b00000000000000000010100000000000),
    .o(\u2_Display/n5539 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt173  (
    .ci(1'b0),
    .i0({\u2_Display/n5542 ,\u2_Display/n5543 ,\u2_Display/n5544 ,\u2_Display/n5545 ,\u2_Display/n5546 ,\u2_Display/n5547 ,\u2_Display/n5548 ,\u2_Display/n5549 ,\u2_Display/n5550 ,\u2_Display/n5551 ,\u2_Display/n5552 ,\u2_Display/n5553 ,\u2_Display/n5554 ,\u2_Display/n5555 ,\u2_Display/n5556 ,\u2_Display/n5557 ,\u2_Display/n5558 ,\u2_Display/n5559 ,\u2_Display/n5560 ,\u2_Display/n5561 ,\u2_Display/n5562 ,\u2_Display/n5563 ,\u2_Display/n5564 ,\u2_Display/n5565 ,\u2_Display/n5566 ,\u2_Display/n5567 ,\u2_Display/n5568 ,\u2_Display/n5569 ,\u2_Display/n5570 ,\u2_Display/n5571 ,\u2_Display/n5572 ,\u2_Display/n5573 }),
    .i1(32'b00000000000000000001010000000000),
    .o(\u2_Display/n5574 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt174  (
    .ci(1'b0),
    .i0({\u2_Display/n5577 ,\u2_Display/n5578 ,\u2_Display/n5579 ,\u2_Display/n5580 ,\u2_Display/n5581 ,\u2_Display/n5582 ,\u2_Display/n5583 ,\u2_Display/n5584 ,\u2_Display/n5585 ,\u2_Display/n5586 ,\u2_Display/n5587 ,\u2_Display/n5588 ,\u2_Display/n5589 ,\u2_Display/n5590 ,\u2_Display/n5591 ,\u2_Display/n5592 ,\u2_Display/n5593 ,\u2_Display/n5594 ,\u2_Display/n5595 ,\u2_Display/n5596 ,\u2_Display/n5597 ,\u2_Display/n5598 ,\u2_Display/n5599 ,\u2_Display/n5600 ,\u2_Display/n5601 ,\u2_Display/n5602 ,\u2_Display/n5603 ,\u2_Display/n5604 ,\u2_Display/n5605 ,\u2_Display/n5606 ,\u2_Display/n5607 ,\u2_Display/n5608 }),
    .i1(32'b00000000000000000000101000000000),
    .o(\u2_Display/n5609 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt175  (
    .ci(1'b0),
    .i0({\u2_Display/n5612 ,\u2_Display/n5613 ,\u2_Display/n5614 ,\u2_Display/n5615 ,\u2_Display/n5616 ,\u2_Display/n5617 ,\u2_Display/n5618 ,\u2_Display/n5619 ,\u2_Display/n5620 ,\u2_Display/n5621 ,\u2_Display/n5622 ,\u2_Display/n5623 ,\u2_Display/n5624 ,\u2_Display/n5625 ,\u2_Display/n5626 ,\u2_Display/n5627 ,\u2_Display/n5628 ,\u2_Display/n5629 ,\u2_Display/n5630 ,\u2_Display/n5631 ,\u2_Display/n5632 ,\u2_Display/n5633 ,\u2_Display/n5634 ,\u2_Display/n5635 ,\u2_Display/n5636 ,\u2_Display/n5637 ,\u2_Display/n5638 ,\u2_Display/n5639 ,\u2_Display/n5640 ,\u2_Display/n5641 ,\u2_Display/n5642 ,\u2_Display/n5643 }),
    .i1(32'b00000000000000000000010100000000),
    .o(\u2_Display/n5644 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt176  (
    .ci(1'b0),
    .i0({\u2_Display/n5647 ,\u2_Display/n5648 ,\u2_Display/n5649 ,\u2_Display/n5650 ,\u2_Display/n5651 ,\u2_Display/n5652 ,\u2_Display/n5653 ,\u2_Display/n5654 ,\u2_Display/n5655 ,\u2_Display/n5656 ,\u2_Display/n5657 ,\u2_Display/n5658 ,\u2_Display/n5659 ,\u2_Display/n5660 ,\u2_Display/n5661 ,\u2_Display/n5662 ,\u2_Display/n5663 ,\u2_Display/n5664 ,\u2_Display/n5665 ,\u2_Display/n5666 ,\u2_Display/n5667 ,\u2_Display/n5668 ,\u2_Display/n5669 ,\u2_Display/n5670 ,\u2_Display/n5671 ,\u2_Display/n5672 ,\u2_Display/n5673 ,\u2_Display/n5674 ,\u2_Display/n5675 ,\u2_Display/n5676 ,\u2_Display/n5677 ,\u2_Display/n5678 }),
    .i1(32'b00000000000000000000001010000000),
    .o(\u2_Display/n5679 ));  // source/rtl/Display.v(179)
  lt_u32_u32 \u2_Display/lt22  (
    .ci(1'b0),
    .i0(\u2_Display/counta ),
    .i1(32'b11111010000000000000000000000000),
    .o(\u2_Display/n417 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt23  (
    .ci(1'b0),
    .i0({\u2_Display/n420 ,\u2_Display/n421 ,\u2_Display/n422 ,\u2_Display/n423 ,\u2_Display/n424 ,\u2_Display/n425 ,\u2_Display/n426 ,\u2_Display/n427 ,\u2_Display/n428 ,\u2_Display/n429 ,\u2_Display/n430 ,\u2_Display/n431 ,\u2_Display/n432 ,\u2_Display/n433 ,\u2_Display/n434 ,\u2_Display/n435 ,\u2_Display/n436 ,\u2_Display/n437 ,\u2_Display/n438 ,\u2_Display/n439 ,\u2_Display/n440 ,\u2_Display/n441 ,\u2_Display/n442 ,\u2_Display/n443 ,\u2_Display/n444 ,\u2_Display/n445 ,\u2_Display/n446 ,\u2_Display/n447 ,\u2_Display/n448 ,\u2_Display/n449 ,\u2_Display/n450 ,\u2_Display/n451 }),
    .i1(32'b01111101000000000000000000000000),
    .o(\u2_Display/n452 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt24  (
    .ci(1'b0),
    .i0({\u2_Display/n455 ,\u2_Display/n456 ,\u2_Display/n457 ,\u2_Display/n458 ,\u2_Display/n459 ,\u2_Display/n460 ,\u2_Display/n461 ,\u2_Display/n462 ,\u2_Display/n463 ,\u2_Display/n464 ,\u2_Display/n465 ,\u2_Display/n466 ,\u2_Display/n467 ,\u2_Display/n468 ,\u2_Display/n469 ,\u2_Display/n470 ,\u2_Display/n471 ,\u2_Display/n472 ,\u2_Display/n473 ,\u2_Display/n474 ,\u2_Display/n475 ,\u2_Display/n476 ,\u2_Display/n477 ,\u2_Display/n478 ,\u2_Display/n479 ,\u2_Display/n480 ,\u2_Display/n481 ,\u2_Display/n482 ,\u2_Display/n483 ,\u2_Display/n484 ,\u2_Display/n485 ,\u2_Display/n486 }),
    .i1(32'b00111110100000000000000000000000),
    .o(\u2_Display/n487 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt25  (
    .ci(1'b0),
    .i0({\u2_Display/n490 ,\u2_Display/n491 ,\u2_Display/n492 ,\u2_Display/n493 ,\u2_Display/n494 ,\u2_Display/n495 ,\u2_Display/n496 ,\u2_Display/n497 ,\u2_Display/n498 ,\u2_Display/n499 ,\u2_Display/n500 ,\u2_Display/n501 ,\u2_Display/n502 ,\u2_Display/n503 ,\u2_Display/n504 ,\u2_Display/n505 ,\u2_Display/n506 ,\u2_Display/n507 ,\u2_Display/n508 ,\u2_Display/n509 ,\u2_Display/n510 ,\u2_Display/n511 ,\u2_Display/n512 ,\u2_Display/n513 ,\u2_Display/n514 ,\u2_Display/n515 ,\u2_Display/n516 ,\u2_Display/n517 ,\u2_Display/n518 ,\u2_Display/n519 ,\u2_Display/n520 ,\u2_Display/n521 }),
    .i1(32'b00011111010000000000000000000000),
    .o(\u2_Display/n522 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt26  (
    .ci(1'b0),
    .i0({\u2_Display/n525 ,\u2_Display/n526 ,\u2_Display/n527 ,\u2_Display/n528 ,\u2_Display/n529 ,\u2_Display/n530 ,\u2_Display/n531 ,\u2_Display/n532 ,\u2_Display/n533 ,\u2_Display/n534 ,\u2_Display/n535 ,\u2_Display/n536 ,\u2_Display/n537 ,\u2_Display/n538 ,\u2_Display/n539 ,\u2_Display/n540 ,\u2_Display/n541 ,\u2_Display/n542 ,\u2_Display/n543 ,\u2_Display/n544 ,\u2_Display/n545 ,\u2_Display/n546 ,\u2_Display/n547 ,\u2_Display/n548 ,\u2_Display/n549 ,\u2_Display/n550 ,\u2_Display/n551 ,\u2_Display/n552 ,\u2_Display/n553 ,\u2_Display/n554 ,\u2_Display/n555 ,\u2_Display/n556 }),
    .i1(32'b00001111101000000000000000000000),
    .o(\u2_Display/n557 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt27  (
    .ci(1'b0),
    .i0({\u2_Display/n560 ,\u2_Display/n561 ,\u2_Display/n562 ,\u2_Display/n563 ,\u2_Display/n564 ,\u2_Display/n565 ,\u2_Display/n566 ,\u2_Display/n567 ,\u2_Display/n568 ,\u2_Display/n569 ,\u2_Display/n570 ,\u2_Display/n571 ,\u2_Display/n572 ,\u2_Display/n573 ,\u2_Display/n574 ,\u2_Display/n575 ,\u2_Display/n576 ,\u2_Display/n577 ,\u2_Display/n578 ,\u2_Display/n579 ,\u2_Display/n580 ,\u2_Display/n581 ,\u2_Display/n582 ,\u2_Display/n583 ,\u2_Display/n584 ,\u2_Display/n585 ,\u2_Display/n586 ,\u2_Display/n587 ,\u2_Display/n588 ,\u2_Display/n589 ,\u2_Display/n590 ,\u2_Display/n591 }),
    .i1(32'b00000111110100000000000000000000),
    .o(\u2_Display/n592 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt28  (
    .ci(1'b0),
    .i0({\u2_Display/n595 ,\u2_Display/n596 ,\u2_Display/n597 ,\u2_Display/n598 ,\u2_Display/n599 ,\u2_Display/n600 ,\u2_Display/n601 ,\u2_Display/n602 ,\u2_Display/n603 ,\u2_Display/n604 ,\u2_Display/n605 ,\u2_Display/n606 ,\u2_Display/n607 ,\u2_Display/n608 ,\u2_Display/n609 ,\u2_Display/n610 ,\u2_Display/n611 ,\u2_Display/n612 ,\u2_Display/n613 ,\u2_Display/n614 ,\u2_Display/n615 ,\u2_Display/n616 ,\u2_Display/n617 ,\u2_Display/n618 ,\u2_Display/n619 ,\u2_Display/n620 ,\u2_Display/n621 ,\u2_Display/n622 ,\u2_Display/n623 ,\u2_Display/n624 ,\u2_Display/n625 ,\u2_Display/n626 }),
    .i1(32'b00000011111010000000000000000000),
    .o(\u2_Display/n627 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt29  (
    .ci(1'b0),
    .i0({\u2_Display/n630 ,\u2_Display/n631 ,\u2_Display/n632 ,\u2_Display/n633 ,\u2_Display/n634 ,\u2_Display/n635 ,\u2_Display/n636 ,\u2_Display/n637 ,\u2_Display/n638 ,\u2_Display/n639 ,\u2_Display/n640 ,\u2_Display/n641 ,\u2_Display/n642 ,\u2_Display/n643 ,\u2_Display/n644 ,\u2_Display/n645 ,\u2_Display/n646 ,\u2_Display/n647 ,\u2_Display/n648 ,\u2_Display/n649 ,\u2_Display/n650 ,\u2_Display/n651 ,\u2_Display/n652 ,\u2_Display/n653 ,\u2_Display/n654 ,\u2_Display/n655 ,\u2_Display/n656 ,\u2_Display/n657 ,\u2_Display/n658 ,\u2_Display/n659 ,\u2_Display/n660 ,\u2_Display/n661 }),
    .i1(32'b00000001111101000000000000000000),
    .o(\u2_Display/n662 ));  // source/rtl/Display.v(230)
  lt_u12_u12 \u2_Display/lt2_2  (
    .ci(1'b0),
    .i0(lcd_ypos),
    .i1({2'b01,\u2_Display/j [9:0]}),
    .o(\u2_Display/n48 ));  // source/rtl/Display.v(165)
  lt_u12_u12 \u2_Display/lt3  (
    .ci(1'b0),
    .i0({2'b00,\u2_Display/j [9:0]}),
    .i1(lcd_ypos),
    .o(\u2_Display/n50 ));  // source/rtl/Display.v(165)
  lt_u32_u32 \u2_Display/lt30  (
    .ci(1'b0),
    .i0({\u2_Display/n665 ,\u2_Display/n666 ,\u2_Display/n667 ,\u2_Display/n668 ,\u2_Display/n669 ,\u2_Display/n670 ,\u2_Display/n671 ,\u2_Display/n672 ,\u2_Display/n673 ,\u2_Display/n674 ,\u2_Display/n675 ,\u2_Display/n676 ,\u2_Display/n677 ,\u2_Display/n678 ,\u2_Display/n679 ,\u2_Display/n680 ,\u2_Display/n681 ,\u2_Display/n682 ,\u2_Display/n683 ,\u2_Display/n684 ,\u2_Display/n685 ,\u2_Display/n686 ,\u2_Display/n687 ,\u2_Display/n688 ,\u2_Display/n689 ,\u2_Display/n690 ,\u2_Display/n691 ,\u2_Display/n692 ,\u2_Display/n693 ,\u2_Display/n694 ,\u2_Display/n695 ,\u2_Display/n696 }),
    .i1(32'b00000000111110100000000000000000),
    .o(\u2_Display/n697 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt31  (
    .ci(1'b0),
    .i0({\u2_Display/n700 ,\u2_Display/n701 ,\u2_Display/n702 ,\u2_Display/n703 ,\u2_Display/n704 ,\u2_Display/n705 ,\u2_Display/n706 ,\u2_Display/n707 ,\u2_Display/n708 ,\u2_Display/n709 ,\u2_Display/n710 ,\u2_Display/n711 ,\u2_Display/n712 ,\u2_Display/n713 ,\u2_Display/n714 ,\u2_Display/n715 ,\u2_Display/n716 ,\u2_Display/n717 ,\u2_Display/n718 ,\u2_Display/n719 ,\u2_Display/n720 ,\u2_Display/n721 ,\u2_Display/n722 ,\u2_Display/n723 ,\u2_Display/n724 ,\u2_Display/n725 ,\u2_Display/n726 ,\u2_Display/n727 ,\u2_Display/n728 ,\u2_Display/n729 ,\u2_Display/n730 ,\u2_Display/n731 }),
    .i1(32'b00000000011111010000000000000000),
    .o(\u2_Display/n732 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt32  (
    .ci(1'b0),
    .i0({\u2_Display/n735 ,\u2_Display/n736 ,\u2_Display/n737 ,\u2_Display/n738 ,\u2_Display/n739 ,\u2_Display/n740 ,\u2_Display/n741 ,\u2_Display/n742 ,\u2_Display/n743 ,\u2_Display/n744 ,\u2_Display/n745 ,\u2_Display/n746 ,\u2_Display/n747 ,\u2_Display/n748 ,\u2_Display/n749 ,\u2_Display/n750 ,\u2_Display/n751 ,\u2_Display/n752 ,\u2_Display/n753 ,\u2_Display/n754 ,\u2_Display/n755 ,\u2_Display/n756 ,\u2_Display/n757 ,\u2_Display/n758 ,\u2_Display/n759 ,\u2_Display/n760 ,\u2_Display/n761 ,\u2_Display/n762 ,\u2_Display/n763 ,\u2_Display/n764 ,\u2_Display/n765 ,\u2_Display/n766 }),
    .i1(32'b00000000001111101000000000000000),
    .o(\u2_Display/n767 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt33  (
    .ci(1'b0),
    .i0({\u2_Display/n770 ,\u2_Display/n771 ,\u2_Display/n772 ,\u2_Display/n773 ,\u2_Display/n774 ,\u2_Display/n775 ,\u2_Display/n776 ,\u2_Display/n777 ,\u2_Display/n778 ,\u2_Display/n779 ,\u2_Display/n780 ,\u2_Display/n781 ,\u2_Display/n782 ,\u2_Display/n783 ,\u2_Display/n784 ,\u2_Display/n785 ,\u2_Display/n786 ,\u2_Display/n787 ,\u2_Display/n788 ,\u2_Display/n789 ,\u2_Display/n790 ,\u2_Display/n791 ,\u2_Display/n792 ,\u2_Display/n793 ,\u2_Display/n794 ,\u2_Display/n795 ,\u2_Display/n796 ,\u2_Display/n797 ,\u2_Display/n798 ,\u2_Display/n799 ,\u2_Display/n800 ,\u2_Display/n801 }),
    .i1(32'b00000000000111110100000000000000),
    .o(\u2_Display/n802 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt34  (
    .ci(1'b0),
    .i0({\u2_Display/n805 ,\u2_Display/n806 ,\u2_Display/n807 ,\u2_Display/n808 ,\u2_Display/n809 ,\u2_Display/n810 ,\u2_Display/n811 ,\u2_Display/n812 ,\u2_Display/n813 ,\u2_Display/n814 ,\u2_Display/n815 ,\u2_Display/n816 ,\u2_Display/n817 ,\u2_Display/n818 ,\u2_Display/n819 ,\u2_Display/n820 ,\u2_Display/n821 ,\u2_Display/n822 ,\u2_Display/n823 ,\u2_Display/n824 ,\u2_Display/n825 ,\u2_Display/n826 ,\u2_Display/n827 ,\u2_Display/n828 ,\u2_Display/n829 ,\u2_Display/n830 ,\u2_Display/n831 ,\u2_Display/n832 ,\u2_Display/n833 ,\u2_Display/n834 ,\u2_Display/n835 ,\u2_Display/n836 }),
    .i1(32'b00000000000011111010000000000000),
    .o(\u2_Display/n837 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt35  (
    .ci(1'b0),
    .i0({\u2_Display/n840 ,\u2_Display/n841 ,\u2_Display/n842 ,\u2_Display/n843 ,\u2_Display/n844 ,\u2_Display/n845 ,\u2_Display/n846 ,\u2_Display/n847 ,\u2_Display/n848 ,\u2_Display/n849 ,\u2_Display/n850 ,\u2_Display/n851 ,\u2_Display/n852 ,\u2_Display/n853 ,\u2_Display/n854 ,\u2_Display/n855 ,\u2_Display/n856 ,\u2_Display/n857 ,\u2_Display/n858 ,\u2_Display/n859 ,\u2_Display/n860 ,\u2_Display/n861 ,\u2_Display/n862 ,\u2_Display/n863 ,\u2_Display/n864 ,\u2_Display/n865 ,\u2_Display/n866 ,\u2_Display/n867 ,\u2_Display/n868 ,\u2_Display/n869 ,\u2_Display/n870 ,\u2_Display/n871 }),
    .i1(32'b00000000000001111101000000000000),
    .o(\u2_Display/n872 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt36  (
    .ci(1'b0),
    .i0({\u2_Display/n875 ,\u2_Display/n876 ,\u2_Display/n877 ,\u2_Display/n878 ,\u2_Display/n879 ,\u2_Display/n880 ,\u2_Display/n881 ,\u2_Display/n882 ,\u2_Display/n883 ,\u2_Display/n884 ,\u2_Display/n885 ,\u2_Display/n886 ,\u2_Display/n887 ,\u2_Display/n888 ,\u2_Display/n889 ,\u2_Display/n890 ,\u2_Display/n891 ,\u2_Display/n892 ,\u2_Display/n893 ,\u2_Display/n894 ,\u2_Display/n895 ,\u2_Display/n896 ,\u2_Display/n897 ,\u2_Display/n898 ,\u2_Display/n899 ,\u2_Display/n900 ,\u2_Display/n901 ,\u2_Display/n902 ,\u2_Display/n903 ,\u2_Display/n904 ,\u2_Display/n905 ,\u2_Display/n906 }),
    .i1(32'b00000000000000111110100000000000),
    .o(\u2_Display/n907 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt37  (
    .ci(1'b0),
    .i0({\u2_Display/n910 ,\u2_Display/n911 ,\u2_Display/n912 ,\u2_Display/n913 ,\u2_Display/n914 ,\u2_Display/n915 ,\u2_Display/n916 ,\u2_Display/n917 ,\u2_Display/n918 ,\u2_Display/n919 ,\u2_Display/n920 ,\u2_Display/n921 ,\u2_Display/n922 ,\u2_Display/n923 ,\u2_Display/n924 ,\u2_Display/n925 ,\u2_Display/n926 ,\u2_Display/n927 ,\u2_Display/n928 ,\u2_Display/n929 ,\u2_Display/n930 ,\u2_Display/n931 ,\u2_Display/n932 ,\u2_Display/n933 ,\u2_Display/n934 ,\u2_Display/n935 ,\u2_Display/n936 ,\u2_Display/n937 ,\u2_Display/n938 ,\u2_Display/n939 ,\u2_Display/n940 ,\u2_Display/n941 }),
    .i1(32'b00000000000000011111010000000000),
    .o(\u2_Display/n942 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt38  (
    .ci(1'b0),
    .i0({\u2_Display/n945 ,\u2_Display/n946 ,\u2_Display/n947 ,\u2_Display/n948 ,\u2_Display/n949 ,\u2_Display/n950 ,\u2_Display/n951 ,\u2_Display/n952 ,\u2_Display/n953 ,\u2_Display/n954 ,\u2_Display/n955 ,\u2_Display/n956 ,\u2_Display/n957 ,\u2_Display/n958 ,\u2_Display/n959 ,\u2_Display/n960 ,\u2_Display/n961 ,\u2_Display/n962 ,\u2_Display/n963 ,\u2_Display/n964 ,\u2_Display/n965 ,\u2_Display/n966 ,\u2_Display/n967 ,\u2_Display/n968 ,\u2_Display/n969 ,\u2_Display/n970 ,\u2_Display/n971 ,\u2_Display/n972 ,\u2_Display/n973 ,\u2_Display/n974 ,\u2_Display/n975 ,\u2_Display/n976 }),
    .i1(32'b00000000000000001111101000000000),
    .o(\u2_Display/n977 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt39  (
    .ci(1'b0),
    .i0({\u2_Display/n980 ,\u2_Display/n981 ,\u2_Display/n982 ,\u2_Display/n983 ,\u2_Display/n984 ,\u2_Display/n985 ,\u2_Display/n986 ,\u2_Display/n987 ,\u2_Display/n988 ,\u2_Display/n989 ,\u2_Display/n990 ,\u2_Display/n991 ,\u2_Display/n992 ,\u2_Display/n993 ,\u2_Display/n994 ,\u2_Display/n995 ,\u2_Display/n996 ,\u2_Display/n997 ,\u2_Display/n998 ,\u2_Display/n999 ,\u2_Display/n1000 ,\u2_Display/n1001 ,\u2_Display/n1002 ,\u2_Display/n1003 ,\u2_Display/n1004 ,\u2_Display/n1005 ,\u2_Display/n1006 ,\u2_Display/n1007 ,\u2_Display/n1008 ,\u2_Display/n1009 ,\u2_Display/n1010 ,\u2_Display/n1011 }),
    .i1(32'b00000000000000000111110100000000),
    .o(\u2_Display/n1012 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt40  (
    .ci(1'b0),
    .i0({\u2_Display/n1015 ,\u2_Display/n1016 ,\u2_Display/n1017 ,\u2_Display/n1018 ,\u2_Display/n1019 ,\u2_Display/n1020 ,\u2_Display/n1021 ,\u2_Display/n1022 ,\u2_Display/n1023 ,\u2_Display/n1024 ,\u2_Display/n1025 ,\u2_Display/n1026 ,\u2_Display/n1027 ,\u2_Display/n1028 ,\u2_Display/n1029 ,\u2_Display/n1030 ,\u2_Display/n1031 ,\u2_Display/n1032 ,\u2_Display/n1033 ,\u2_Display/n1034 ,\u2_Display/n1035 ,\u2_Display/n1036 ,\u2_Display/n1037 ,\u2_Display/n1038 ,\u2_Display/n1039 ,\u2_Display/n1040 ,\u2_Display/n1041 ,\u2_Display/n1042 ,\u2_Display/n1043 ,\u2_Display/n1044 ,\u2_Display/n1045 ,\u2_Display/n1046 }),
    .i1(32'b00000000000000000011111010000000),
    .o(\u2_Display/n1047 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt41  (
    .ci(1'b0),
    .i0({\u2_Display/n1050 ,\u2_Display/n1051 ,\u2_Display/n1052 ,\u2_Display/n1053 ,\u2_Display/n1054 ,\u2_Display/n1055 ,\u2_Display/n1056 ,\u2_Display/n1057 ,\u2_Display/n1058 ,\u2_Display/n1059 ,\u2_Display/n1060 ,\u2_Display/n1061 ,\u2_Display/n1062 ,\u2_Display/n1063 ,\u2_Display/n1064 ,\u2_Display/n1065 ,\u2_Display/n1066 ,\u2_Display/n1067 ,\u2_Display/n1068 ,\u2_Display/n1069 ,\u2_Display/n1070 ,\u2_Display/n1071 ,\u2_Display/n1072 ,\u2_Display/n1073 ,\u2_Display/n1074 ,\u2_Display/n1075 ,\u2_Display/n1076 ,\u2_Display/n1077 ,\u2_Display/n1078 ,\u2_Display/n1079 ,\u2_Display/n1080 ,\u2_Display/n1081 }),
    .i1(32'b00000000000000000001111101000000),
    .o(\u2_Display/n1082 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt42  (
    .ci(1'b0),
    .i0({\u2_Display/n1085 ,\u2_Display/n1086 ,\u2_Display/n1087 ,\u2_Display/n1088 ,\u2_Display/n1089 ,\u2_Display/n1090 ,\u2_Display/n1091 ,\u2_Display/n1092 ,\u2_Display/n1093 ,\u2_Display/n1094 ,\u2_Display/n1095 ,\u2_Display/n1096 ,\u2_Display/n1097 ,\u2_Display/n1098 ,\u2_Display/n1099 ,\u2_Display/n1100 ,\u2_Display/n1101 ,\u2_Display/n1102 ,\u2_Display/n1103 ,\u2_Display/n1104 ,\u2_Display/n1105 ,\u2_Display/n1106 ,\u2_Display/n1107 ,\u2_Display/n1108 ,\u2_Display/n1109 ,\u2_Display/n1110 ,\u2_Display/n1111 ,\u2_Display/n1112 ,\u2_Display/n1113 ,\u2_Display/n1114 ,\u2_Display/n1115 ,\u2_Display/n1116 }),
    .i1(32'b00000000000000000000111110100000),
    .o(\u2_Display/n1117 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt43  (
    .ci(1'b0),
    .i0({\u2_Display/n1120 ,\u2_Display/n1121 ,\u2_Display/n1122 ,\u2_Display/n1123 ,\u2_Display/n1124 ,\u2_Display/n1125 ,\u2_Display/n1126 ,\u2_Display/n1127 ,\u2_Display/n1128 ,\u2_Display/n1129 ,\u2_Display/n1130 ,\u2_Display/n1131 ,\u2_Display/n1132 ,\u2_Display/n1133 ,\u2_Display/n1134 ,\u2_Display/n1135 ,\u2_Display/n1136 ,\u2_Display/n1137 ,\u2_Display/n1138 ,\u2_Display/n1139 ,\u2_Display/n1140 ,\u2_Display/n1141 ,\u2_Display/n1142 ,\u2_Display/n1143 ,\u2_Display/n1144 ,\u2_Display/n1145 ,\u2_Display/n1146 ,\u2_Display/n1147 ,\u2_Display/n1148 ,\u2_Display/n1149 ,\u2_Display/n1150 ,\u2_Display/n1151 }),
    .i1(32'b00000000000000000000011111010000),
    .o(\u2_Display/n1152 ));  // source/rtl/Display.v(230)
  lt_u32_u32 \u2_Display/lt44  (
    .ci(1'b0),
    .i0({\u2_Display/n1155 ,\u2_Display/n1156 ,\u2_Display/n1157 ,\u2_Display/n1158 ,\u2_Display/n1159 ,\u2_Display/n1160 ,\u2_Display/n1161 ,\u2_Display/n1162 ,\u2_Display/n1163 ,\u2_Display/n1164 ,\u2_Display/n1165 ,\u2_Display/n1166 ,\u2_Display/n1167 ,\u2_Display/n1168 ,\u2_Display/n1169 ,\u2_Display/n1170 ,\u2_Display/n1171 ,\u2_Display/n1172 ,\u2_Display/n1173 ,\u2_Display/n1174 ,\u2_Display/n1175 ,\u2_Display/n1176 ,\u2_Display/n1177 ,\u2_Display/n1178 ,\u2_Display/n1179 ,\u2_Display/n1180 ,\u2_Display/n1181 ,\u2_Display/n1182 ,\u2_Display/n1183 ,\u2_Display/n1184 ,\u2_Display/n1185 ,\u2_Display/n1186 }),
    .i1(32'b00000000000000000000001111101000),
    .o(\u2_Display/n1187 ));  // source/rtl/Display.v(230)
  lt_u12_u12 \u2_Display/lt4_2  (
    .ci(1'b0),
    .i0(lcd_xpos),
    .i1({\u2_Display/add4_2_co ,\u2_Display/n94 [3:0],\u2_Display/i [6:0]}),
    .o(\u2_Display/n95 ));  // source/rtl/Display.v(181)
  lt_u32_u32 \u2_Display/lt55  (
    .ci(1'b0),
    .i0(\u2_Display/counta ),
    .i1(32'b11100001000000000000000000000000),
    .o(\u2_Display/n1540 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt56  (
    .ci(1'b0),
    .i0({\u2_Display/n1543 ,\u2_Display/n1544 ,\u2_Display/n1545 ,\u2_Display/n1546 ,\u2_Display/n1547 ,\u2_Display/n1548 ,\u2_Display/n1549 ,\u2_Display/n1550 ,\u2_Display/n1551 ,\u2_Display/n1552 ,\u2_Display/n1553 ,\u2_Display/n1554 ,\u2_Display/n1555 ,\u2_Display/n1556 ,\u2_Display/n1557 ,\u2_Display/n1558 ,\u2_Display/n1559 ,\u2_Display/n1560 ,\u2_Display/n1561 ,\u2_Display/n1562 ,\u2_Display/n1563 ,\u2_Display/n1564 ,\u2_Display/n1565 ,\u2_Display/n1566 ,\u2_Display/n1567 ,\u2_Display/n1568 ,\u2_Display/n1569 ,\u2_Display/n1570 ,\u2_Display/n1571 ,\u2_Display/n1572 ,\u2_Display/n1573 ,\u2_Display/n1574 }),
    .i1(32'b01110000100000000000000000000000),
    .o(\u2_Display/n1575 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt57  (
    .ci(1'b0),
    .i0({\u2_Display/n1578 ,\u2_Display/n1579 ,\u2_Display/n1580 ,\u2_Display/n1581 ,\u2_Display/n1582 ,\u2_Display/n1583 ,\u2_Display/n1584 ,\u2_Display/n1585 ,\u2_Display/n1586 ,\u2_Display/n1587 ,\u2_Display/n1588 ,\u2_Display/n1589 ,\u2_Display/n1590 ,\u2_Display/n1591 ,\u2_Display/n1592 ,\u2_Display/n1593 ,\u2_Display/n1594 ,\u2_Display/n1595 ,\u2_Display/n1596 ,\u2_Display/n1597 ,\u2_Display/n1598 ,\u2_Display/n1599 ,\u2_Display/n1600 ,\u2_Display/n1601 ,\u2_Display/n1602 ,\u2_Display/n1603 ,\u2_Display/n1604 ,\u2_Display/n1605 ,\u2_Display/n1606 ,\u2_Display/n1607 ,\u2_Display/n1608 ,\u2_Display/n1609 }),
    .i1(32'b00111000010000000000000000000000),
    .o(\u2_Display/n1610 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt58  (
    .ci(1'b0),
    .i0({\u2_Display/n1613 ,\u2_Display/n1614 ,\u2_Display/n1615 ,\u2_Display/n1616 ,\u2_Display/n1617 ,\u2_Display/n1618 ,\u2_Display/n1619 ,\u2_Display/n1620 ,\u2_Display/n1621 ,\u2_Display/n1622 ,\u2_Display/n1623 ,\u2_Display/n1624 ,\u2_Display/n1625 ,\u2_Display/n1626 ,\u2_Display/n1627 ,\u2_Display/n1628 ,\u2_Display/n1629 ,\u2_Display/n1630 ,\u2_Display/n1631 ,\u2_Display/n1632 ,\u2_Display/n1633 ,\u2_Display/n1634 ,\u2_Display/n1635 ,\u2_Display/n1636 ,\u2_Display/n1637 ,\u2_Display/n1638 ,\u2_Display/n1639 ,\u2_Display/n1640 ,\u2_Display/n1641 ,\u2_Display/n1642 ,\u2_Display/n1643 ,\u2_Display/n1644 }),
    .i1(32'b00011100001000000000000000000000),
    .o(\u2_Display/n1645 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt59  (
    .ci(1'b0),
    .i0({\u2_Display/n1648 ,\u2_Display/n1649 ,\u2_Display/n1650 ,\u2_Display/n1651 ,\u2_Display/n1652 ,\u2_Display/n1653 ,\u2_Display/n1654 ,\u2_Display/n1655 ,\u2_Display/n1656 ,\u2_Display/n1657 ,\u2_Display/n1658 ,\u2_Display/n1659 ,\u2_Display/n1660 ,\u2_Display/n1661 ,\u2_Display/n1662 ,\u2_Display/n1663 ,\u2_Display/n1664 ,\u2_Display/n1665 ,\u2_Display/n1666 ,\u2_Display/n1667 ,\u2_Display/n1668 ,\u2_Display/n1669 ,\u2_Display/n1670 ,\u2_Display/n1671 ,\u2_Display/n1672 ,\u2_Display/n1673 ,\u2_Display/n1674 ,\u2_Display/n1675 ,\u2_Display/n1676 ,\u2_Display/n1677 ,\u2_Display/n1678 ,\u2_Display/n1679 }),
    .i1(32'b00001110000100000000000000000000),
    .o(\u2_Display/n1680 ));  // source/rtl/Display.v(213)
  lt_u13_u13 \u2_Display/lt5_2  (
    .ci(1'b0),
    .i0({\u2_Display/n96 [31],\u2_Display/n96 [31],\u2_Display/n96 [10:0]}),
    .i1({1'b0,lcd_xpos}),
    .o(\u2_Display/n97 ));  // source/rtl/Display.v(181)
  lt_u32_u32 \u2_Display/lt60  (
    .ci(1'b0),
    .i0({\u2_Display/n1683 ,\u2_Display/n1684 ,\u2_Display/n1685 ,\u2_Display/n1686 ,\u2_Display/n1687 ,\u2_Display/n1688 ,\u2_Display/n1689 ,\u2_Display/n1690 ,\u2_Display/n1691 ,\u2_Display/n1692 ,\u2_Display/n1693 ,\u2_Display/n1694 ,\u2_Display/n1695 ,\u2_Display/n1696 ,\u2_Display/n1697 ,\u2_Display/n1698 ,\u2_Display/n1699 ,\u2_Display/n1700 ,\u2_Display/n1701 ,\u2_Display/n1702 ,\u2_Display/n1703 ,\u2_Display/n1704 ,\u2_Display/n1705 ,\u2_Display/n1706 ,\u2_Display/n1707 ,\u2_Display/n1708 ,\u2_Display/n1709 ,\u2_Display/n1710 ,\u2_Display/n1711 ,\u2_Display/n1712 ,\u2_Display/n1713 ,\u2_Display/n1714 }),
    .i1(32'b00000111000010000000000000000000),
    .o(\u2_Display/n1715 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt61  (
    .ci(1'b0),
    .i0({\u2_Display/n1718 ,\u2_Display/n1719 ,\u2_Display/n1720 ,\u2_Display/n1721 ,\u2_Display/n1722 ,\u2_Display/n1723 ,\u2_Display/n1724 ,\u2_Display/n1725 ,\u2_Display/n1726 ,\u2_Display/n1727 ,\u2_Display/n1728 ,\u2_Display/n1729 ,\u2_Display/n1730 ,\u2_Display/n1731 ,\u2_Display/n1732 ,\u2_Display/n1733 ,\u2_Display/n1734 ,\u2_Display/n1735 ,\u2_Display/n1736 ,\u2_Display/n1737 ,\u2_Display/n1738 ,\u2_Display/n1739 ,\u2_Display/n1740 ,\u2_Display/n1741 ,\u2_Display/n1742 ,\u2_Display/n1743 ,\u2_Display/n1744 ,\u2_Display/n1745 ,\u2_Display/n1746 ,\u2_Display/n1747 ,\u2_Display/n1748 ,\u2_Display/n1749 }),
    .i1(32'b00000011100001000000000000000000),
    .o(\u2_Display/n1750 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt62  (
    .ci(1'b0),
    .i0({\u2_Display/n1753 ,\u2_Display/n1754 ,\u2_Display/n1755 ,\u2_Display/n1756 ,\u2_Display/n1757 ,\u2_Display/n1758 ,\u2_Display/n1759 ,\u2_Display/n1760 ,\u2_Display/n1761 ,\u2_Display/n1762 ,\u2_Display/n1763 ,\u2_Display/n1764 ,\u2_Display/n1765 ,\u2_Display/n1766 ,\u2_Display/n1767 ,\u2_Display/n1768 ,\u2_Display/n1769 ,\u2_Display/n1770 ,\u2_Display/n1771 ,\u2_Display/n1772 ,\u2_Display/n1773 ,\u2_Display/n1774 ,\u2_Display/n1775 ,\u2_Display/n1776 ,\u2_Display/n1777 ,\u2_Display/n1778 ,\u2_Display/n1779 ,\u2_Display/n1780 ,\u2_Display/n1781 ,\u2_Display/n1782 ,\u2_Display/n1783 ,\u2_Display/n1784 }),
    .i1(32'b00000001110000100000000000000000),
    .o(\u2_Display/n1785 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt63  (
    .ci(1'b0),
    .i0({\u2_Display/n1788 ,\u2_Display/n1789 ,\u2_Display/n1790 ,\u2_Display/n1791 ,\u2_Display/n1792 ,\u2_Display/n1793 ,\u2_Display/n1794 ,\u2_Display/n1795 ,\u2_Display/n1796 ,\u2_Display/n1797 ,\u2_Display/n1798 ,\u2_Display/n1799 ,\u2_Display/n1800 ,\u2_Display/n1801 ,\u2_Display/n1802 ,\u2_Display/n1803 ,\u2_Display/n1804 ,\u2_Display/n1805 ,\u2_Display/n1806 ,\u2_Display/n1807 ,\u2_Display/n1808 ,\u2_Display/n1809 ,\u2_Display/n1810 ,\u2_Display/n1811 ,\u2_Display/n1812 ,\u2_Display/n1813 ,\u2_Display/n1814 ,\u2_Display/n1815 ,\u2_Display/n1816 ,\u2_Display/n1817 ,\u2_Display/n1818 ,\u2_Display/n1819 }),
    .i1(32'b00000000111000010000000000000000),
    .o(\u2_Display/n1820 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt64  (
    .ci(1'b0),
    .i0({\u2_Display/n1823 ,\u2_Display/n1824 ,\u2_Display/n1825 ,\u2_Display/n1826 ,\u2_Display/n1827 ,\u2_Display/n1828 ,\u2_Display/n1829 ,\u2_Display/n1830 ,\u2_Display/n1831 ,\u2_Display/n1832 ,\u2_Display/n1833 ,\u2_Display/n1834 ,\u2_Display/n1835 ,\u2_Display/n1836 ,\u2_Display/n1837 ,\u2_Display/n1838 ,\u2_Display/n1839 ,\u2_Display/n1840 ,\u2_Display/n1841 ,\u2_Display/n1842 ,\u2_Display/n1843 ,\u2_Display/n1844 ,\u2_Display/n1845 ,\u2_Display/n1846 ,\u2_Display/n1847 ,\u2_Display/n1848 ,\u2_Display/n1849 ,\u2_Display/n1850 ,\u2_Display/n1851 ,\u2_Display/n1852 ,\u2_Display/n1853 ,\u2_Display/n1854 }),
    .i1(32'b00000000011100001000000000000000),
    .o(\u2_Display/n1855 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt65  (
    .ci(1'b0),
    .i0({\u2_Display/n1858 ,\u2_Display/n1859 ,\u2_Display/n1860 ,\u2_Display/n1861 ,\u2_Display/n1862 ,\u2_Display/n1863 ,\u2_Display/n1864 ,\u2_Display/n1865 ,\u2_Display/n1866 ,\u2_Display/n1867 ,\u2_Display/n1868 ,\u2_Display/n1869 ,\u2_Display/n1870 ,\u2_Display/n1871 ,\u2_Display/n1872 ,\u2_Display/n1873 ,\u2_Display/n1874 ,\u2_Display/n1875 ,\u2_Display/n1876 ,\u2_Display/n1877 ,\u2_Display/n1878 ,\u2_Display/n1879 ,\u2_Display/n1880 ,\u2_Display/n1881 ,\u2_Display/n1882 ,\u2_Display/n1883 ,\u2_Display/n1884 ,\u2_Display/n1885 ,\u2_Display/n1886 ,\u2_Display/n1887 ,\u2_Display/n1888 ,\u2_Display/n1889 }),
    .i1(32'b00000000001110000100000000000000),
    .o(\u2_Display/n1890 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt66  (
    .ci(1'b0),
    .i0({\u2_Display/n1893 ,\u2_Display/n1894 ,\u2_Display/n1895 ,\u2_Display/n1896 ,\u2_Display/n1897 ,\u2_Display/n1898 ,\u2_Display/n1899 ,\u2_Display/n1900 ,\u2_Display/n1901 ,\u2_Display/n1902 ,\u2_Display/n1903 ,\u2_Display/n1904 ,\u2_Display/n1905 ,\u2_Display/n1906 ,\u2_Display/n1907 ,\u2_Display/n1908 ,\u2_Display/n1909 ,\u2_Display/n1910 ,\u2_Display/n1911 ,\u2_Display/n1912 ,\u2_Display/n1913 ,\u2_Display/n1914 ,\u2_Display/n1915 ,\u2_Display/n1916 ,\u2_Display/n1917 ,\u2_Display/n1918 ,\u2_Display/n1919 ,\u2_Display/n1920 ,\u2_Display/n1921 ,\u2_Display/n1922 ,\u2_Display/n1923 ,\u2_Display/n1924 }),
    .i1(32'b00000000000111000010000000000000),
    .o(\u2_Display/n1925 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt67  (
    .ci(1'b0),
    .i0({\u2_Display/n1928 ,\u2_Display/n1929 ,\u2_Display/n1930 ,\u2_Display/n1931 ,\u2_Display/n1932 ,\u2_Display/n1933 ,\u2_Display/n1934 ,\u2_Display/n1935 ,\u2_Display/n1936 ,\u2_Display/n1937 ,\u2_Display/n1938 ,\u2_Display/n1939 ,\u2_Display/n1940 ,\u2_Display/n1941 ,\u2_Display/n1942 ,\u2_Display/n1943 ,\u2_Display/n1944 ,\u2_Display/n1945 ,\u2_Display/n1946 ,\u2_Display/n1947 ,\u2_Display/n1948 ,\u2_Display/n1949 ,\u2_Display/n1950 ,\u2_Display/n1951 ,\u2_Display/n1952 ,\u2_Display/n1953 ,\u2_Display/n1954 ,\u2_Display/n1955 ,\u2_Display/n1956 ,\u2_Display/n1957 ,\u2_Display/n1958 ,\u2_Display/n1959 }),
    .i1(32'b00000000000011100001000000000000),
    .o(\u2_Display/n1960 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt68  (
    .ci(1'b0),
    .i0({\u2_Display/n1963 ,\u2_Display/n1964 ,\u2_Display/n1965 ,\u2_Display/n1966 ,\u2_Display/n1967 ,\u2_Display/n1968 ,\u2_Display/n1969 ,\u2_Display/n1970 ,\u2_Display/n1971 ,\u2_Display/n1972 ,\u2_Display/n1973 ,\u2_Display/n1974 ,\u2_Display/n1975 ,\u2_Display/n1976 ,\u2_Display/n1977 ,\u2_Display/n1978 ,\u2_Display/n1979 ,\u2_Display/n1980 ,\u2_Display/n1981 ,\u2_Display/n1982 ,\u2_Display/n1983 ,\u2_Display/n1984 ,\u2_Display/n1985 ,\u2_Display/n1986 ,\u2_Display/n1987 ,\u2_Display/n1988 ,\u2_Display/n1989 ,\u2_Display/n1990 ,\u2_Display/n1991 ,\u2_Display/n1992 ,\u2_Display/n1993 ,\u2_Display/n1994 }),
    .i1(32'b00000000000001110000100000000000),
    .o(\u2_Display/n1995 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt69  (
    .ci(1'b0),
    .i0({\u2_Display/n1998 ,\u2_Display/n1999 ,\u2_Display/n2000 ,\u2_Display/n2001 ,\u2_Display/n2002 ,\u2_Display/n2003 ,\u2_Display/n2004 ,\u2_Display/n2005 ,\u2_Display/n2006 ,\u2_Display/n2007 ,\u2_Display/n2008 ,\u2_Display/n2009 ,\u2_Display/n2010 ,\u2_Display/n2011 ,\u2_Display/n2012 ,\u2_Display/n2013 ,\u2_Display/n2014 ,\u2_Display/n2015 ,\u2_Display/n2016 ,\u2_Display/n2017 ,\u2_Display/n2018 ,\u2_Display/n2019 ,\u2_Display/n2020 ,\u2_Display/n2021 ,\u2_Display/n2022 ,\u2_Display/n2023 ,\u2_Display/n2024 ,\u2_Display/n2025 ,\u2_Display/n2026 ,\u2_Display/n2027 ,\u2_Display/n2028 ,\u2_Display/n2029 }),
    .i1(32'b00000000000000111000010000000000),
    .o(\u2_Display/n2030 ));  // source/rtl/Display.v(213)
  lt_u12_u12 \u2_Display/lt6_2  (
    .ci(1'b0),
    .i0(lcd_ypos),
    .i1({1'b0,\u2_Display/add5_2_co ,\u2_Display/n99 [0],\u2_Display/j [8:0]}),
    .o(\u2_Display/n100 ));  // source/rtl/Display.v(181)
  lt_u32_u32 \u2_Display/lt70  (
    .ci(1'b0),
    .i0({\u2_Display/n2033 ,\u2_Display/n2034 ,\u2_Display/n2035 ,\u2_Display/n2036 ,\u2_Display/n2037 ,\u2_Display/n2038 ,\u2_Display/n2039 ,\u2_Display/n2040 ,\u2_Display/n2041 ,\u2_Display/n2042 ,\u2_Display/n2043 ,\u2_Display/n2044 ,\u2_Display/n2045 ,\u2_Display/n2046 ,\u2_Display/n2047 ,\u2_Display/n2048 ,\u2_Display/n2049 ,\u2_Display/n2050 ,\u2_Display/n2051 ,\u2_Display/n2052 ,\u2_Display/n2053 ,\u2_Display/n2054 ,\u2_Display/n2055 ,\u2_Display/n2056 ,\u2_Display/n2057 ,\u2_Display/n2058 ,\u2_Display/n2059 ,\u2_Display/n2060 ,\u2_Display/n2061 ,\u2_Display/n2062 ,\u2_Display/n2063 ,\u2_Display/n2064 }),
    .i1(32'b00000000000000011100001000000000),
    .o(\u2_Display/n2065 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt71  (
    .ci(1'b0),
    .i0({\u2_Display/n2068 ,\u2_Display/n2069 ,\u2_Display/n2070 ,\u2_Display/n2071 ,\u2_Display/n2072 ,\u2_Display/n2073 ,\u2_Display/n2074 ,\u2_Display/n2075 ,\u2_Display/n2076 ,\u2_Display/n2077 ,\u2_Display/n2078 ,\u2_Display/n2079 ,\u2_Display/n2080 ,\u2_Display/n2081 ,\u2_Display/n2082 ,\u2_Display/n2083 ,\u2_Display/n2084 ,\u2_Display/n2085 ,\u2_Display/n2086 ,\u2_Display/n2087 ,\u2_Display/n2088 ,\u2_Display/n2089 ,\u2_Display/n2090 ,\u2_Display/n2091 ,\u2_Display/n2092 ,\u2_Display/n2093 ,\u2_Display/n2094 ,\u2_Display/n2095 ,\u2_Display/n2096 ,\u2_Display/n2097 ,\u2_Display/n2098 ,\u2_Display/n2099 }),
    .i1(32'b00000000000000001110000100000000),
    .o(\u2_Display/n2100 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt72  (
    .ci(1'b0),
    .i0({\u2_Display/n2103 ,\u2_Display/n2104 ,\u2_Display/n2105 ,\u2_Display/n2106 ,\u2_Display/n2107 ,\u2_Display/n2108 ,\u2_Display/n2109 ,\u2_Display/n2110 ,\u2_Display/n2111 ,\u2_Display/n2112 ,\u2_Display/n2113 ,\u2_Display/n2114 ,\u2_Display/n2115 ,\u2_Display/n2116 ,\u2_Display/n2117 ,\u2_Display/n2118 ,\u2_Display/n2119 ,\u2_Display/n2120 ,\u2_Display/n2121 ,\u2_Display/n2122 ,\u2_Display/n2123 ,\u2_Display/n2124 ,\u2_Display/n2125 ,\u2_Display/n2126 ,\u2_Display/n2127 ,\u2_Display/n2128 ,\u2_Display/n2129 ,\u2_Display/n2130 ,\u2_Display/n2131 ,\u2_Display/n2132 ,\u2_Display/n2133 ,\u2_Display/n2134 }),
    .i1(32'b00000000000000000111000010000000),
    .o(\u2_Display/n2135 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt73  (
    .ci(1'b0),
    .i0({\u2_Display/n2138 ,\u2_Display/n2139 ,\u2_Display/n2140 ,\u2_Display/n2141 ,\u2_Display/n2142 ,\u2_Display/n2143 ,\u2_Display/n2144 ,\u2_Display/n2145 ,\u2_Display/n2146 ,\u2_Display/n2147 ,\u2_Display/n2148 ,\u2_Display/n2149 ,\u2_Display/n2150 ,\u2_Display/n2151 ,\u2_Display/n2152 ,\u2_Display/n2153 ,\u2_Display/n2154 ,\u2_Display/n2155 ,\u2_Display/n2156 ,\u2_Display/n2157 ,\u2_Display/n2158 ,\u2_Display/n2159 ,\u2_Display/n2160 ,\u2_Display/n2161 ,\u2_Display/n2162 ,\u2_Display/n2163 ,\u2_Display/n2164 ,\u2_Display/n2165 ,\u2_Display/n2166 ,\u2_Display/n2167 ,\u2_Display/n2168 ,\u2_Display/n2169 }),
    .i1(32'b00000000000000000011100001000000),
    .o(\u2_Display/n2170 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt74  (
    .ci(1'b0),
    .i0({\u2_Display/n2173 ,\u2_Display/n2174 ,\u2_Display/n2175 ,\u2_Display/n2176 ,\u2_Display/n2177 ,\u2_Display/n2178 ,\u2_Display/n2179 ,\u2_Display/n2180 ,\u2_Display/n2181 ,\u2_Display/n2182 ,\u2_Display/n2183 ,\u2_Display/n2184 ,\u2_Display/n2185 ,\u2_Display/n2186 ,\u2_Display/n2187 ,\u2_Display/n2188 ,\u2_Display/n2189 ,\u2_Display/n2190 ,\u2_Display/n2191 ,\u2_Display/n2192 ,\u2_Display/n2193 ,\u2_Display/n2194 ,\u2_Display/n2195 ,\u2_Display/n2196 ,\u2_Display/n2197 ,\u2_Display/n2198 ,\u2_Display/n2199 ,\u2_Display/n2200 ,\u2_Display/n2201 ,\u2_Display/n2202 ,\u2_Display/n2203 ,\u2_Display/n2204 }),
    .i1(32'b00000000000000000001110000100000),
    .o(\u2_Display/n2205 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt75  (
    .ci(1'b0),
    .i0({\u2_Display/n2208 ,\u2_Display/n2209 ,\u2_Display/n2210 ,\u2_Display/n2211 ,\u2_Display/n2212 ,\u2_Display/n2213 ,\u2_Display/n2214 ,\u2_Display/n2215 ,\u2_Display/n2216 ,\u2_Display/n2217 ,\u2_Display/n2218 ,\u2_Display/n2219 ,\u2_Display/n2220 ,\u2_Display/n2221 ,\u2_Display/n2222 ,\u2_Display/n2223 ,\u2_Display/n2224 ,\u2_Display/n2225 ,\u2_Display/n2226 ,\u2_Display/n2227 ,\u2_Display/n2228 ,\u2_Display/n2229 ,\u2_Display/n2230 ,\u2_Display/n2231 ,\u2_Display/n2232 ,\u2_Display/n2233 ,\u2_Display/n2234 ,\u2_Display/n2235 ,\u2_Display/n2236 ,\u2_Display/n2237 ,\u2_Display/n2238 ,\u2_Display/n2239 }),
    .i1(32'b00000000000000000000111000010000),
    .o(\u2_Display/n2240 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt76  (
    .ci(1'b0),
    .i0({\u2_Display/n2243 ,\u2_Display/n2244 ,\u2_Display/n2245 ,\u2_Display/n2246 ,\u2_Display/n2247 ,\u2_Display/n2248 ,\u2_Display/n2249 ,\u2_Display/n2250 ,\u2_Display/n2251 ,\u2_Display/n2252 ,\u2_Display/n2253 ,\u2_Display/n2254 ,\u2_Display/n2255 ,\u2_Display/n2256 ,\u2_Display/n2257 ,\u2_Display/n2258 ,\u2_Display/n2259 ,\u2_Display/n2260 ,\u2_Display/n2261 ,\u2_Display/n2262 ,\u2_Display/n2263 ,\u2_Display/n2264 ,\u2_Display/n2265 ,\u2_Display/n2266 ,\u2_Display/n2267 ,\u2_Display/n2268 ,\u2_Display/n2269 ,\u2_Display/n2270 ,\u2_Display/n2271 ,\u2_Display/n2272 ,\u2_Display/n2273 ,\u2_Display/n2274 }),
    .i1(32'b00000000000000000000011100001000),
    .o(\u2_Display/n2275 ));  // source/rtl/Display.v(213)
  lt_u32_u32 \u2_Display/lt77  (
    .ci(1'b0),
    .i0({\u2_Display/n2278 ,\u2_Display/n2279 ,\u2_Display/n2280 ,\u2_Display/n2281 ,\u2_Display/n2282 ,\u2_Display/n2283 ,\u2_Display/n2284 ,\u2_Display/n2285 ,\u2_Display/n2286 ,\u2_Display/n2287 ,\u2_Display/n2288 ,\u2_Display/n2289 ,\u2_Display/n2290 ,\u2_Display/n2291 ,\u2_Display/n2292 ,\u2_Display/n2293 ,\u2_Display/n2294 ,\u2_Display/n2295 ,\u2_Display/n2296 ,\u2_Display/n2297 ,\u2_Display/n2298 ,\u2_Display/n2299 ,\u2_Display/n2300 ,\u2_Display/n2301 ,\u2_Display/n2302 ,\u2_Display/n2303 ,\u2_Display/n2304 ,\u2_Display/n2305 ,\u2_Display/n2306 ,\u2_Display/n2307 ,\u2_Display/n2308 ,\u2_Display/n2309 }),
    .i1(32'b00000000000000000000001110000100),
    .o(\u2_Display/n2310 ));  // source/rtl/Display.v(213)
  lt_u13_u13 \u2_Display/lt7_2  (
    .ci(1'b0),
    .i0({\u2_Display/n102 [31],\u2_Display/n102 [31],\u2_Display/n102 [31],\u2_Display/n102 [9:0]}),
    .i1({1'b0,lcd_ypos}),
    .o(\u2_Display/n103 ));  // source/rtl/Display.v(181)
  lt_u32_u32 \u2_Display/lt88  (
    .ci(1'b0),
    .i0(\u2_Display/counta ),
    .i1(32'b10010110000000000000000000000000),
    .o(\u2_Display/n2663 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt89  (
    .ci(1'b0),
    .i0({\u2_Display/n2666 ,\u2_Display/n2667 ,\u2_Display/n2668 ,\u2_Display/n2669 ,\u2_Display/n2670 ,\u2_Display/n2671 ,\u2_Display/n2672 ,\u2_Display/n2673 ,\u2_Display/n2674 ,\u2_Display/n2675 ,\u2_Display/n2676 ,\u2_Display/n2677 ,\u2_Display/n2678 ,\u2_Display/n2679 ,\u2_Display/n2680 ,\u2_Display/n2681 ,\u2_Display/n2682 ,\u2_Display/n2683 ,\u2_Display/n2684 ,\u2_Display/n2685 ,\u2_Display/n2686 ,\u2_Display/n2687 ,\u2_Display/n2688 ,\u2_Display/n2689 ,\u2_Display/n2690 ,\u2_Display/n2691 ,\u2_Display/n2692 ,\u2_Display/n2693 ,\u2_Display/n2694 ,\u2_Display/n2695 ,\u2_Display/n2696 ,\u2_Display/n2697 }),
    .i1(32'b01001011000000000000000000000000),
    .o(\u2_Display/n2698 ));  // source/rtl/Display.v(196)
  lt_u12_u12 \u2_Display/lt8_2  (
    .ci(1'b0),
    .i0(lcd_xpos),
    .i1({1'b0,\u2_Display/add6_2_co ,\u2_Display/n135 [2:0],\u2_Display/j [6:0]}),
    .o(\u2_Display/n136 ));  // source/rtl/Display.v(197)
  lt_u32_u32 \u2_Display/lt90  (
    .ci(1'b0),
    .i0({\u2_Display/n2701 ,\u2_Display/n2702 ,\u2_Display/n2703 ,\u2_Display/n2704 ,\u2_Display/n2705 ,\u2_Display/n2706 ,\u2_Display/n2707 ,\u2_Display/n2708 ,\u2_Display/n2709 ,\u2_Display/n2710 ,\u2_Display/n2711 ,\u2_Display/n2712 ,\u2_Display/n2713 ,\u2_Display/n2714 ,\u2_Display/n2715 ,\u2_Display/n2716 ,\u2_Display/n2717 ,\u2_Display/n2718 ,\u2_Display/n2719 ,\u2_Display/n2720 ,\u2_Display/n2721 ,\u2_Display/n2722 ,\u2_Display/n2723 ,\u2_Display/n2724 ,\u2_Display/n2725 ,\u2_Display/n2726 ,\u2_Display/n2727 ,\u2_Display/n2728 ,\u2_Display/n2729 ,\u2_Display/n2730 ,\u2_Display/n2731 ,\u2_Display/n2732 }),
    .i1(32'b00100101100000000000000000000000),
    .o(\u2_Display/n2733 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt91  (
    .ci(1'b0),
    .i0({\u2_Display/n2736 ,\u2_Display/n2737 ,\u2_Display/n2738 ,\u2_Display/n2739 ,\u2_Display/n2740 ,\u2_Display/n2741 ,\u2_Display/n2742 ,\u2_Display/n2743 ,\u2_Display/n2744 ,\u2_Display/n2745 ,\u2_Display/n2746 ,\u2_Display/n2747 ,\u2_Display/n2748 ,\u2_Display/n2749 ,\u2_Display/n2750 ,\u2_Display/n2751 ,\u2_Display/n2752 ,\u2_Display/n2753 ,\u2_Display/n2754 ,\u2_Display/n2755 ,\u2_Display/n2756 ,\u2_Display/n2757 ,\u2_Display/n2758 ,\u2_Display/n2759 ,\u2_Display/n2760 ,\u2_Display/n2761 ,\u2_Display/n2762 ,\u2_Display/n2763 ,\u2_Display/n2764 ,\u2_Display/n2765 ,\u2_Display/n2766 ,\u2_Display/n2767 }),
    .i1(32'b00010010110000000000000000000000),
    .o(\u2_Display/n2768 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt92  (
    .ci(1'b0),
    .i0({\u2_Display/n2771 ,\u2_Display/n2772 ,\u2_Display/n2773 ,\u2_Display/n2774 ,\u2_Display/n2775 ,\u2_Display/n2776 ,\u2_Display/n2777 ,\u2_Display/n2778 ,\u2_Display/n2779 ,\u2_Display/n2780 ,\u2_Display/n2781 ,\u2_Display/n2782 ,\u2_Display/n2783 ,\u2_Display/n2784 ,\u2_Display/n2785 ,\u2_Display/n2786 ,\u2_Display/n2787 ,\u2_Display/n2788 ,\u2_Display/n2789 ,\u2_Display/n2790 ,\u2_Display/n2791 ,\u2_Display/n2792 ,\u2_Display/n2793 ,\u2_Display/n2794 ,\u2_Display/n2795 ,\u2_Display/n2796 ,\u2_Display/n2797 ,\u2_Display/n2798 ,\u2_Display/n2799 ,\u2_Display/n2800 ,\u2_Display/n2801 ,\u2_Display/n2802 }),
    .i1(32'b00001001011000000000000000000000),
    .o(\u2_Display/n2803 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt93  (
    .ci(1'b0),
    .i0({\u2_Display/n2806 ,\u2_Display/n2807 ,\u2_Display/n2808 ,\u2_Display/n2809 ,\u2_Display/n2810 ,\u2_Display/n2811 ,\u2_Display/n2812 ,\u2_Display/n2813 ,\u2_Display/n2814 ,\u2_Display/n2815 ,\u2_Display/n2816 ,\u2_Display/n2817 ,\u2_Display/n2818 ,\u2_Display/n2819 ,\u2_Display/n2820 ,\u2_Display/n2821 ,\u2_Display/n2822 ,\u2_Display/n2823 ,\u2_Display/n2824 ,\u2_Display/n2825 ,\u2_Display/n2826 ,\u2_Display/n2827 ,\u2_Display/n2828 ,\u2_Display/n2829 ,\u2_Display/n2830 ,\u2_Display/n2831 ,\u2_Display/n2832 ,\u2_Display/n2833 ,\u2_Display/n2834 ,\u2_Display/n2835 ,\u2_Display/n2836 ,\u2_Display/n2837 }),
    .i1(32'b00000100101100000000000000000000),
    .o(\u2_Display/n2838 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt94  (
    .ci(1'b0),
    .i0({\u2_Display/n2841 ,\u2_Display/n2842 ,\u2_Display/n2843 ,\u2_Display/n2844 ,\u2_Display/n2845 ,\u2_Display/n2846 ,\u2_Display/n2847 ,\u2_Display/n2848 ,\u2_Display/n2849 ,\u2_Display/n2850 ,\u2_Display/n2851 ,\u2_Display/n2852 ,\u2_Display/n2853 ,\u2_Display/n2854 ,\u2_Display/n2855 ,\u2_Display/n2856 ,\u2_Display/n2857 ,\u2_Display/n2858 ,\u2_Display/n2859 ,\u2_Display/n2860 ,\u2_Display/n2861 ,\u2_Display/n2862 ,\u2_Display/n2863 ,\u2_Display/n2864 ,\u2_Display/n2865 ,\u2_Display/n2866 ,\u2_Display/n2867 ,\u2_Display/n2868 ,\u2_Display/n2869 ,\u2_Display/n2870 ,\u2_Display/n2871 ,\u2_Display/n2872 }),
    .i1(32'b00000010010110000000000000000000),
    .o(\u2_Display/n2873 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt95  (
    .ci(1'b0),
    .i0({\u2_Display/n2876 ,\u2_Display/n2877 ,\u2_Display/n2878 ,\u2_Display/n2879 ,\u2_Display/n2880 ,\u2_Display/n2881 ,\u2_Display/n2882 ,\u2_Display/n2883 ,\u2_Display/n2884 ,\u2_Display/n2885 ,\u2_Display/n2886 ,\u2_Display/n2887 ,\u2_Display/n2888 ,\u2_Display/n2889 ,\u2_Display/n2890 ,\u2_Display/n2891 ,\u2_Display/n2892 ,\u2_Display/n2893 ,\u2_Display/n2894 ,\u2_Display/n2895 ,\u2_Display/n2896 ,\u2_Display/n2897 ,\u2_Display/n2898 ,\u2_Display/n2899 ,\u2_Display/n2900 ,\u2_Display/n2901 ,\u2_Display/n2902 ,\u2_Display/n2903 ,\u2_Display/n2904 ,\u2_Display/n2905 ,\u2_Display/n2906 ,\u2_Display/n2907 }),
    .i1(32'b00000001001011000000000000000000),
    .o(\u2_Display/n2908 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt96  (
    .ci(1'b0),
    .i0({\u2_Display/n2911 ,\u2_Display/n2912 ,\u2_Display/n2913 ,\u2_Display/n2914 ,\u2_Display/n2915 ,\u2_Display/n2916 ,\u2_Display/n2917 ,\u2_Display/n2918 ,\u2_Display/n2919 ,\u2_Display/n2920 ,\u2_Display/n2921 ,\u2_Display/n2922 ,\u2_Display/n2923 ,\u2_Display/n2924 ,\u2_Display/n2925 ,\u2_Display/n2926 ,\u2_Display/n2927 ,\u2_Display/n2928 ,\u2_Display/n2929 ,\u2_Display/n2930 ,\u2_Display/n2931 ,\u2_Display/n2932 ,\u2_Display/n2933 ,\u2_Display/n2934 ,\u2_Display/n2935 ,\u2_Display/n2936 ,\u2_Display/n2937 ,\u2_Display/n2938 ,\u2_Display/n2939 ,\u2_Display/n2940 ,\u2_Display/n2941 ,\u2_Display/n2942 }),
    .i1(32'b00000000100101100000000000000000),
    .o(\u2_Display/n2943 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt97  (
    .ci(1'b0),
    .i0({\u2_Display/n2946 ,\u2_Display/n2947 ,\u2_Display/n2948 ,\u2_Display/n2949 ,\u2_Display/n2950 ,\u2_Display/n2951 ,\u2_Display/n2952 ,\u2_Display/n2953 ,\u2_Display/n2954 ,\u2_Display/n2955 ,\u2_Display/n2956 ,\u2_Display/n2957 ,\u2_Display/n2958 ,\u2_Display/n2959 ,\u2_Display/n2960 ,\u2_Display/n2961 ,\u2_Display/n2962 ,\u2_Display/n2963 ,\u2_Display/n2964 ,\u2_Display/n2965 ,\u2_Display/n2966 ,\u2_Display/n2967 ,\u2_Display/n2968 ,\u2_Display/n2969 ,\u2_Display/n2970 ,\u2_Display/n2971 ,\u2_Display/n2972 ,\u2_Display/n2973 ,\u2_Display/n2974 ,\u2_Display/n2975 ,\u2_Display/n2976 ,\u2_Display/n2977 }),
    .i1(32'b00000000010010110000000000000000),
    .o(\u2_Display/n2978 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt98  (
    .ci(1'b0),
    .i0({\u2_Display/n2981 ,\u2_Display/n2982 ,\u2_Display/n2983 ,\u2_Display/n2984 ,\u2_Display/n2985 ,\u2_Display/n2986 ,\u2_Display/n2987 ,\u2_Display/n2988 ,\u2_Display/n2989 ,\u2_Display/n2990 ,\u2_Display/n2991 ,\u2_Display/n2992 ,\u2_Display/n2993 ,\u2_Display/n2994 ,\u2_Display/n2995 ,\u2_Display/n2996 ,\u2_Display/n2997 ,\u2_Display/n2998 ,\u2_Display/n2999 ,\u2_Display/n3000 ,\u2_Display/n3001 ,\u2_Display/n3002 ,\u2_Display/n3003 ,\u2_Display/n3004 ,\u2_Display/n3005 ,\u2_Display/n3006 ,\u2_Display/n3007 ,\u2_Display/n3008 ,\u2_Display/n3009 ,\u2_Display/n3010 ,\u2_Display/n3011 ,\u2_Display/n3012 }),
    .i1(32'b00000000001001011000000000000000),
    .o(\u2_Display/n3013 ));  // source/rtl/Display.v(196)
  lt_u32_u32 \u2_Display/lt99  (
    .ci(1'b0),
    .i0({\u2_Display/n3016 ,\u2_Display/n3017 ,\u2_Display/n3018 ,\u2_Display/n3019 ,\u2_Display/n3020 ,\u2_Display/n3021 ,\u2_Display/n3022 ,\u2_Display/n3023 ,\u2_Display/n3024 ,\u2_Display/n3025 ,\u2_Display/n3026 ,\u2_Display/n3027 ,\u2_Display/n3028 ,\u2_Display/n3029 ,\u2_Display/n3030 ,\u2_Display/n3031 ,\u2_Display/n3032 ,\u2_Display/n3033 ,\u2_Display/n3034 ,\u2_Display/n3035 ,\u2_Display/n3036 ,\u2_Display/n3037 ,\u2_Display/n3038 ,\u2_Display/n3039 ,\u2_Display/n3040 ,\u2_Display/n3041 ,\u2_Display/n3042 ,\u2_Display/n3043 ,\u2_Display/n3044 ,\u2_Display/n3045 ,\u2_Display/n3046 ,\u2_Display/n3047 }),
    .i1(32'b00000000000100101100000000000000),
    .o(\u2_Display/n3048 ));  // source/rtl/Display.v(196)
  lt_u13_u13 \u2_Display/lt9_2  (
    .ci(1'b0),
    .i0({\u2_Display/n137 [31],\u2_Display/n137 [31],\u2_Display/n137 [31],\u2_Display/n137 [9:0]}),
    .i1({1'b0,lcd_xpos}),
    .o(\u2_Display/n138 ));  // source/rtl/Display.v(197)
  binary_mux_s1_w1 \u2_Display/mux10_b0  (
    .i0(\u2_Display/n226 [0]),
    .i1(\u2_Display/n133 [0]),
    .sel(on_off[2]),
    .o(\u2_Display/n230 [0]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux10_b1  (
    .i0(\u2_Display/n226 [1]),
    .i1(\u2_Display/n133 [1]),
    .sel(on_off[2]),
    .o(\u2_Display/n230 [1]));  // source/rtl/Display.v(242)
  and \u2_Display/mux10_b10_sel_is_2  (\u2_Display/mux10_b10_sel_is_2_o , \on_off[2]_neg , \u2_Display/mux5_b0_sel_is_0_o );
  binary_mux_s1_w1 \u2_Display/mux10_b2  (
    .i0(\u2_Display/n226 [2]),
    .i1(\u2_Display/n133 [2]),
    .sel(on_off[2]),
    .o(\u2_Display/n230 [2]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux10_b3  (
    .i0(\u2_Display/n226 [3]),
    .i1(\u2_Display/n133 [3]),
    .sel(on_off[2]),
    .o(\u2_Display/n230 [3]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux10_b4  (
    .i0(\u2_Display/n226 [4]),
    .i1(\u2_Display/n133 [4]),
    .sel(on_off[2]),
    .o(\u2_Display/n230 [4]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux10_b5  (
    .i0(\u2_Display/n226 [5]),
    .i1(\u2_Display/n133 [5]),
    .sel(on_off[2]),
    .o(\u2_Display/n230 [5]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux10_b6  (
    .i0(\u2_Display/n226 [6]),
    .i1(\u2_Display/n133 [6]),
    .sel(on_off[2]),
    .o(\u2_Display/n230 [6]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux10_b7  (
    .i0(\u2_Display/n226 [7]),
    .i1(\u2_Display/n133 [7]),
    .sel(on_off[2]),
    .o(\u2_Display/n230 [7]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux10_b8  (
    .i0(\u2_Display/n226 [8]),
    .i1(\u2_Display/n133 [8]),
    .sel(on_off[2]),
    .o(\u2_Display/n230 [8]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux10_b9  (
    .i0(\u2_Display/n226 [9]),
    .i1(\u2_Display/n133 [9]),
    .sel(on_off[2]),
    .o(\u2_Display/n230 [9]));  // source/rtl/Display.v(242)
  AL_MUX \u2_Display/mux11_b0  (
    .i0(\u2_Display/n134 [0]),
    .i1(\u2_Display/n223 [0]),
    .sel(\u2_Display/mux11_b0_sel_is_0_o ),
    .o(\u2_Display/n231 [0]));
  and \u2_Display/mux11_b0_sel_is_0  (\u2_Display/mux11_b0_sel_is_0_o , \on_off[2]_neg , \on_off[3]_neg );
  AL_MUX \u2_Display/mux11_b1  (
    .i0(\u2_Display/n134 [1]),
    .i1(\u2_Display/n223 [1]),
    .sel(\u2_Display/mux11_b0_sel_is_0_o ),
    .o(\u2_Display/n231 [1]));
  AL_MUX \u2_Display/mux11_b2  (
    .i0(\u2_Display/n134 [2]),
    .i1(\u2_Display/n223 [2]),
    .sel(\u2_Display/mux11_b0_sel_is_0_o ),
    .o(\u2_Display/n231 [2]));
  AL_MUX \u2_Display/mux11_b3  (
    .i0(\u2_Display/n134 [3]),
    .i1(\u2_Display/n223 [3]),
    .sel(\u2_Display/mux11_b0_sel_is_0_o ),
    .o(\u2_Display/n231 [3]));
  AL_MUX \u2_Display/mux11_b4  (
    .i0(\u2_Display/n134 [4]),
    .i1(\u2_Display/n223 [4]),
    .sel(\u2_Display/mux11_b0_sel_is_0_o ),
    .o(\u2_Display/n231 [4]));
  AL_MUX \u2_Display/mux11_b5  (
    .i0(\u2_Display/n134 [5]),
    .i1(\u2_Display/n223 [5]),
    .sel(\u2_Display/mux11_b0_sel_is_0_o ),
    .o(\u2_Display/n231 [5]));
  AL_MUX \u2_Display/mux11_b6  (
    .i0(\u2_Display/n134 [6]),
    .i1(\u2_Display/n223 [6]),
    .sel(\u2_Display/mux11_b0_sel_is_0_o ),
    .o(\u2_Display/n231 [6]));
  AL_MUX \u2_Display/mux11_b7  (
    .i0(\u2_Display/n134 [7]),
    .i1(\u2_Display/n223 [7]),
    .sel(\u2_Display/mux11_b0_sel_is_0_o ),
    .o(\u2_Display/n231 [7]));
  AL_MUX \u2_Display/mux11_b8  (
    .i0(\u2_Display/n134 [8]),
    .i1(\u2_Display/n223 [8]),
    .sel(\u2_Display/mux11_b0_sel_is_0_o ),
    .o(\u2_Display/n231 [8]));
  AL_MUX \u2_Display/mux11_b9  (
    .i0(\u2_Display/n134 [9]),
    .i1(\u2_Display/n223 [9]),
    .sel(\u2_Display/mux11_b0_sel_is_0_o ),
    .o(\u2_Display/n231 [9]));
  AL_MUX \u2_Display/mux12_b0  (
    .i0(\u2_Display/n145 ),
    .i1(1'b0),
    .sel(\u2_Display/mux10_b10_sel_is_2_o ),
    .o(\u2_Display/n232 [0]));
  and \u2_Display/mux13_b0_sel_is_2  (\u2_Display/mux13_b0_sel_is_2_o , \on_off[1]_neg , \u2_Display/mux10_b10_sel_is_2_o );
  binary_mux_s1_w1 \u2_Display/mux14_b0  (
    .i0(\u2_Display/n230 [0]),
    .i1(\u2_Display/n93 [0]),
    .sel(on_off[1]),
    .o(\u2_Display/n234 [0]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux14_b1  (
    .i0(\u2_Display/n230 [1]),
    .i1(\u2_Display/n93 [1]),
    .sel(on_off[1]),
    .o(\u2_Display/n234 [1]));  // source/rtl/Display.v(242)
  AL_MUX \u2_Display/mux14_b10  (
    .i0(1'b0),
    .i1(\u2_Display/i [10]),
    .sel(\u2_Display/mux13_b0_sel_is_2_o ),
    .o(\u2_Display/n234 [10]));
  binary_mux_s1_w1 \u2_Display/mux14_b2  (
    .i0(\u2_Display/n230 [2]),
    .i1(\u2_Display/n93 [2]),
    .sel(on_off[1]),
    .o(\u2_Display/n234 [2]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux14_b3  (
    .i0(\u2_Display/n230 [3]),
    .i1(\u2_Display/n93 [3]),
    .sel(on_off[1]),
    .o(\u2_Display/n234 [3]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux14_b4  (
    .i0(\u2_Display/n230 [4]),
    .i1(\u2_Display/n93 [4]),
    .sel(on_off[1]),
    .o(\u2_Display/n234 [4]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux14_b5  (
    .i0(\u2_Display/n230 [5]),
    .i1(\u2_Display/n93 [5]),
    .sel(on_off[1]),
    .o(\u2_Display/n234 [5]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux14_b6  (
    .i0(\u2_Display/n230 [6]),
    .i1(\u2_Display/n93 [6]),
    .sel(on_off[1]),
    .o(\u2_Display/n234 [6]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux14_b7  (
    .i0(\u2_Display/n230 [7]),
    .i1(\u2_Display/n93 [7]),
    .sel(on_off[1]),
    .o(\u2_Display/n234 [7]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux14_b8  (
    .i0(\u2_Display/n230 [8]),
    .i1(\u2_Display/n93 [8]),
    .sel(on_off[1]),
    .o(\u2_Display/n234 [8]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux14_b9  (
    .i0(\u2_Display/n230 [9]),
    .i1(\u2_Display/n93 [9]),
    .sel(on_off[1]),
    .o(\u2_Display/n234 [9]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux15_b9  (
    .i0(\u2_Display/n231 [9]),
    .i1(1'b0),
    .sel(on_off[1]),
    .o(\u2_Display/n235 [9]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux16_b0  (
    .i0(\u2_Display/n232 [0]),
    .i1(\u2_Display/n104 ),
    .sel(on_off[1]),
    .o(\u2_Display/n236 [0]));  // source/rtl/Display.v(242)
  and \u2_Display/mux17_b0_sel_is_2  (\u2_Display/mux17_b0_sel_is_2_o , \on_off[0]_neg , \u2_Display/mux13_b0_sel_is_2_o );
  not \u2_Display/mux17_b0_sel_is_2_o_inv  (\u2_Display/mux17_b0_sel_is_2_o_neg , \u2_Display/mux17_b0_sel_is_2_o );
  binary_mux_s1_w1 \u2_Display/mux18_b0  (
    .i0(\u2_Display/n234 [0]),
    .i1(\u2_Display/n42 [0]),
    .sel(on_off[0]),
    .o(\u2_Display/n238 [0]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux18_b1  (
    .i0(\u2_Display/n234 [1]),
    .i1(\u2_Display/n42 [1]),
    .sel(on_off[0]),
    .o(\u2_Display/n238 [1]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux18_b10  (
    .i0(\u2_Display/n234 [10]),
    .i1(\u2_Display/n42 [10]),
    .sel(on_off[0]),
    .o(\u2_Display/n238 [10]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux18_b2  (
    .i0(\u2_Display/n234 [2]),
    .i1(\u2_Display/n42 [2]),
    .sel(on_off[0]),
    .o(\u2_Display/n238 [2]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux18_b3  (
    .i0(\u2_Display/n234 [3]),
    .i1(\u2_Display/n42 [3]),
    .sel(on_off[0]),
    .o(\u2_Display/n238 [3]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux18_b4  (
    .i0(\u2_Display/n234 [4]),
    .i1(\u2_Display/n42 [4]),
    .sel(on_off[0]),
    .o(\u2_Display/n238 [4]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux18_b5  (
    .i0(\u2_Display/n234 [5]),
    .i1(\u2_Display/n42 [5]),
    .sel(on_off[0]),
    .o(\u2_Display/n238 [5]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux18_b6  (
    .i0(\u2_Display/n234 [6]),
    .i1(\u2_Display/n42 [6]),
    .sel(on_off[0]),
    .o(\u2_Display/n238 [6]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux18_b7  (
    .i0(\u2_Display/n234 [7]),
    .i1(\u2_Display/n42 [7]),
    .sel(on_off[0]),
    .o(\u2_Display/n238 [7]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux18_b8  (
    .i0(\u2_Display/n234 [8]),
    .i1(\u2_Display/n42 [8]),
    .sel(on_off[0]),
    .o(\u2_Display/n238 [8]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux18_b9  (
    .i0(\u2_Display/n234 [9]),
    .i1(\u2_Display/n42 [9]),
    .sel(on_off[0]),
    .o(\u2_Display/n238 [9]));  // source/rtl/Display.v(242)
  AL_MUX \u2_Display/mux19_b0  (
    .i0(\u2_Display/counta [0]),
    .i1(\u2_Display/n231 [0]),
    .sel(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n239 [0]));
  and \u2_Display/mux19_b0_sel_is_0  (\u2_Display/mux19_b0_sel_is_0_o , \on_off[0]_neg , \on_off[1]_neg );
  AL_MUX \u2_Display/mux19_b1  (
    .i0(\u2_Display/counta [1]),
    .i1(\u2_Display/n231 [1]),
    .sel(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n239 [1]));
  AL_MUX \u2_Display/mux19_b2  (
    .i0(\u2_Display/counta [2]),
    .i1(\u2_Display/n231 [2]),
    .sel(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n239 [2]));
  AL_MUX \u2_Display/mux19_b3  (
    .i0(\u2_Display/counta [3]),
    .i1(\u2_Display/n231 [3]),
    .sel(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n239 [3]));
  AL_MUX \u2_Display/mux19_b4  (
    .i0(\u2_Display/counta [4]),
    .i1(\u2_Display/n231 [4]),
    .sel(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n239 [4]));
  AL_MUX \u2_Display/mux19_b5  (
    .i0(\u2_Display/counta [5]),
    .i1(\u2_Display/n231 [5]),
    .sel(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n239 [5]));
  AL_MUX \u2_Display/mux19_b6  (
    .i0(\u2_Display/counta [6]),
    .i1(\u2_Display/n231 [6]),
    .sel(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n239 [6]));
  AL_MUX \u2_Display/mux19_b7  (
    .i0(\u2_Display/counta [7]),
    .i1(\u2_Display/n231 [7]),
    .sel(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n239 [7]));
  AL_MUX \u2_Display/mux19_b8  (
    .i0(\u2_Display/counta [8]),
    .i1(\u2_Display/n231 [8]),
    .sel(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n239 [8]));
  binary_mux_s1_w1 \u2_Display/mux19_b9  (
    .i0(\u2_Display/n235 [9]),
    .i1(\u2_Display/counta [9]),
    .sel(on_off[0]),
    .o(\u2_Display/n239 [9]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux20_b0  (
    .i0(\u2_Display/n236 [0]),
    .i1(\u2_Display/n51 ),
    .sel(on_off[0]),
    .o(\u2_Display/n240 [0]));  // source/rtl/Display.v(242)
  and \u2_Display/mux21_b0_sel_is_0  (\u2_Display/mux21_b0_sel_is_0_o , rst_n, \u2_Display/mux17_b0_sel_is_2_o_neg );
  binary_mux_s1_w1 \u2_Display/mux3_b0  (
    .i0(\u2_Display/j [0]),
    .i1(\u2_Display/n196 [0]),
    .sel(on_off[4]),
    .o(\u2_Display/n223 [0]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux3_b1  (
    .i0(\u2_Display/j [1]),
    .i1(\u2_Display/n196 [1]),
    .sel(on_off[4]),
    .o(\u2_Display/n223 [1]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux3_b2  (
    .i0(\u2_Display/j [2]),
    .i1(\u2_Display/n196 [2]),
    .sel(on_off[4]),
    .o(\u2_Display/n223 [2]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux3_b3  (
    .i0(\u2_Display/j [3]),
    .i1(\u2_Display/n196 [3]),
    .sel(on_off[4]),
    .o(\u2_Display/n223 [3]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux3_b4  (
    .i0(\u2_Display/j [4]),
    .i1(\u2_Display/n196 [4]),
    .sel(on_off[4]),
    .o(\u2_Display/n223 [4]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux3_b5  (
    .i0(\u2_Display/j [5]),
    .i1(\u2_Display/n196 [5]),
    .sel(on_off[4]),
    .o(\u2_Display/n223 [5]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux3_b6  (
    .i0(\u2_Display/j [6]),
    .i1(\u2_Display/n196 [6]),
    .sel(on_off[4]),
    .o(\u2_Display/n223 [6]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux3_b7  (
    .i0(\u2_Display/j [7]),
    .i1(\u2_Display/n196 [7]),
    .sel(on_off[4]),
    .o(\u2_Display/n223 [7]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux3_b8  (
    .i0(\u2_Display/j [8]),
    .i1(\u2_Display/n196 [8]),
    .sel(on_off[4]),
    .o(\u2_Display/n223 [8]));  // source/rtl/Display.v(242)
  binary_mux_s1_w1 \u2_Display/mux3_b9  (
    .i0(\u2_Display/j [9]),
    .i1(\u2_Display/n196 [9]),
    .sel(on_off[4]),
    .o(\u2_Display/n223 [9]));  // source/rtl/Display.v(242)
  and \u2_Display/mux5_b0_sel_is_0  (\u2_Display/mux5_b0_sel_is_0_o , \on_off[3]_neg , \on_off[4]_neg );
  AL_MUX \u2_Display/mux6_b0  (
    .i0(\u2_Display/n147 [0]),
    .i1(\u2_Display/i [0]),
    .sel(\u2_Display/mux5_b0_sel_is_0_o ),
    .o(\u2_Display/n226 [0]));
  AL_MUX \u2_Display/mux6_b1  (
    .i0(\u2_Display/n147 [1]),
    .i1(\u2_Display/i [1]),
    .sel(\u2_Display/mux5_b0_sel_is_0_o ),
    .o(\u2_Display/n226 [1]));
  AL_MUX \u2_Display/mux6_b2  (
    .i0(\u2_Display/n147 [2]),
    .i1(\u2_Display/i [2]),
    .sel(\u2_Display/mux5_b0_sel_is_0_o ),
    .o(\u2_Display/n226 [2]));
  AL_MUX \u2_Display/mux6_b3  (
    .i0(\u2_Display/n147 [3]),
    .i1(\u2_Display/i [3]),
    .sel(\u2_Display/mux5_b0_sel_is_0_o ),
    .o(\u2_Display/n226 [3]));
  AL_MUX \u2_Display/mux6_b4  (
    .i0(\u2_Display/n147 [4]),
    .i1(\u2_Display/i [4]),
    .sel(\u2_Display/mux5_b0_sel_is_0_o ),
    .o(\u2_Display/n226 [4]));
  AL_MUX \u2_Display/mux6_b5  (
    .i0(\u2_Display/n147 [5]),
    .i1(\u2_Display/i [5]),
    .sel(\u2_Display/mux5_b0_sel_is_0_o ),
    .o(\u2_Display/n226 [5]));
  AL_MUX \u2_Display/mux6_b6  (
    .i0(\u2_Display/n147 [6]),
    .i1(\u2_Display/i [6]),
    .sel(\u2_Display/mux5_b0_sel_is_0_o ),
    .o(\u2_Display/n226 [6]));
  AL_MUX \u2_Display/mux6_b7  (
    .i0(\u2_Display/n147 [7]),
    .i1(\u2_Display/i [7]),
    .sel(\u2_Display/mux5_b0_sel_is_0_o ),
    .o(\u2_Display/n226 [7]));
  AL_MUX \u2_Display/mux6_b8  (
    .i0(\u2_Display/n147 [8]),
    .i1(\u2_Display/i [8]),
    .sel(\u2_Display/mux5_b0_sel_is_0_o ),
    .o(\u2_Display/n226 [8]));
  AL_MUX \u2_Display/mux6_b9  (
    .i0(\u2_Display/n147 [9]),
    .i1(\u2_Display/i [9]),
    .sel(\u2_Display/mux5_b0_sel_is_0_o ),
    .o(\u2_Display/n226 [9]));
  reg_sr_as_w1 \u2_Display/reg0_b0  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [0]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [0]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b1  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [1]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [1]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b10  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [10]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [10]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b11  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [11]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [11]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b12  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [12]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [12]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b13  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [13]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [13]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b14  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [14]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [14]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b15  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [15]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [15]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b16  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [16]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [16]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b17  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [17]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [17]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b18  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [18]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [18]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b19  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [19]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [19]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b2  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [2]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [2]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b20  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [20]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [20]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b21  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [21]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [21]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b22  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [22]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [22]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b23  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [23]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [23]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b24  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [24]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [24]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b25  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [25]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [25]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b26  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [26]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [26]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b27  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [27]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [27]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b28  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [28]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [28]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b29  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [29]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [29]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b3  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [3]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [3]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b30  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [30]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [30]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b4  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [4]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [4]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b5  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [5]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [5]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b6  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [6]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [6]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b7  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [7]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [7]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b8  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [8]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [8]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b9  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [9]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [9]));  // source/rtl/Display.v(61)
  reg_ar_as_w1 \u2_Display/reg1_b0  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n240 [0]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(lcd_data[23]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b0  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [0]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [0]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b1  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [1]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [1]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b10  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [10]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [10]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b11  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [11]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [11]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b12  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [12]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [12]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b13  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [13]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [13]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b14  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [14]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [14]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b15  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [15]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [15]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b16  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [16]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [16]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b17  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [17]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [17]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b18  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [18]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [18]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b19  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [19]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [19]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b2  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [2]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [2]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b20  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [20]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [20]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b21  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [21]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [21]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b22  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [22]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [22]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b23  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [23]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [23]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b24  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [24]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [24]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b25  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [25]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [25]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b26  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [26]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [26]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b27  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [27]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [27]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b28  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [28]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [28]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b29  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [29]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [29]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b3  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [3]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [3]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b30  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [30]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [30]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b31  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [31]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [31]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b4  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [4]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [4]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b5  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [5]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [5]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b6  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [6]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [6]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b7  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [7]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [7]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b8  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [8]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [8]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b9  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [9]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [9]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b0  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [0]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [0]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b1  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [1]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [1]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b10  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [10]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [10]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b2  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [2]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [2]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b3  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [3]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [3]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b4  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [4]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [4]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b5  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [5]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [5]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b6  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [6]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [6]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b7  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [7]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [7]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b8  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [8]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [8]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b9  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [9]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [9]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b0  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [0]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [0]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b1  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [1]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [1]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b2  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [2]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [2]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b3  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [3]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [3]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b4  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [4]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [4]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b5  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [5]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [5]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b6  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [6]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [6]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b7  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [7]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [7]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b8  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [8]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [8]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b9  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [9]),
    .en(rst_n),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [9]));  // source/rtl/Display.v(252)
  add_pu11_mu11_o12 \u2_Display/sub0_2  (
    .i0(11'b01010000000),
    .i1(\u2_Display/i [10:0]),
    .o({\u2_Display/n96 [31],\u2_Display/n96 [10:0]}));  // source/rtl/Display.v(181)
  add_pu10_mu10_o11 \u2_Display/sub1_2  (
    .i0(10'b1000000000),
    .i1(\u2_Display/j [9:0]),
    .o({\u2_Display/n102 [31],\u2_Display/n102 [9:0]}));  // source/rtl/Display.v(181)
  add_pu10_mu10_o11 \u2_Display/sub2_2  (
    .i0(10'b1010000000),
    .i1(\u2_Display/j [9:0]),
    .o({\u2_Display/n137 [31],\u2_Display/n137 [9:0]}));  // source/rtl/Display.v(197)
  add_pu11_mu11_o12 \u2_Display/sub3_2  (
    .i0(11'b01000000000),
    .i1(\u2_Display/i [10:0]),
    .o({\u2_Display/n143 [31],\u2_Display/n143 [10:0]}));  // source/rtl/Display.v(197)
  and \u2_Display/u10  (\u2_Display/n49 , \u2_Display/n46 , \u2_Display/n48 );  // source/rtl/Display.v(165)
  AL_MUX \u2_Display/u10000  (
    .i0(\u2_Display/n6319 ),
    .i1(\u2_Display/n5191 [27]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5196 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10001  (
    .i0(\u2_Display/n6320 ),
    .i1(\u2_Display/n5191 [26]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5197 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10002  (
    .i0(\u2_Display/n6321 ),
    .i1(\u2_Display/n5191 [25]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5198 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10003  (
    .i0(\u2_Display/n6322 ),
    .i1(\u2_Display/n5191 [24]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5199 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10004  (
    .i0(\u2_Display/n6323 ),
    .i1(\u2_Display/n5191 [23]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5200 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10005  (
    .i0(\u2_Display/n6324 ),
    .i1(\u2_Display/n5191 [22]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5201 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10006  (
    .i0(\u2_Display/n6325 ),
    .i1(\u2_Display/n5191 [21]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5202 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10007  (
    .i0(\u2_Display/n6326 ),
    .i1(\u2_Display/n5191 [20]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5203 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10008  (
    .i0(\u2_Display/n6327 ),
    .i1(\u2_Display/n5191 [19]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5204 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10009  (
    .i0(\u2_Display/n6328 ),
    .i1(\u2_Display/n5191 [18]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5205 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10010  (
    .i0(\u2_Display/n6329 ),
    .i1(\u2_Display/n5191 [17]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5206 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10011  (
    .i0(\u2_Display/n6330 ),
    .i1(\u2_Display/n5191 [16]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5207 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10012  (
    .i0(\u2_Display/n6331 ),
    .i1(\u2_Display/n5191 [15]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5208 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10013  (
    .i0(\u2_Display/n6332 ),
    .i1(\u2_Display/n5191 [14]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5209 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10014  (
    .i0(\u2_Display/n6333 ),
    .i1(\u2_Display/n5191 [13]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5210 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10015  (
    .i0(\u2_Display/n6334 ),
    .i1(\u2_Display/n5191 [12]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5211 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10016  (
    .i0(\u2_Display/n6335 ),
    .i1(\u2_Display/n5191 [11]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5212 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10017  (
    .i0(\u2_Display/n6336 ),
    .i1(\u2_Display/n5191 [10]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5213 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10018  (
    .i0(\u2_Display/n6337 ),
    .i1(\u2_Display/n5191 [9]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5214 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10019  (
    .i0(\u2_Display/n6338 ),
    .i1(\u2_Display/n5191 [8]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5215 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10020  (
    .i0(\u2_Display/n6339 ),
    .i1(\u2_Display/n5191 [7]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5216 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10021  (
    .i0(\u2_Display/n6340 ),
    .i1(\u2_Display/n5191 [6]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5217 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10022  (
    .i0(\u2_Display/n6341 ),
    .i1(\u2_Display/n5191 [5]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5218 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10023  (
    .i0(\u2_Display/n6342 ),
    .i1(\u2_Display/n5191 [4]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5219 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10024  (
    .i0(\u2_Display/n6343 ),
    .i1(\u2_Display/n5191 [3]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5220 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10025  (
    .i0(\u2_Display/n6344 ),
    .i1(\u2_Display/n5191 [2]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5221 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10026  (
    .i0(\u2_Display/n6345 ),
    .i1(\u2_Display/n5191 [1]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5222 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10027  (
    .i0(\u2_Display/n6346 ),
    .i1(\u2_Display/n5191 [0]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n5223 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10028  (\u2_Display/n5225 , \u2_Display/n5224 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10061  (
    .i0(\u2_Display/n6350 ),
    .i1(\u2_Display/n5226 [31]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5227 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10062  (
    .i0(\u2_Display/n6351 ),
    .i1(\u2_Display/n5226 [30]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5228 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10063  (
    .i0(\u2_Display/n6352 ),
    .i1(\u2_Display/n5226 [29]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5229 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10064  (
    .i0(\u2_Display/n6353 ),
    .i1(\u2_Display/n5226 [28]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5230 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10065  (
    .i0(\u2_Display/n5196 ),
    .i1(\u2_Display/n5226 [27]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5231 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10066  (
    .i0(\u2_Display/n5197 ),
    .i1(\u2_Display/n5226 [26]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5232 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10067  (
    .i0(\u2_Display/n5198 ),
    .i1(\u2_Display/n5226 [25]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5233 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10068  (
    .i0(\u2_Display/n5199 ),
    .i1(\u2_Display/n5226 [24]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5234 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10069  (
    .i0(\u2_Display/n5200 ),
    .i1(\u2_Display/n5226 [23]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5235 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10070  (
    .i0(\u2_Display/n5201 ),
    .i1(\u2_Display/n5226 [22]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5236 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10071  (
    .i0(\u2_Display/n5202 ),
    .i1(\u2_Display/n5226 [21]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5237 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10072  (
    .i0(\u2_Display/n5203 ),
    .i1(\u2_Display/n5226 [20]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5238 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10073  (
    .i0(\u2_Display/n5204 ),
    .i1(\u2_Display/n5226 [19]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5239 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10074  (
    .i0(\u2_Display/n5205 ),
    .i1(\u2_Display/n5226 [18]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5240 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10075  (
    .i0(\u2_Display/n5206 ),
    .i1(\u2_Display/n5226 [17]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5241 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10076  (
    .i0(\u2_Display/n5207 ),
    .i1(\u2_Display/n5226 [16]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5242 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10077  (
    .i0(\u2_Display/n5208 ),
    .i1(\u2_Display/n5226 [15]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5243 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10078  (
    .i0(\u2_Display/n5209 ),
    .i1(\u2_Display/n5226 [14]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5244 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10079  (
    .i0(\u2_Display/n5210 ),
    .i1(\u2_Display/n5226 [13]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5245 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10080  (
    .i0(\u2_Display/n5211 ),
    .i1(\u2_Display/n5226 [12]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5246 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10081  (
    .i0(\u2_Display/n5212 ),
    .i1(\u2_Display/n5226 [11]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5247 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10082  (
    .i0(\u2_Display/n5213 ),
    .i1(\u2_Display/n5226 [10]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5248 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10083  (
    .i0(\u2_Display/n5214 ),
    .i1(\u2_Display/n5226 [9]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5249 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10084  (
    .i0(\u2_Display/n5215 ),
    .i1(\u2_Display/n5226 [8]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5250 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10085  (
    .i0(\u2_Display/n5216 ),
    .i1(\u2_Display/n5226 [7]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5251 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10086  (
    .i0(\u2_Display/n5217 ),
    .i1(\u2_Display/n5226 [6]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5252 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10087  (
    .i0(\u2_Display/n5218 ),
    .i1(\u2_Display/n5226 [5]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5253 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10088  (
    .i0(\u2_Display/n5219 ),
    .i1(\u2_Display/n5226 [4]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5254 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10089  (
    .i0(\u2_Display/n5220 ),
    .i1(\u2_Display/n5226 [3]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5255 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10090  (
    .i0(\u2_Display/n5221 ),
    .i1(\u2_Display/n5226 [2]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5256 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10091  (
    .i0(\u2_Display/n5222 ),
    .i1(\u2_Display/n5226 [1]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5257 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10092  (
    .i0(\u2_Display/n5223 ),
    .i1(\u2_Display/n5226 [0]),
    .sel(\u2_Display/n5225 ),
    .o(\u2_Display/n5258 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10093  (\u2_Display/n5260 , \u2_Display/n5259 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10126  (
    .i0(\u2_Display/n5227 ),
    .i1(\u2_Display/n5261 [31]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5262 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10127  (
    .i0(\u2_Display/n5228 ),
    .i1(\u2_Display/n5261 [30]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5263 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10128  (
    .i0(\u2_Display/n5229 ),
    .i1(\u2_Display/n5261 [29]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5264 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10129  (
    .i0(\u2_Display/n5230 ),
    .i1(\u2_Display/n5261 [28]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5265 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10130  (
    .i0(\u2_Display/n5231 ),
    .i1(\u2_Display/n5261 [27]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5266 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10131  (
    .i0(\u2_Display/n5232 ),
    .i1(\u2_Display/n5261 [26]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5267 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10132  (
    .i0(\u2_Display/n5233 ),
    .i1(\u2_Display/n5261 [25]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5268 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10133  (
    .i0(\u2_Display/n5234 ),
    .i1(\u2_Display/n5261 [24]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5269 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10134  (
    .i0(\u2_Display/n5235 ),
    .i1(\u2_Display/n5261 [23]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5270 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10135  (
    .i0(\u2_Display/n5236 ),
    .i1(\u2_Display/n5261 [22]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5271 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10136  (
    .i0(\u2_Display/n5237 ),
    .i1(\u2_Display/n5261 [21]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5272 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10137  (
    .i0(\u2_Display/n5238 ),
    .i1(\u2_Display/n5261 [20]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5273 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10138  (
    .i0(\u2_Display/n5239 ),
    .i1(\u2_Display/n5261 [19]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5274 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10139  (
    .i0(\u2_Display/n5240 ),
    .i1(\u2_Display/n5261 [18]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5275 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10140  (
    .i0(\u2_Display/n5241 ),
    .i1(\u2_Display/n5261 [17]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5276 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10141  (
    .i0(\u2_Display/n5242 ),
    .i1(\u2_Display/n5261 [16]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5277 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10142  (
    .i0(\u2_Display/n5243 ),
    .i1(\u2_Display/n5261 [15]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5278 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10143  (
    .i0(\u2_Display/n5244 ),
    .i1(\u2_Display/n5261 [14]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5279 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10144  (
    .i0(\u2_Display/n5245 ),
    .i1(\u2_Display/n5261 [13]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5280 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10145  (
    .i0(\u2_Display/n5246 ),
    .i1(\u2_Display/n5261 [12]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5281 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10146  (
    .i0(\u2_Display/n5247 ),
    .i1(\u2_Display/n5261 [11]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5282 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10147  (
    .i0(\u2_Display/n5248 ),
    .i1(\u2_Display/n5261 [10]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5283 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10148  (
    .i0(\u2_Display/n5249 ),
    .i1(\u2_Display/n5261 [9]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5284 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10149  (
    .i0(\u2_Display/n5250 ),
    .i1(\u2_Display/n5261 [8]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5285 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10150  (
    .i0(\u2_Display/n5251 ),
    .i1(\u2_Display/n5261 [7]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5286 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10151  (
    .i0(\u2_Display/n5252 ),
    .i1(\u2_Display/n5261 [6]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5287 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10152  (
    .i0(\u2_Display/n5253 ),
    .i1(\u2_Display/n5261 [5]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5288 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10153  (
    .i0(\u2_Display/n5254 ),
    .i1(\u2_Display/n5261 [4]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5289 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10154  (
    .i0(\u2_Display/n5255 ),
    .i1(\u2_Display/n5261 [3]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5290 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10155  (
    .i0(\u2_Display/n5256 ),
    .i1(\u2_Display/n5261 [2]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5291 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10156  (
    .i0(\u2_Display/n5257 ),
    .i1(\u2_Display/n5261 [1]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5292 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10157  (
    .i0(\u2_Display/n5258 ),
    .i1(\u2_Display/n5261 [0]),
    .sel(\u2_Display/n5260 ),
    .o(\u2_Display/n5293 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10158  (\u2_Display/n5295 , \u2_Display/n5294 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10191  (
    .i0(\u2_Display/n5262 ),
    .i1(\u2_Display/n5296 [31]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5297 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10192  (
    .i0(\u2_Display/n5263 ),
    .i1(\u2_Display/n5296 [30]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5298 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10193  (
    .i0(\u2_Display/n5264 ),
    .i1(\u2_Display/n5296 [29]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5299 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10194  (
    .i0(\u2_Display/n5265 ),
    .i1(\u2_Display/n5296 [28]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5300 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10195  (
    .i0(\u2_Display/n5266 ),
    .i1(\u2_Display/n5296 [27]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5301 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10196  (
    .i0(\u2_Display/n5267 ),
    .i1(\u2_Display/n5296 [26]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5302 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10197  (
    .i0(\u2_Display/n5268 ),
    .i1(\u2_Display/n5296 [25]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5303 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10198  (
    .i0(\u2_Display/n5269 ),
    .i1(\u2_Display/n5296 [24]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5304 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10199  (
    .i0(\u2_Display/n5270 ),
    .i1(\u2_Display/n5296 [23]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5305 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1020  (
    .i0(\u2_Display/n525 ),
    .i1(\u2_Display/n559 [31]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n560 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10200  (
    .i0(\u2_Display/n5271 ),
    .i1(\u2_Display/n5296 [22]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5306 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10201  (
    .i0(\u2_Display/n5272 ),
    .i1(\u2_Display/n5296 [21]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5307 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10202  (
    .i0(\u2_Display/n5273 ),
    .i1(\u2_Display/n5296 [20]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5308 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10203  (
    .i0(\u2_Display/n5274 ),
    .i1(\u2_Display/n5296 [19]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5309 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10204  (
    .i0(\u2_Display/n5275 ),
    .i1(\u2_Display/n5296 [18]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5310 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10205  (
    .i0(\u2_Display/n5276 ),
    .i1(\u2_Display/n5296 [17]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5311 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10206  (
    .i0(\u2_Display/n5277 ),
    .i1(\u2_Display/n5296 [16]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5312 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10207  (
    .i0(\u2_Display/n5278 ),
    .i1(\u2_Display/n5296 [15]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5313 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10208  (
    .i0(\u2_Display/n5279 ),
    .i1(\u2_Display/n5296 [14]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5314 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10209  (
    .i0(\u2_Display/n5280 ),
    .i1(\u2_Display/n5296 [13]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5315 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1021  (
    .i0(\u2_Display/n526 ),
    .i1(\u2_Display/n559 [30]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n561 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10210  (
    .i0(\u2_Display/n5281 ),
    .i1(\u2_Display/n5296 [12]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5316 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10211  (
    .i0(\u2_Display/n5282 ),
    .i1(\u2_Display/n5296 [11]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5317 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10212  (
    .i0(\u2_Display/n5283 ),
    .i1(\u2_Display/n5296 [10]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5318 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10213  (
    .i0(\u2_Display/n5284 ),
    .i1(\u2_Display/n5296 [9]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5319 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10214  (
    .i0(\u2_Display/n5285 ),
    .i1(\u2_Display/n5296 [8]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5320 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10215  (
    .i0(\u2_Display/n5286 ),
    .i1(\u2_Display/n5296 [7]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5321 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10216  (
    .i0(\u2_Display/n5287 ),
    .i1(\u2_Display/n5296 [6]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5322 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10217  (
    .i0(\u2_Display/n5288 ),
    .i1(\u2_Display/n5296 [5]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5323 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10218  (
    .i0(\u2_Display/n5289 ),
    .i1(\u2_Display/n5296 [4]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5324 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10219  (
    .i0(\u2_Display/n5290 ),
    .i1(\u2_Display/n5296 [3]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5325 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1022  (
    .i0(\u2_Display/n527 ),
    .i1(\u2_Display/n559 [29]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n562 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10220  (
    .i0(\u2_Display/n5291 ),
    .i1(\u2_Display/n5296 [2]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5326 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10221  (
    .i0(\u2_Display/n5292 ),
    .i1(\u2_Display/n5296 [1]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5327 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10222  (
    .i0(\u2_Display/n5293 ),
    .i1(\u2_Display/n5296 [0]),
    .sel(\u2_Display/n5295 ),
    .o(\u2_Display/n5328 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10223  (\u2_Display/n5330 , \u2_Display/n5329 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1023  (
    .i0(\u2_Display/n528 ),
    .i1(\u2_Display/n559 [28]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n563 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1024  (
    .i0(\u2_Display/n529 ),
    .i1(\u2_Display/n559 [27]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n564 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1025  (
    .i0(\u2_Display/n530 ),
    .i1(\u2_Display/n559 [26]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n565 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10256  (
    .i0(\u2_Display/n5297 ),
    .i1(\u2_Display/n5331 [31]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5332 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10257  (
    .i0(\u2_Display/n5298 ),
    .i1(\u2_Display/n5331 [30]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5333 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10258  (
    .i0(\u2_Display/n5299 ),
    .i1(\u2_Display/n5331 [29]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5334 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10259  (
    .i0(\u2_Display/n5300 ),
    .i1(\u2_Display/n5331 [28]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5335 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1026  (
    .i0(\u2_Display/n531 ),
    .i1(\u2_Display/n559 [25]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n566 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10260  (
    .i0(\u2_Display/n5301 ),
    .i1(\u2_Display/n5331 [27]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5336 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10261  (
    .i0(\u2_Display/n5302 ),
    .i1(\u2_Display/n5331 [26]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5337 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10262  (
    .i0(\u2_Display/n5303 ),
    .i1(\u2_Display/n5331 [25]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5338 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10263  (
    .i0(\u2_Display/n5304 ),
    .i1(\u2_Display/n5331 [24]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5339 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10264  (
    .i0(\u2_Display/n5305 ),
    .i1(\u2_Display/n5331 [23]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5340 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10265  (
    .i0(\u2_Display/n5306 ),
    .i1(\u2_Display/n5331 [22]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5341 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10266  (
    .i0(\u2_Display/n5307 ),
    .i1(\u2_Display/n5331 [21]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5342 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10267  (
    .i0(\u2_Display/n5308 ),
    .i1(\u2_Display/n5331 [20]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5343 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10268  (
    .i0(\u2_Display/n5309 ),
    .i1(\u2_Display/n5331 [19]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5344 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10269  (
    .i0(\u2_Display/n5310 ),
    .i1(\u2_Display/n5331 [18]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5345 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1027  (
    .i0(\u2_Display/n532 ),
    .i1(\u2_Display/n559 [24]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n567 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10270  (
    .i0(\u2_Display/n5311 ),
    .i1(\u2_Display/n5331 [17]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5346 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10271  (
    .i0(\u2_Display/n5312 ),
    .i1(\u2_Display/n5331 [16]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5347 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10272  (
    .i0(\u2_Display/n5313 ),
    .i1(\u2_Display/n5331 [15]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5348 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10273  (
    .i0(\u2_Display/n5314 ),
    .i1(\u2_Display/n5331 [14]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5349 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10274  (
    .i0(\u2_Display/n5315 ),
    .i1(\u2_Display/n5331 [13]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5350 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10275  (
    .i0(\u2_Display/n5316 ),
    .i1(\u2_Display/n5331 [12]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5351 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10276  (
    .i0(\u2_Display/n5317 ),
    .i1(\u2_Display/n5331 [11]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5352 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10277  (
    .i0(\u2_Display/n5318 ),
    .i1(\u2_Display/n5331 [10]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5353 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10278  (
    .i0(\u2_Display/n5319 ),
    .i1(\u2_Display/n5331 [9]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5354 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10279  (
    .i0(\u2_Display/n5320 ),
    .i1(\u2_Display/n5331 [8]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5355 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1028  (
    .i0(\u2_Display/n533 ),
    .i1(\u2_Display/n559 [23]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n568 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10280  (
    .i0(\u2_Display/n5321 ),
    .i1(\u2_Display/n5331 [7]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5356 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10281  (
    .i0(\u2_Display/n5322 ),
    .i1(\u2_Display/n5331 [6]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5357 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10282  (
    .i0(\u2_Display/n5323 ),
    .i1(\u2_Display/n5331 [5]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5358 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10283  (
    .i0(\u2_Display/n5324 ),
    .i1(\u2_Display/n5331 [4]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5359 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10284  (
    .i0(\u2_Display/n5325 ),
    .i1(\u2_Display/n5331 [3]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5360 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10285  (
    .i0(\u2_Display/n5326 ),
    .i1(\u2_Display/n5331 [2]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5361 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10286  (
    .i0(\u2_Display/n5327 ),
    .i1(\u2_Display/n5331 [1]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5362 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10287  (
    .i0(\u2_Display/n5328 ),
    .i1(\u2_Display/n5331 [0]),
    .sel(\u2_Display/n5330 ),
    .o(\u2_Display/n5363 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10288  (\u2_Display/n5365 , \u2_Display/n5364 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1029  (
    .i0(\u2_Display/n534 ),
    .i1(\u2_Display/n559 [22]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n569 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1030  (
    .i0(\u2_Display/n535 ),
    .i1(\u2_Display/n559 [21]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n570 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1031  (
    .i0(\u2_Display/n536 ),
    .i1(\u2_Display/n559 [20]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n571 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1032  (
    .i0(\u2_Display/n537 ),
    .i1(\u2_Display/n559 [19]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n572 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10321  (
    .i0(\u2_Display/n5332 ),
    .i1(\u2_Display/n5366 [31]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5367 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10322  (
    .i0(\u2_Display/n5333 ),
    .i1(\u2_Display/n5366 [30]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5368 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10323  (
    .i0(\u2_Display/n5334 ),
    .i1(\u2_Display/n5366 [29]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5369 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10324  (
    .i0(\u2_Display/n5335 ),
    .i1(\u2_Display/n5366 [28]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5370 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10325  (
    .i0(\u2_Display/n5336 ),
    .i1(\u2_Display/n5366 [27]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5371 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10326  (
    .i0(\u2_Display/n5337 ),
    .i1(\u2_Display/n5366 [26]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5372 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10327  (
    .i0(\u2_Display/n5338 ),
    .i1(\u2_Display/n5366 [25]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5373 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10328  (
    .i0(\u2_Display/n5339 ),
    .i1(\u2_Display/n5366 [24]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5374 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10329  (
    .i0(\u2_Display/n5340 ),
    .i1(\u2_Display/n5366 [23]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5375 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1033  (
    .i0(\u2_Display/n538 ),
    .i1(\u2_Display/n559 [18]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n573 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10330  (
    .i0(\u2_Display/n5341 ),
    .i1(\u2_Display/n5366 [22]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5376 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10331  (
    .i0(\u2_Display/n5342 ),
    .i1(\u2_Display/n5366 [21]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5377 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10332  (
    .i0(\u2_Display/n5343 ),
    .i1(\u2_Display/n5366 [20]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5378 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10333  (
    .i0(\u2_Display/n5344 ),
    .i1(\u2_Display/n5366 [19]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5379 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10334  (
    .i0(\u2_Display/n5345 ),
    .i1(\u2_Display/n5366 [18]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5380 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10335  (
    .i0(\u2_Display/n5346 ),
    .i1(\u2_Display/n5366 [17]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5381 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10336  (
    .i0(\u2_Display/n5347 ),
    .i1(\u2_Display/n5366 [16]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5382 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10337  (
    .i0(\u2_Display/n5348 ),
    .i1(\u2_Display/n5366 [15]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5383 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10338  (
    .i0(\u2_Display/n5349 ),
    .i1(\u2_Display/n5366 [14]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5384 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10339  (
    .i0(\u2_Display/n5350 ),
    .i1(\u2_Display/n5366 [13]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5385 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1034  (
    .i0(\u2_Display/n539 ),
    .i1(\u2_Display/n559 [17]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n574 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10340  (
    .i0(\u2_Display/n5351 ),
    .i1(\u2_Display/n5366 [12]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5386 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10341  (
    .i0(\u2_Display/n5352 ),
    .i1(\u2_Display/n5366 [11]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5387 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10342  (
    .i0(\u2_Display/n5353 ),
    .i1(\u2_Display/n5366 [10]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5388 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10343  (
    .i0(\u2_Display/n5354 ),
    .i1(\u2_Display/n5366 [9]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5389 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10344  (
    .i0(\u2_Display/n5355 ),
    .i1(\u2_Display/n5366 [8]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5390 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10345  (
    .i0(\u2_Display/n5356 ),
    .i1(\u2_Display/n5366 [7]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5391 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10346  (
    .i0(\u2_Display/n5357 ),
    .i1(\u2_Display/n5366 [6]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5392 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10347  (
    .i0(\u2_Display/n5358 ),
    .i1(\u2_Display/n5366 [5]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5393 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10348  (
    .i0(\u2_Display/n5359 ),
    .i1(\u2_Display/n5366 [4]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5394 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10349  (
    .i0(\u2_Display/n5360 ),
    .i1(\u2_Display/n5366 [3]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5395 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1035  (
    .i0(\u2_Display/n540 ),
    .i1(\u2_Display/n559 [16]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n575 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10350  (
    .i0(\u2_Display/n5361 ),
    .i1(\u2_Display/n5366 [2]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5396 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10351  (
    .i0(\u2_Display/n5362 ),
    .i1(\u2_Display/n5366 [1]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5397 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10352  (
    .i0(\u2_Display/n5363 ),
    .i1(\u2_Display/n5366 [0]),
    .sel(\u2_Display/n5365 ),
    .o(\u2_Display/n5398 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10353  (\u2_Display/n5400 , \u2_Display/n5399 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1036  (
    .i0(\u2_Display/n541 ),
    .i1(\u2_Display/n559 [15]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n576 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1037  (
    .i0(\u2_Display/n542 ),
    .i1(\u2_Display/n559 [14]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n577 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1038  (
    .i0(\u2_Display/n543 ),
    .i1(\u2_Display/n559 [13]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n578 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10386  (
    .i0(\u2_Display/n5367 ),
    .i1(\u2_Display/n5401 [31]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5402 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10387  (
    .i0(\u2_Display/n5368 ),
    .i1(\u2_Display/n5401 [30]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5403 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10388  (
    .i0(\u2_Display/n5369 ),
    .i1(\u2_Display/n5401 [29]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5404 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10389  (
    .i0(\u2_Display/n5370 ),
    .i1(\u2_Display/n5401 [28]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5405 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1039  (
    .i0(\u2_Display/n544 ),
    .i1(\u2_Display/n559 [12]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n579 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10390  (
    .i0(\u2_Display/n5371 ),
    .i1(\u2_Display/n5401 [27]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5406 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10391  (
    .i0(\u2_Display/n5372 ),
    .i1(\u2_Display/n5401 [26]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5407 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10392  (
    .i0(\u2_Display/n5373 ),
    .i1(\u2_Display/n5401 [25]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5408 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10393  (
    .i0(\u2_Display/n5374 ),
    .i1(\u2_Display/n5401 [24]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5409 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10394  (
    .i0(\u2_Display/n5375 ),
    .i1(\u2_Display/n5401 [23]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5410 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10395  (
    .i0(\u2_Display/n5376 ),
    .i1(\u2_Display/n5401 [22]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5411 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10396  (
    .i0(\u2_Display/n5377 ),
    .i1(\u2_Display/n5401 [21]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5412 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10397  (
    .i0(\u2_Display/n5378 ),
    .i1(\u2_Display/n5401 [20]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5413 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10398  (
    .i0(\u2_Display/n5379 ),
    .i1(\u2_Display/n5401 [19]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5414 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10399  (
    .i0(\u2_Display/n5380 ),
    .i1(\u2_Display/n5401 [18]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5415 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1040  (
    .i0(\u2_Display/n545 ),
    .i1(\u2_Display/n559 [11]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n580 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10400  (
    .i0(\u2_Display/n5381 ),
    .i1(\u2_Display/n5401 [17]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5416 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10401  (
    .i0(\u2_Display/n5382 ),
    .i1(\u2_Display/n5401 [16]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5417 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10402  (
    .i0(\u2_Display/n5383 ),
    .i1(\u2_Display/n5401 [15]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5418 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10403  (
    .i0(\u2_Display/n5384 ),
    .i1(\u2_Display/n5401 [14]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5419 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10404  (
    .i0(\u2_Display/n5385 ),
    .i1(\u2_Display/n5401 [13]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5420 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10405  (
    .i0(\u2_Display/n5386 ),
    .i1(\u2_Display/n5401 [12]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5421 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10406  (
    .i0(\u2_Display/n5387 ),
    .i1(\u2_Display/n5401 [11]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5422 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10407  (
    .i0(\u2_Display/n5388 ),
    .i1(\u2_Display/n5401 [10]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5423 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10408  (
    .i0(\u2_Display/n5389 ),
    .i1(\u2_Display/n5401 [9]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5424 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10409  (
    .i0(\u2_Display/n5390 ),
    .i1(\u2_Display/n5401 [8]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5425 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1041  (
    .i0(\u2_Display/n546 ),
    .i1(\u2_Display/n559 [10]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n581 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10410  (
    .i0(\u2_Display/n5391 ),
    .i1(\u2_Display/n5401 [7]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5426 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10411  (
    .i0(\u2_Display/n5392 ),
    .i1(\u2_Display/n5401 [6]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5427 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10412  (
    .i0(\u2_Display/n5393 ),
    .i1(\u2_Display/n5401 [5]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5428 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10413  (
    .i0(\u2_Display/n5394 ),
    .i1(\u2_Display/n5401 [4]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5429 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10414  (
    .i0(\u2_Display/n5395 ),
    .i1(\u2_Display/n5401 [3]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5430 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10415  (
    .i0(\u2_Display/n5396 ),
    .i1(\u2_Display/n5401 [2]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5431 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10416  (
    .i0(\u2_Display/n5397 ),
    .i1(\u2_Display/n5401 [1]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5432 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10417  (
    .i0(\u2_Display/n5398 ),
    .i1(\u2_Display/n5401 [0]),
    .sel(\u2_Display/n5400 ),
    .o(\u2_Display/n5433 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10418  (\u2_Display/n5435 , \u2_Display/n5434 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1042  (
    .i0(\u2_Display/n547 ),
    .i1(\u2_Display/n559 [9]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n582 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1043  (
    .i0(\u2_Display/n548 ),
    .i1(\u2_Display/n559 [8]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n583 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1044  (
    .i0(\u2_Display/n549 ),
    .i1(\u2_Display/n559 [7]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n584 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1045  (
    .i0(\u2_Display/n550 ),
    .i1(\u2_Display/n559 [6]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n585 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10451  (
    .i0(\u2_Display/n5402 ),
    .i1(\u2_Display/n5436 [31]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5437 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10452  (
    .i0(\u2_Display/n5403 ),
    .i1(\u2_Display/n5436 [30]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5438 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10453  (
    .i0(\u2_Display/n5404 ),
    .i1(\u2_Display/n5436 [29]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5439 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10454  (
    .i0(\u2_Display/n5405 ),
    .i1(\u2_Display/n5436 [28]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5440 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10455  (
    .i0(\u2_Display/n5406 ),
    .i1(\u2_Display/n5436 [27]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5441 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10456  (
    .i0(\u2_Display/n5407 ),
    .i1(\u2_Display/n5436 [26]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5442 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10457  (
    .i0(\u2_Display/n5408 ),
    .i1(\u2_Display/n5436 [25]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5443 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10458  (
    .i0(\u2_Display/n5409 ),
    .i1(\u2_Display/n5436 [24]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5444 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10459  (
    .i0(\u2_Display/n5410 ),
    .i1(\u2_Display/n5436 [23]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5445 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1046  (
    .i0(\u2_Display/n551 ),
    .i1(\u2_Display/n559 [5]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n586 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10460  (
    .i0(\u2_Display/n5411 ),
    .i1(\u2_Display/n5436 [22]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5446 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10461  (
    .i0(\u2_Display/n5412 ),
    .i1(\u2_Display/n5436 [21]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5447 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10462  (
    .i0(\u2_Display/n5413 ),
    .i1(\u2_Display/n5436 [20]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5448 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10463  (
    .i0(\u2_Display/n5414 ),
    .i1(\u2_Display/n5436 [19]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5449 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10464  (
    .i0(\u2_Display/n5415 ),
    .i1(\u2_Display/n5436 [18]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5450 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10465  (
    .i0(\u2_Display/n5416 ),
    .i1(\u2_Display/n5436 [17]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5451 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10466  (
    .i0(\u2_Display/n5417 ),
    .i1(\u2_Display/n5436 [16]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5452 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10467  (
    .i0(\u2_Display/n5418 ),
    .i1(\u2_Display/n5436 [15]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5453 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10468  (
    .i0(\u2_Display/n5419 ),
    .i1(\u2_Display/n5436 [14]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5454 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10469  (
    .i0(\u2_Display/n5420 ),
    .i1(\u2_Display/n5436 [13]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5455 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1047  (
    .i0(\u2_Display/n552 ),
    .i1(\u2_Display/n559 [4]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n587 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10470  (
    .i0(\u2_Display/n5421 ),
    .i1(\u2_Display/n5436 [12]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5456 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10471  (
    .i0(\u2_Display/n5422 ),
    .i1(\u2_Display/n5436 [11]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5457 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10472  (
    .i0(\u2_Display/n5423 ),
    .i1(\u2_Display/n5436 [10]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5458 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10473  (
    .i0(\u2_Display/n5424 ),
    .i1(\u2_Display/n5436 [9]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5459 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10474  (
    .i0(\u2_Display/n5425 ),
    .i1(\u2_Display/n5436 [8]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5460 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10475  (
    .i0(\u2_Display/n5426 ),
    .i1(\u2_Display/n5436 [7]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5461 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10476  (
    .i0(\u2_Display/n5427 ),
    .i1(\u2_Display/n5436 [6]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5462 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10477  (
    .i0(\u2_Display/n5428 ),
    .i1(\u2_Display/n5436 [5]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5463 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10478  (
    .i0(\u2_Display/n5429 ),
    .i1(\u2_Display/n5436 [4]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5464 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10479  (
    .i0(\u2_Display/n5430 ),
    .i1(\u2_Display/n5436 [3]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5465 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1048  (
    .i0(\u2_Display/n553 ),
    .i1(\u2_Display/n559 [3]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n588 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10480  (
    .i0(\u2_Display/n5431 ),
    .i1(\u2_Display/n5436 [2]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5466 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10481  (
    .i0(\u2_Display/n5432 ),
    .i1(\u2_Display/n5436 [1]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5467 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10482  (
    .i0(\u2_Display/n5433 ),
    .i1(\u2_Display/n5436 [0]),
    .sel(\u2_Display/n5435 ),
    .o(\u2_Display/n5468 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10483  (\u2_Display/n5470 , \u2_Display/n5469 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1049  (
    .i0(\u2_Display/n554 ),
    .i1(\u2_Display/n559 [2]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n589 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1050  (
    .i0(\u2_Display/n555 ),
    .i1(\u2_Display/n559 [1]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n590 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1051  (
    .i0(\u2_Display/n556 ),
    .i1(\u2_Display/n559 [0]),
    .sel(\u2_Display/n558 ),
    .o(\u2_Display/n591 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10516  (
    .i0(\u2_Display/n5437 ),
    .i1(\u2_Display/n5471 [31]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5472 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10517  (
    .i0(\u2_Display/n5438 ),
    .i1(\u2_Display/n5471 [30]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5473 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10518  (
    .i0(\u2_Display/n5439 ),
    .i1(\u2_Display/n5471 [29]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5474 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10519  (
    .i0(\u2_Display/n5440 ),
    .i1(\u2_Display/n5471 [28]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5475 ));  // source/rtl/Display.v(179)
  not \u2_Display/u1052  (\u2_Display/n593 , \u2_Display/n592 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10520  (
    .i0(\u2_Display/n5441 ),
    .i1(\u2_Display/n5471 [27]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5476 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10521  (
    .i0(\u2_Display/n5442 ),
    .i1(\u2_Display/n5471 [26]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5477 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10522  (
    .i0(\u2_Display/n5443 ),
    .i1(\u2_Display/n5471 [25]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5478 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10523  (
    .i0(\u2_Display/n5444 ),
    .i1(\u2_Display/n5471 [24]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5479 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10524  (
    .i0(\u2_Display/n5445 ),
    .i1(\u2_Display/n5471 [23]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5480 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10525  (
    .i0(\u2_Display/n5446 ),
    .i1(\u2_Display/n5471 [22]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5481 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10526  (
    .i0(\u2_Display/n5447 ),
    .i1(\u2_Display/n5471 [21]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5482 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10527  (
    .i0(\u2_Display/n5448 ),
    .i1(\u2_Display/n5471 [20]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5483 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10528  (
    .i0(\u2_Display/n5449 ),
    .i1(\u2_Display/n5471 [19]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5484 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10529  (
    .i0(\u2_Display/n5450 ),
    .i1(\u2_Display/n5471 [18]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5485 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10530  (
    .i0(\u2_Display/n5451 ),
    .i1(\u2_Display/n5471 [17]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5486 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10531  (
    .i0(\u2_Display/n5452 ),
    .i1(\u2_Display/n5471 [16]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5487 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10532  (
    .i0(\u2_Display/n5453 ),
    .i1(\u2_Display/n5471 [15]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5488 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10533  (
    .i0(\u2_Display/n5454 ),
    .i1(\u2_Display/n5471 [14]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5489 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10534  (
    .i0(\u2_Display/n5455 ),
    .i1(\u2_Display/n5471 [13]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5490 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10535  (
    .i0(\u2_Display/n5456 ),
    .i1(\u2_Display/n5471 [12]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5491 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10536  (
    .i0(\u2_Display/n5457 ),
    .i1(\u2_Display/n5471 [11]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5492 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10537  (
    .i0(\u2_Display/n5458 ),
    .i1(\u2_Display/n5471 [10]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5493 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10538  (
    .i0(\u2_Display/n5459 ),
    .i1(\u2_Display/n5471 [9]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5494 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10539  (
    .i0(\u2_Display/n5460 ),
    .i1(\u2_Display/n5471 [8]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5495 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10540  (
    .i0(\u2_Display/n5461 ),
    .i1(\u2_Display/n5471 [7]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5496 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10541  (
    .i0(\u2_Display/n5462 ),
    .i1(\u2_Display/n5471 [6]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5497 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10542  (
    .i0(\u2_Display/n5463 ),
    .i1(\u2_Display/n5471 [5]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5498 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10543  (
    .i0(\u2_Display/n5464 ),
    .i1(\u2_Display/n5471 [4]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5499 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10544  (
    .i0(\u2_Display/n5465 ),
    .i1(\u2_Display/n5471 [3]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5500 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10545  (
    .i0(\u2_Display/n5466 ),
    .i1(\u2_Display/n5471 [2]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5501 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10546  (
    .i0(\u2_Display/n5467 ),
    .i1(\u2_Display/n5471 [1]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5502 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10547  (
    .i0(\u2_Display/n5468 ),
    .i1(\u2_Display/n5471 [0]),
    .sel(\u2_Display/n5470 ),
    .o(\u2_Display/n5503 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10548  (\u2_Display/n5505 , \u2_Display/n5504 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10581  (
    .i0(\u2_Display/n5472 ),
    .i1(\u2_Display/n5506 [31]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5507 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10582  (
    .i0(\u2_Display/n5473 ),
    .i1(\u2_Display/n5506 [30]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5508 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10583  (
    .i0(\u2_Display/n5474 ),
    .i1(\u2_Display/n5506 [29]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5509 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10584  (
    .i0(\u2_Display/n5475 ),
    .i1(\u2_Display/n5506 [28]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5510 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10585  (
    .i0(\u2_Display/n5476 ),
    .i1(\u2_Display/n5506 [27]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5511 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10586  (
    .i0(\u2_Display/n5477 ),
    .i1(\u2_Display/n5506 [26]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5512 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10587  (
    .i0(\u2_Display/n5478 ),
    .i1(\u2_Display/n5506 [25]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5513 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10588  (
    .i0(\u2_Display/n5479 ),
    .i1(\u2_Display/n5506 [24]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5514 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10589  (
    .i0(\u2_Display/n5480 ),
    .i1(\u2_Display/n5506 [23]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5515 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10590  (
    .i0(\u2_Display/n5481 ),
    .i1(\u2_Display/n5506 [22]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5516 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10591  (
    .i0(\u2_Display/n5482 ),
    .i1(\u2_Display/n5506 [21]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5517 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10592  (
    .i0(\u2_Display/n5483 ),
    .i1(\u2_Display/n5506 [20]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5518 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10593  (
    .i0(\u2_Display/n5484 ),
    .i1(\u2_Display/n5506 [19]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5519 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10594  (
    .i0(\u2_Display/n5485 ),
    .i1(\u2_Display/n5506 [18]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5520 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10595  (
    .i0(\u2_Display/n5486 ),
    .i1(\u2_Display/n5506 [17]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5521 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10596  (
    .i0(\u2_Display/n5487 ),
    .i1(\u2_Display/n5506 [16]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5522 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10597  (
    .i0(\u2_Display/n5488 ),
    .i1(\u2_Display/n5506 [15]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5523 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10598  (
    .i0(\u2_Display/n5489 ),
    .i1(\u2_Display/n5506 [14]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5524 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10599  (
    .i0(\u2_Display/n5490 ),
    .i1(\u2_Display/n5506 [13]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5525 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10600  (
    .i0(\u2_Display/n5491 ),
    .i1(\u2_Display/n5506 [12]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5526 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10601  (
    .i0(\u2_Display/n5492 ),
    .i1(\u2_Display/n5506 [11]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5527 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10602  (
    .i0(\u2_Display/n5493 ),
    .i1(\u2_Display/n5506 [10]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5528 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10603  (
    .i0(\u2_Display/n5494 ),
    .i1(\u2_Display/n5506 [9]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5529 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10604  (
    .i0(\u2_Display/n5495 ),
    .i1(\u2_Display/n5506 [8]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5530 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10605  (
    .i0(\u2_Display/n5496 ),
    .i1(\u2_Display/n5506 [7]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5531 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10606  (
    .i0(\u2_Display/n5497 ),
    .i1(\u2_Display/n5506 [6]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5532 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10607  (
    .i0(\u2_Display/n5498 ),
    .i1(\u2_Display/n5506 [5]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5533 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10608  (
    .i0(\u2_Display/n5499 ),
    .i1(\u2_Display/n5506 [4]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5534 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10609  (
    .i0(\u2_Display/n5500 ),
    .i1(\u2_Display/n5506 [3]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5535 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10610  (
    .i0(\u2_Display/n5501 ),
    .i1(\u2_Display/n5506 [2]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5536 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10611  (
    .i0(\u2_Display/n5502 ),
    .i1(\u2_Display/n5506 [1]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5537 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10612  (
    .i0(\u2_Display/n5503 ),
    .i1(\u2_Display/n5506 [0]),
    .sel(\u2_Display/n5505 ),
    .o(\u2_Display/n5538 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10613  (\u2_Display/n5540 , \u2_Display/n5539 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10646  (
    .i0(\u2_Display/n5507 ),
    .i1(\u2_Display/n5541 [31]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5542 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10647  (
    .i0(\u2_Display/n5508 ),
    .i1(\u2_Display/n5541 [30]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5543 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10648  (
    .i0(\u2_Display/n5509 ),
    .i1(\u2_Display/n5541 [29]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5544 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10649  (
    .i0(\u2_Display/n5510 ),
    .i1(\u2_Display/n5541 [28]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5545 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10650  (
    .i0(\u2_Display/n5511 ),
    .i1(\u2_Display/n5541 [27]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5546 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10651  (
    .i0(\u2_Display/n5512 ),
    .i1(\u2_Display/n5541 [26]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5547 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10652  (
    .i0(\u2_Display/n5513 ),
    .i1(\u2_Display/n5541 [25]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5548 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10653  (
    .i0(\u2_Display/n5514 ),
    .i1(\u2_Display/n5541 [24]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5549 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10654  (
    .i0(\u2_Display/n5515 ),
    .i1(\u2_Display/n5541 [23]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5550 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10655  (
    .i0(\u2_Display/n5516 ),
    .i1(\u2_Display/n5541 [22]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5551 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10656  (
    .i0(\u2_Display/n5517 ),
    .i1(\u2_Display/n5541 [21]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5552 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10657  (
    .i0(\u2_Display/n5518 ),
    .i1(\u2_Display/n5541 [20]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5553 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10658  (
    .i0(\u2_Display/n5519 ),
    .i1(\u2_Display/n5541 [19]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5554 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10659  (
    .i0(\u2_Display/n5520 ),
    .i1(\u2_Display/n5541 [18]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5555 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10660  (
    .i0(\u2_Display/n5521 ),
    .i1(\u2_Display/n5541 [17]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5556 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10661  (
    .i0(\u2_Display/n5522 ),
    .i1(\u2_Display/n5541 [16]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5557 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10662  (
    .i0(\u2_Display/n5523 ),
    .i1(\u2_Display/n5541 [15]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5558 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10663  (
    .i0(\u2_Display/n5524 ),
    .i1(\u2_Display/n5541 [14]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5559 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10664  (
    .i0(\u2_Display/n5525 ),
    .i1(\u2_Display/n5541 [13]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5560 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10665  (
    .i0(\u2_Display/n5526 ),
    .i1(\u2_Display/n5541 [12]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5561 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10666  (
    .i0(\u2_Display/n5527 ),
    .i1(\u2_Display/n5541 [11]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5562 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10667  (
    .i0(\u2_Display/n5528 ),
    .i1(\u2_Display/n5541 [10]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5563 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10668  (
    .i0(\u2_Display/n5529 ),
    .i1(\u2_Display/n5541 [9]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5564 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10669  (
    .i0(\u2_Display/n5530 ),
    .i1(\u2_Display/n5541 [8]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5565 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10670  (
    .i0(\u2_Display/n5531 ),
    .i1(\u2_Display/n5541 [7]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5566 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10671  (
    .i0(\u2_Display/n5532 ),
    .i1(\u2_Display/n5541 [6]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5567 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10672  (
    .i0(\u2_Display/n5533 ),
    .i1(\u2_Display/n5541 [5]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5568 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10673  (
    .i0(\u2_Display/n5534 ),
    .i1(\u2_Display/n5541 [4]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5569 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10674  (
    .i0(\u2_Display/n5535 ),
    .i1(\u2_Display/n5541 [3]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5570 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10675  (
    .i0(\u2_Display/n5536 ),
    .i1(\u2_Display/n5541 [2]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5571 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10676  (
    .i0(\u2_Display/n5537 ),
    .i1(\u2_Display/n5541 [1]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5572 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10677  (
    .i0(\u2_Display/n5538 ),
    .i1(\u2_Display/n5541 [0]),
    .sel(\u2_Display/n5540 ),
    .o(\u2_Display/n5573 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10678  (\u2_Display/n5575 , \u2_Display/n5574 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10711  (
    .i0(\u2_Display/n5542 ),
    .i1(\u2_Display/n5576 [31]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5577 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10712  (
    .i0(\u2_Display/n5543 ),
    .i1(\u2_Display/n5576 [30]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5578 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10713  (
    .i0(\u2_Display/n5544 ),
    .i1(\u2_Display/n5576 [29]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5579 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10714  (
    .i0(\u2_Display/n5545 ),
    .i1(\u2_Display/n5576 [28]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5580 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10715  (
    .i0(\u2_Display/n5546 ),
    .i1(\u2_Display/n5576 [27]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5581 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10716  (
    .i0(\u2_Display/n5547 ),
    .i1(\u2_Display/n5576 [26]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5582 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10717  (
    .i0(\u2_Display/n5548 ),
    .i1(\u2_Display/n5576 [25]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5583 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10718  (
    .i0(\u2_Display/n5549 ),
    .i1(\u2_Display/n5576 [24]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5584 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10719  (
    .i0(\u2_Display/n5550 ),
    .i1(\u2_Display/n5576 [23]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5585 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10720  (
    .i0(\u2_Display/n5551 ),
    .i1(\u2_Display/n5576 [22]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5586 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10721  (
    .i0(\u2_Display/n5552 ),
    .i1(\u2_Display/n5576 [21]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5587 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10722  (
    .i0(\u2_Display/n5553 ),
    .i1(\u2_Display/n5576 [20]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5588 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10723  (
    .i0(\u2_Display/n5554 ),
    .i1(\u2_Display/n5576 [19]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5589 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10724  (
    .i0(\u2_Display/n5555 ),
    .i1(\u2_Display/n5576 [18]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5590 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10725  (
    .i0(\u2_Display/n5556 ),
    .i1(\u2_Display/n5576 [17]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5591 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10726  (
    .i0(\u2_Display/n5557 ),
    .i1(\u2_Display/n5576 [16]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5592 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10727  (
    .i0(\u2_Display/n5558 ),
    .i1(\u2_Display/n5576 [15]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5593 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10728  (
    .i0(\u2_Display/n5559 ),
    .i1(\u2_Display/n5576 [14]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5594 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10729  (
    .i0(\u2_Display/n5560 ),
    .i1(\u2_Display/n5576 [13]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5595 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10730  (
    .i0(\u2_Display/n5561 ),
    .i1(\u2_Display/n5576 [12]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5596 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10731  (
    .i0(\u2_Display/n5562 ),
    .i1(\u2_Display/n5576 [11]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5597 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10732  (
    .i0(\u2_Display/n5563 ),
    .i1(\u2_Display/n5576 [10]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5598 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10733  (
    .i0(\u2_Display/n5564 ),
    .i1(\u2_Display/n5576 [9]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5599 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10734  (
    .i0(\u2_Display/n5565 ),
    .i1(\u2_Display/n5576 [8]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5600 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10735  (
    .i0(\u2_Display/n5566 ),
    .i1(\u2_Display/n5576 [7]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5601 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10736  (
    .i0(\u2_Display/n5567 ),
    .i1(\u2_Display/n5576 [6]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5602 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10737  (
    .i0(\u2_Display/n5568 ),
    .i1(\u2_Display/n5576 [5]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5603 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10738  (
    .i0(\u2_Display/n5569 ),
    .i1(\u2_Display/n5576 [4]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5604 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10739  (
    .i0(\u2_Display/n5570 ),
    .i1(\u2_Display/n5576 [3]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5605 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10740  (
    .i0(\u2_Display/n5571 ),
    .i1(\u2_Display/n5576 [2]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5606 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10741  (
    .i0(\u2_Display/n5572 ),
    .i1(\u2_Display/n5576 [1]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5607 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10742  (
    .i0(\u2_Display/n5573 ),
    .i1(\u2_Display/n5576 [0]),
    .sel(\u2_Display/n5575 ),
    .o(\u2_Display/n5608 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10743  (\u2_Display/n5610 , \u2_Display/n5609 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10776  (
    .i0(\u2_Display/n5577 ),
    .i1(\u2_Display/n5611 [31]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5612 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10777  (
    .i0(\u2_Display/n5578 ),
    .i1(\u2_Display/n5611 [30]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5613 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10778  (
    .i0(\u2_Display/n5579 ),
    .i1(\u2_Display/n5611 [29]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5614 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10779  (
    .i0(\u2_Display/n5580 ),
    .i1(\u2_Display/n5611 [28]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5615 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10780  (
    .i0(\u2_Display/n5581 ),
    .i1(\u2_Display/n5611 [27]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5616 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10781  (
    .i0(\u2_Display/n5582 ),
    .i1(\u2_Display/n5611 [26]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5617 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10782  (
    .i0(\u2_Display/n5583 ),
    .i1(\u2_Display/n5611 [25]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5618 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10783  (
    .i0(\u2_Display/n5584 ),
    .i1(\u2_Display/n5611 [24]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5619 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10784  (
    .i0(\u2_Display/n5585 ),
    .i1(\u2_Display/n5611 [23]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5620 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10785  (
    .i0(\u2_Display/n5586 ),
    .i1(\u2_Display/n5611 [22]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5621 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10786  (
    .i0(\u2_Display/n5587 ),
    .i1(\u2_Display/n5611 [21]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5622 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10787  (
    .i0(\u2_Display/n5588 ),
    .i1(\u2_Display/n5611 [20]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5623 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10788  (
    .i0(\u2_Display/n5589 ),
    .i1(\u2_Display/n5611 [19]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5624 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10789  (
    .i0(\u2_Display/n5590 ),
    .i1(\u2_Display/n5611 [18]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5625 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10790  (
    .i0(\u2_Display/n5591 ),
    .i1(\u2_Display/n5611 [17]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5626 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10791  (
    .i0(\u2_Display/n5592 ),
    .i1(\u2_Display/n5611 [16]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5627 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10792  (
    .i0(\u2_Display/n5593 ),
    .i1(\u2_Display/n5611 [15]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5628 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10793  (
    .i0(\u2_Display/n5594 ),
    .i1(\u2_Display/n5611 [14]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5629 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10794  (
    .i0(\u2_Display/n5595 ),
    .i1(\u2_Display/n5611 [13]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5630 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10795  (
    .i0(\u2_Display/n5596 ),
    .i1(\u2_Display/n5611 [12]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5631 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10796  (
    .i0(\u2_Display/n5597 ),
    .i1(\u2_Display/n5611 [11]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5632 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10797  (
    .i0(\u2_Display/n5598 ),
    .i1(\u2_Display/n5611 [10]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5633 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10798  (
    .i0(\u2_Display/n5599 ),
    .i1(\u2_Display/n5611 [9]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5634 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10799  (
    .i0(\u2_Display/n5600 ),
    .i1(\u2_Display/n5611 [8]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5635 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10800  (
    .i0(\u2_Display/n5601 ),
    .i1(\u2_Display/n5611 [7]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5636 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10801  (
    .i0(\u2_Display/n5602 ),
    .i1(\u2_Display/n5611 [6]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5637 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10802  (
    .i0(\u2_Display/n5603 ),
    .i1(\u2_Display/n5611 [5]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5638 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10803  (
    .i0(\u2_Display/n5604 ),
    .i1(\u2_Display/n5611 [4]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5639 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10804  (
    .i0(\u2_Display/n5605 ),
    .i1(\u2_Display/n5611 [3]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5640 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10805  (
    .i0(\u2_Display/n5606 ),
    .i1(\u2_Display/n5611 [2]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5641 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10806  (
    .i0(\u2_Display/n5607 ),
    .i1(\u2_Display/n5611 [1]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5642 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10807  (
    .i0(\u2_Display/n5608 ),
    .i1(\u2_Display/n5611 [0]),
    .sel(\u2_Display/n5610 ),
    .o(\u2_Display/n5643 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10808  (\u2_Display/n5645 , \u2_Display/n5644 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10841  (
    .i0(\u2_Display/n5612 ),
    .i1(\u2_Display/n5646 [31]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5647 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10842  (
    .i0(\u2_Display/n5613 ),
    .i1(\u2_Display/n5646 [30]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5648 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10843  (
    .i0(\u2_Display/n5614 ),
    .i1(\u2_Display/n5646 [29]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5649 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10844  (
    .i0(\u2_Display/n5615 ),
    .i1(\u2_Display/n5646 [28]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5650 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10845  (
    .i0(\u2_Display/n5616 ),
    .i1(\u2_Display/n5646 [27]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5651 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10846  (
    .i0(\u2_Display/n5617 ),
    .i1(\u2_Display/n5646 [26]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5652 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10847  (
    .i0(\u2_Display/n5618 ),
    .i1(\u2_Display/n5646 [25]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5653 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10848  (
    .i0(\u2_Display/n5619 ),
    .i1(\u2_Display/n5646 [24]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5654 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10849  (
    .i0(\u2_Display/n5620 ),
    .i1(\u2_Display/n5646 [23]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5655 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1085  (
    .i0(\u2_Display/n560 ),
    .i1(\u2_Display/n594 [31]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n595 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10850  (
    .i0(\u2_Display/n5621 ),
    .i1(\u2_Display/n5646 [22]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5656 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10851  (
    .i0(\u2_Display/n5622 ),
    .i1(\u2_Display/n5646 [21]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5657 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10852  (
    .i0(\u2_Display/n5623 ),
    .i1(\u2_Display/n5646 [20]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5658 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10853  (
    .i0(\u2_Display/n5624 ),
    .i1(\u2_Display/n5646 [19]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5659 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10854  (
    .i0(\u2_Display/n5625 ),
    .i1(\u2_Display/n5646 [18]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5660 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10855  (
    .i0(\u2_Display/n5626 ),
    .i1(\u2_Display/n5646 [17]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5661 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10856  (
    .i0(\u2_Display/n5627 ),
    .i1(\u2_Display/n5646 [16]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5662 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10857  (
    .i0(\u2_Display/n5628 ),
    .i1(\u2_Display/n5646 [15]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5663 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10858  (
    .i0(\u2_Display/n5629 ),
    .i1(\u2_Display/n5646 [14]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5664 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10859  (
    .i0(\u2_Display/n5630 ),
    .i1(\u2_Display/n5646 [13]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5665 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1086  (
    .i0(\u2_Display/n561 ),
    .i1(\u2_Display/n594 [30]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n596 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10860  (
    .i0(\u2_Display/n5631 ),
    .i1(\u2_Display/n5646 [12]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5666 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10861  (
    .i0(\u2_Display/n5632 ),
    .i1(\u2_Display/n5646 [11]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5667 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10862  (
    .i0(\u2_Display/n5633 ),
    .i1(\u2_Display/n5646 [10]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5668 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10863  (
    .i0(\u2_Display/n5634 ),
    .i1(\u2_Display/n5646 [9]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5669 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10864  (
    .i0(\u2_Display/n5635 ),
    .i1(\u2_Display/n5646 [8]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5670 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10865  (
    .i0(\u2_Display/n5636 ),
    .i1(\u2_Display/n5646 [7]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5671 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10866  (
    .i0(\u2_Display/n5637 ),
    .i1(\u2_Display/n5646 [6]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5672 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10867  (
    .i0(\u2_Display/n5638 ),
    .i1(\u2_Display/n5646 [5]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5673 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10868  (
    .i0(\u2_Display/n5639 ),
    .i1(\u2_Display/n5646 [4]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5674 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10869  (
    .i0(\u2_Display/n5640 ),
    .i1(\u2_Display/n5646 [3]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5675 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1087  (
    .i0(\u2_Display/n562 ),
    .i1(\u2_Display/n594 [29]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n597 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10870  (
    .i0(\u2_Display/n5641 ),
    .i1(\u2_Display/n5646 [2]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5676 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10871  (
    .i0(\u2_Display/n5642 ),
    .i1(\u2_Display/n5646 [1]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5677 ));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10872  (
    .i0(\u2_Display/n5643 ),
    .i1(\u2_Display/n5646 [0]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n5678 ));  // source/rtl/Display.v(179)
  not \u2_Display/u10873  (\u2_Display/n5680 , \u2_Display/n5679 );  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1088  (
    .i0(\u2_Display/n563 ),
    .i1(\u2_Display/n594 [28]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n598 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1089  (
    .i0(\u2_Display/n564 ),
    .i1(\u2_Display/n594 [27]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n599 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1090  (
    .i0(\u2_Display/n565 ),
    .i1(\u2_Display/n594 [26]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n600 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10906  (
    .i0(\u2_Display/n5669 ),
    .i1(\u2_Display/n5681 [9]),
    .sel(\u2_Display/n5680 ),
    .o(\u2_Display/n93 [9]));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10907  (
    .i0(\u2_Display/n5670 ),
    .i1(\u2_Display/n5681 [8]),
    .sel(\u2_Display/n5680 ),
    .o(\u2_Display/n93 [8]));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10908  (
    .i0(\u2_Display/n5671 ),
    .i1(\u2_Display/n5681 [7]),
    .sel(\u2_Display/n5680 ),
    .o(\u2_Display/n93 [7]));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10909  (
    .i0(\u2_Display/n5672 ),
    .i1(\u2_Display/n5681 [6]),
    .sel(\u2_Display/n5680 ),
    .o(\u2_Display/n93 [6]));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1091  (
    .i0(\u2_Display/n566 ),
    .i1(\u2_Display/n594 [25]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n601 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u10910  (
    .i0(\u2_Display/n5673 ),
    .i1(\u2_Display/n5681 [5]),
    .sel(\u2_Display/n5680 ),
    .o(\u2_Display/n93 [5]));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10911  (
    .i0(\u2_Display/n5674 ),
    .i1(\u2_Display/n5681 [4]),
    .sel(\u2_Display/n5680 ),
    .o(\u2_Display/n93 [4]));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10912  (
    .i0(\u2_Display/n5675 ),
    .i1(\u2_Display/n5681 [3]),
    .sel(\u2_Display/n5680 ),
    .o(\u2_Display/n93 [3]));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10913  (
    .i0(\u2_Display/n5676 ),
    .i1(\u2_Display/n5681 [2]),
    .sel(\u2_Display/n5680 ),
    .o(\u2_Display/n93 [2]));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10914  (
    .i0(\u2_Display/n5677 ),
    .i1(\u2_Display/n5681 [1]),
    .sel(\u2_Display/n5680 ),
    .o(\u2_Display/n93 [1]));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u10915  (
    .i0(\u2_Display/n5678 ),
    .i1(\u2_Display/n5681 [0]),
    .sel(\u2_Display/n5680 ),
    .o(\u2_Display/n93 [0]));  // source/rtl/Display.v(179)
  AL_MUX \u2_Display/u1092  (
    .i0(\u2_Display/n567 ),
    .i1(\u2_Display/n594 [24]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n602 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1093  (
    .i0(\u2_Display/n568 ),
    .i1(\u2_Display/n594 [23]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n603 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1094  (
    .i0(\u2_Display/n569 ),
    .i1(\u2_Display/n594 [22]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n604 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1095  (
    .i0(\u2_Display/n570 ),
    .i1(\u2_Display/n594 [21]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n605 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1096  (
    .i0(\u2_Display/n571 ),
    .i1(\u2_Display/n594 [20]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n606 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1097  (
    .i0(\u2_Display/n572 ),
    .i1(\u2_Display/n594 [19]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n607 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1098  (
    .i0(\u2_Display/n573 ),
    .i1(\u2_Display/n594 [18]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n608 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1099  (
    .i0(\u2_Display/n574 ),
    .i1(\u2_Display/n594 [17]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n609 ));  // source/rtl/Display.v(230)
  and \u2_Display/u11  (\u2_Display/n51 , \u2_Display/n49 , \u2_Display/n50 );  // source/rtl/Display.v(165)
  AL_MUX \u2_Display/u1100  (
    .i0(\u2_Display/n575 ),
    .i1(\u2_Display/n594 [16]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n610 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1101  (
    .i0(\u2_Display/n576 ),
    .i1(\u2_Display/n594 [15]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n611 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1102  (
    .i0(\u2_Display/n577 ),
    .i1(\u2_Display/n594 [14]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n612 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1103  (
    .i0(\u2_Display/n578 ),
    .i1(\u2_Display/n594 [13]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n613 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1104  (
    .i0(\u2_Display/n579 ),
    .i1(\u2_Display/n594 [12]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n614 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1105  (
    .i0(\u2_Display/n580 ),
    .i1(\u2_Display/n594 [11]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n615 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1106  (
    .i0(\u2_Display/n581 ),
    .i1(\u2_Display/n594 [10]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n616 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1107  (
    .i0(\u2_Display/n582 ),
    .i1(\u2_Display/n594 [9]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n617 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1108  (
    .i0(\u2_Display/n583 ),
    .i1(\u2_Display/n594 [8]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n618 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1109  (
    .i0(\u2_Display/n584 ),
    .i1(\u2_Display/n594 [7]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n619 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1110  (
    .i0(\u2_Display/n585 ),
    .i1(\u2_Display/n594 [6]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n620 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1111  (
    .i0(\u2_Display/n586 ),
    .i1(\u2_Display/n594 [5]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n621 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1112  (
    .i0(\u2_Display/n587 ),
    .i1(\u2_Display/n594 [4]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n622 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1113  (
    .i0(\u2_Display/n588 ),
    .i1(\u2_Display/n594 [3]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n623 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1114  (
    .i0(\u2_Display/n589 ),
    .i1(\u2_Display/n594 [2]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n624 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1115  (
    .i0(\u2_Display/n590 ),
    .i1(\u2_Display/n594 [1]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n625 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1116  (
    .i0(\u2_Display/n591 ),
    .i1(\u2_Display/n594 [0]),
    .sel(\u2_Display/n593 ),
    .o(\u2_Display/n626 ));  // source/rtl/Display.v(230)
  not \u2_Display/u1117  (\u2_Display/n628 , \u2_Display/n627 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1150  (
    .i0(\u2_Display/n595 ),
    .i1(\u2_Display/n629 [31]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n630 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1151  (
    .i0(\u2_Display/n596 ),
    .i1(\u2_Display/n629 [30]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n631 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1152  (
    .i0(\u2_Display/n597 ),
    .i1(\u2_Display/n629 [29]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n632 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1153  (
    .i0(\u2_Display/n598 ),
    .i1(\u2_Display/n629 [28]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n633 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1154  (
    .i0(\u2_Display/n599 ),
    .i1(\u2_Display/n629 [27]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n634 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1155  (
    .i0(\u2_Display/n600 ),
    .i1(\u2_Display/n629 [26]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n635 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1156  (
    .i0(\u2_Display/n601 ),
    .i1(\u2_Display/n629 [25]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n636 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1157  (
    .i0(\u2_Display/n602 ),
    .i1(\u2_Display/n629 [24]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n637 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1158  (
    .i0(\u2_Display/n603 ),
    .i1(\u2_Display/n629 [23]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n638 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1159  (
    .i0(\u2_Display/n604 ),
    .i1(\u2_Display/n629 [22]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n639 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1160  (
    .i0(\u2_Display/n605 ),
    .i1(\u2_Display/n629 [21]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n640 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1161  (
    .i0(\u2_Display/n606 ),
    .i1(\u2_Display/n629 [20]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n641 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1162  (
    .i0(\u2_Display/n607 ),
    .i1(\u2_Display/n629 [19]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n642 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1163  (
    .i0(\u2_Display/n608 ),
    .i1(\u2_Display/n629 [18]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n643 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1164  (
    .i0(\u2_Display/n609 ),
    .i1(\u2_Display/n629 [17]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n644 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1165  (
    .i0(\u2_Display/n610 ),
    .i1(\u2_Display/n629 [16]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n645 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1166  (
    .i0(\u2_Display/n611 ),
    .i1(\u2_Display/n629 [15]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n646 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1167  (
    .i0(\u2_Display/n612 ),
    .i1(\u2_Display/n629 [14]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n647 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1168  (
    .i0(\u2_Display/n613 ),
    .i1(\u2_Display/n629 [13]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n648 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1169  (
    .i0(\u2_Display/n614 ),
    .i1(\u2_Display/n629 [12]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n649 ));  // source/rtl/Display.v(230)
  not \u2_Display/u11698  (\u2_Display/n6068 , \u2_Display/n4909 );  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1170  (
    .i0(\u2_Display/n615 ),
    .i1(\u2_Display/n629 [11]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n650 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1171  (
    .i0(\u2_Display/n616 ),
    .i1(\u2_Display/n629 [10]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n651 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1172  (
    .i0(\u2_Display/n617 ),
    .i1(\u2_Display/n629 [9]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n652 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1173  (
    .i0(\u2_Display/n618 ),
    .i1(\u2_Display/n629 [8]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n653 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u11731  (
    .i0(\u2_Display/counta [31]),
    .i1(\u2_Display/n4911 [31]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6070 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11732  (
    .i0(\u2_Display/counta [30]),
    .i1(\u2_Display/n4911 [30]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6071 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11733  (
    .i0(\u2_Display/counta [29]),
    .i1(\u2_Display/n4911 [29]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6072 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11734  (
    .i0(\u2_Display/counta [28]),
    .i1(\u2_Display/n4911 [28]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6073 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11735  (
    .i0(\u2_Display/counta [27]),
    .i1(\u2_Display/n4911 [27]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6074 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11736  (
    .i0(\u2_Display/counta [26]),
    .i1(\u2_Display/n4911 [26]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6075 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11737  (
    .i0(\u2_Display/counta [25]),
    .i1(\u2_Display/n4911 [25]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6076 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11738  (
    .i0(\u2_Display/counta [24]),
    .i1(\u2_Display/n4911 [24]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6077 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11739  (
    .i0(\u2_Display/counta [23]),
    .i1(\u2_Display/n4911 [23]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6078 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1174  (
    .i0(\u2_Display/n619 ),
    .i1(\u2_Display/n629 [7]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n654 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u11740  (
    .i0(\u2_Display/counta [22]),
    .i1(\u2_Display/n4911 [22]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6079 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11741  (
    .i0(\u2_Display/counta [21]),
    .i1(\u2_Display/n4911 [21]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6080 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11742  (
    .i0(\u2_Display/counta [20]),
    .i1(\u2_Display/n4911 [20]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6081 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11743  (
    .i0(\u2_Display/counta [19]),
    .i1(\u2_Display/n4911 [19]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6082 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11744  (
    .i0(\u2_Display/counta [18]),
    .i1(\u2_Display/n4911 [18]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6083 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11745  (
    .i0(\u2_Display/counta [17]),
    .i1(\u2_Display/n4911 [17]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6084 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11746  (
    .i0(\u2_Display/counta [16]),
    .i1(\u2_Display/n4911 [16]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6085 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11747  (
    .i0(\u2_Display/counta [15]),
    .i1(\u2_Display/n4911 [15]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6086 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11748  (
    .i0(\u2_Display/counta [14]),
    .i1(\u2_Display/n4911 [14]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6087 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11749  (
    .i0(\u2_Display/counta [13]),
    .i1(\u2_Display/n4911 [13]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6088 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1175  (
    .i0(\u2_Display/n620 ),
    .i1(\u2_Display/n629 [6]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n655 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u11750  (
    .i0(\u2_Display/counta [12]),
    .i1(\u2_Display/n4911 [12]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6089 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11751  (
    .i0(\u2_Display/counta [11]),
    .i1(\u2_Display/n4911 [11]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6090 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11752  (
    .i0(\u2_Display/counta [10]),
    .i1(\u2_Display/n4911 [10]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6091 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11753  (
    .i0(\u2_Display/counta [9]),
    .i1(\u2_Display/n4911 [9]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6092 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11754  (
    .i0(\u2_Display/counta [8]),
    .i1(\u2_Display/n4911 [8]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6093 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11755  (
    .i0(\u2_Display/counta [7]),
    .i1(\u2_Display/n4911 [7]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6094 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11756  (
    .i0(\u2_Display/counta [6]),
    .i1(\u2_Display/n4911 [6]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6095 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11757  (
    .i0(\u2_Display/counta [5]),
    .i1(\u2_Display/n4911 [5]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6096 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11758  (
    .i0(\u2_Display/counta [4]),
    .i1(\u2_Display/n4911 [4]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6097 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11759  (
    .i0(\u2_Display/counta [3]),
    .i1(\u2_Display/n4911 [3]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6098 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1176  (
    .i0(\u2_Display/n621 ),
    .i1(\u2_Display/n629 [5]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n656 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u11760  (
    .i0(\u2_Display/counta [2]),
    .i1(\u2_Display/n4911 [2]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6099 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11761  (
    .i0(\u2_Display/counta [1]),
    .i1(\u2_Display/n4911 [1]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6100 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11762  (
    .i0(\u2_Display/counta [0]),
    .i1(\u2_Display/n4911 [0]),
    .sel(\u2_Display/n6068 ),
    .o(\u2_Display/n6101 ));  // source/rtl/Display.v(163)
  not \u2_Display/u11763  (\u2_Display/n6103 , \u2_Display/n4944 );  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1177  (
    .i0(\u2_Display/n622 ),
    .i1(\u2_Display/n629 [4]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n657 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1178  (
    .i0(\u2_Display/n623 ),
    .i1(\u2_Display/n629 [3]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n658 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1179  (
    .i0(\u2_Display/n624 ),
    .i1(\u2_Display/n629 [2]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n659 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u11796  (
    .i0(\u2_Display/n6070 ),
    .i1(\u2_Display/n4946 [31]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6105 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11797  (
    .i0(\u2_Display/n6071 ),
    .i1(\u2_Display/n4946 [30]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6106 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11798  (
    .i0(\u2_Display/n6072 ),
    .i1(\u2_Display/n4946 [29]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6107 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11799  (
    .i0(\u2_Display/n6073 ),
    .i1(\u2_Display/n4946 [28]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6108 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1180  (
    .i0(\u2_Display/n625 ),
    .i1(\u2_Display/n629 [1]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n660 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u11800  (
    .i0(\u2_Display/n6074 ),
    .i1(\u2_Display/n4946 [27]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6109 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11801  (
    .i0(\u2_Display/n6075 ),
    .i1(\u2_Display/n4946 [26]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6110 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11802  (
    .i0(\u2_Display/n6076 ),
    .i1(\u2_Display/n4946 [25]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6111 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11803  (
    .i0(\u2_Display/n6077 ),
    .i1(\u2_Display/n4946 [24]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6112 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11804  (
    .i0(\u2_Display/n6078 ),
    .i1(\u2_Display/n4946 [23]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6113 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11805  (
    .i0(\u2_Display/n6079 ),
    .i1(\u2_Display/n4946 [22]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6114 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11806  (
    .i0(\u2_Display/n6080 ),
    .i1(\u2_Display/n4946 [21]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6115 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11807  (
    .i0(\u2_Display/n6081 ),
    .i1(\u2_Display/n4946 [20]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6116 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11808  (
    .i0(\u2_Display/n6082 ),
    .i1(\u2_Display/n4946 [19]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6117 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11809  (
    .i0(\u2_Display/n6083 ),
    .i1(\u2_Display/n4946 [18]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6118 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1181  (
    .i0(\u2_Display/n626 ),
    .i1(\u2_Display/n629 [0]),
    .sel(\u2_Display/n628 ),
    .o(\u2_Display/n661 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u11810  (
    .i0(\u2_Display/n6084 ),
    .i1(\u2_Display/n4946 [17]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6119 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11811  (
    .i0(\u2_Display/n6085 ),
    .i1(\u2_Display/n4946 [16]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6120 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11812  (
    .i0(\u2_Display/n6086 ),
    .i1(\u2_Display/n4946 [15]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6121 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11813  (
    .i0(\u2_Display/n6087 ),
    .i1(\u2_Display/n4946 [14]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6122 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11814  (
    .i0(\u2_Display/n6088 ),
    .i1(\u2_Display/n4946 [13]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6123 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11815  (
    .i0(\u2_Display/n6089 ),
    .i1(\u2_Display/n4946 [12]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6124 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11816  (
    .i0(\u2_Display/n6090 ),
    .i1(\u2_Display/n4946 [11]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6125 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11817  (
    .i0(\u2_Display/n6091 ),
    .i1(\u2_Display/n4946 [10]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6126 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11818  (
    .i0(\u2_Display/n6092 ),
    .i1(\u2_Display/n4946 [9]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6127 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11819  (
    .i0(\u2_Display/n6093 ),
    .i1(\u2_Display/n4946 [8]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6128 ));  // source/rtl/Display.v(163)
  not \u2_Display/u1182  (\u2_Display/n663 , \u2_Display/n662 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u11820  (
    .i0(\u2_Display/n6094 ),
    .i1(\u2_Display/n4946 [7]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6129 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11821  (
    .i0(\u2_Display/n6095 ),
    .i1(\u2_Display/n4946 [6]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6130 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11822  (
    .i0(\u2_Display/n6096 ),
    .i1(\u2_Display/n4946 [5]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6131 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11823  (
    .i0(\u2_Display/n6097 ),
    .i1(\u2_Display/n4946 [4]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6132 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11824  (
    .i0(\u2_Display/n6098 ),
    .i1(\u2_Display/n4946 [3]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6133 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11825  (
    .i0(\u2_Display/n6099 ),
    .i1(\u2_Display/n4946 [2]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6134 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11826  (
    .i0(\u2_Display/n6100 ),
    .i1(\u2_Display/n4946 [1]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6135 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11827  (
    .i0(\u2_Display/n6101 ),
    .i1(\u2_Display/n4946 [0]),
    .sel(\u2_Display/n6103 ),
    .o(\u2_Display/n6136 ));  // source/rtl/Display.v(163)
  not \u2_Display/u11828  (\u2_Display/n6138 , \u2_Display/n4979 );  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11861  (
    .i0(\u2_Display/n6105 ),
    .i1(\u2_Display/n4981 [31]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6140 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11862  (
    .i0(\u2_Display/n6106 ),
    .i1(\u2_Display/n4981 [30]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6141 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11863  (
    .i0(\u2_Display/n6107 ),
    .i1(\u2_Display/n4981 [29]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6142 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11864  (
    .i0(\u2_Display/n6108 ),
    .i1(\u2_Display/n4981 [28]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6143 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11865  (
    .i0(\u2_Display/n6109 ),
    .i1(\u2_Display/n4981 [27]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6144 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11866  (
    .i0(\u2_Display/n6110 ),
    .i1(\u2_Display/n4981 [26]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6145 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11867  (
    .i0(\u2_Display/n6111 ),
    .i1(\u2_Display/n4981 [25]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6146 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11868  (
    .i0(\u2_Display/n6112 ),
    .i1(\u2_Display/n4981 [24]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6147 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11869  (
    .i0(\u2_Display/n6113 ),
    .i1(\u2_Display/n4981 [23]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6148 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11870  (
    .i0(\u2_Display/n6114 ),
    .i1(\u2_Display/n4981 [22]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6149 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11871  (
    .i0(\u2_Display/n6115 ),
    .i1(\u2_Display/n4981 [21]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6150 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11872  (
    .i0(\u2_Display/n6116 ),
    .i1(\u2_Display/n4981 [20]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6151 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11873  (
    .i0(\u2_Display/n6117 ),
    .i1(\u2_Display/n4981 [19]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6152 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11874  (
    .i0(\u2_Display/n6118 ),
    .i1(\u2_Display/n4981 [18]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6153 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11875  (
    .i0(\u2_Display/n6119 ),
    .i1(\u2_Display/n4981 [17]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6154 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11876  (
    .i0(\u2_Display/n6120 ),
    .i1(\u2_Display/n4981 [16]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6155 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11877  (
    .i0(\u2_Display/n6121 ),
    .i1(\u2_Display/n4981 [15]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6156 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11878  (
    .i0(\u2_Display/n6122 ),
    .i1(\u2_Display/n4981 [14]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6157 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11879  (
    .i0(\u2_Display/n6123 ),
    .i1(\u2_Display/n4981 [13]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6158 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11880  (
    .i0(\u2_Display/n6124 ),
    .i1(\u2_Display/n4981 [12]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6159 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11881  (
    .i0(\u2_Display/n6125 ),
    .i1(\u2_Display/n4981 [11]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6160 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11882  (
    .i0(\u2_Display/n6126 ),
    .i1(\u2_Display/n4981 [10]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6161 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11883  (
    .i0(\u2_Display/n6127 ),
    .i1(\u2_Display/n4981 [9]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6162 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11884  (
    .i0(\u2_Display/n6128 ),
    .i1(\u2_Display/n4981 [8]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6163 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11885  (
    .i0(\u2_Display/n6129 ),
    .i1(\u2_Display/n4981 [7]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6164 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11886  (
    .i0(\u2_Display/n6130 ),
    .i1(\u2_Display/n4981 [6]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6165 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11887  (
    .i0(\u2_Display/n6131 ),
    .i1(\u2_Display/n4981 [5]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6166 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11888  (
    .i0(\u2_Display/n6132 ),
    .i1(\u2_Display/n4981 [4]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6167 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11889  (
    .i0(\u2_Display/n6133 ),
    .i1(\u2_Display/n4981 [3]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6168 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11890  (
    .i0(\u2_Display/n6134 ),
    .i1(\u2_Display/n4981 [2]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6169 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11891  (
    .i0(\u2_Display/n6135 ),
    .i1(\u2_Display/n4981 [1]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6170 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11892  (
    .i0(\u2_Display/n6136 ),
    .i1(\u2_Display/n4981 [0]),
    .sel(\u2_Display/n6138 ),
    .o(\u2_Display/n6171 ));  // source/rtl/Display.v(163)
  not \u2_Display/u11893  (\u2_Display/n6173 , \u2_Display/n5014 );  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11926  (
    .i0(\u2_Display/n6140 ),
    .i1(\u2_Display/n5016 [31]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6175 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11927  (
    .i0(\u2_Display/n6141 ),
    .i1(\u2_Display/n5016 [30]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6176 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11928  (
    .i0(\u2_Display/n6142 ),
    .i1(\u2_Display/n5016 [29]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6177 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11929  (
    .i0(\u2_Display/n6143 ),
    .i1(\u2_Display/n5016 [28]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6178 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11930  (
    .i0(\u2_Display/n6144 ),
    .i1(\u2_Display/n5016 [27]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6179 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11931  (
    .i0(\u2_Display/n6145 ),
    .i1(\u2_Display/n5016 [26]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6180 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11932  (
    .i0(\u2_Display/n6146 ),
    .i1(\u2_Display/n5016 [25]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6181 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11933  (
    .i0(\u2_Display/n6147 ),
    .i1(\u2_Display/n5016 [24]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6182 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11934  (
    .i0(\u2_Display/n6148 ),
    .i1(\u2_Display/n5016 [23]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6183 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11935  (
    .i0(\u2_Display/n6149 ),
    .i1(\u2_Display/n5016 [22]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6184 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11936  (
    .i0(\u2_Display/n6150 ),
    .i1(\u2_Display/n5016 [21]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6185 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11937  (
    .i0(\u2_Display/n6151 ),
    .i1(\u2_Display/n5016 [20]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6186 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11938  (
    .i0(\u2_Display/n6152 ),
    .i1(\u2_Display/n5016 [19]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6187 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11939  (
    .i0(\u2_Display/n6153 ),
    .i1(\u2_Display/n5016 [18]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6188 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11940  (
    .i0(\u2_Display/n6154 ),
    .i1(\u2_Display/n5016 [17]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6189 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11941  (
    .i0(\u2_Display/n6155 ),
    .i1(\u2_Display/n5016 [16]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6190 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11942  (
    .i0(\u2_Display/n6156 ),
    .i1(\u2_Display/n5016 [15]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6191 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11943  (
    .i0(\u2_Display/n6157 ),
    .i1(\u2_Display/n5016 [14]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6192 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11944  (
    .i0(\u2_Display/n6158 ),
    .i1(\u2_Display/n5016 [13]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6193 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11945  (
    .i0(\u2_Display/n6159 ),
    .i1(\u2_Display/n5016 [12]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6194 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11946  (
    .i0(\u2_Display/n6160 ),
    .i1(\u2_Display/n5016 [11]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6195 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11947  (
    .i0(\u2_Display/n6161 ),
    .i1(\u2_Display/n5016 [10]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6196 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11948  (
    .i0(\u2_Display/n6162 ),
    .i1(\u2_Display/n5016 [9]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6197 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11949  (
    .i0(\u2_Display/n6163 ),
    .i1(\u2_Display/n5016 [8]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6198 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11950  (
    .i0(\u2_Display/n6164 ),
    .i1(\u2_Display/n5016 [7]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6199 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11951  (
    .i0(\u2_Display/n6165 ),
    .i1(\u2_Display/n5016 [6]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6200 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11952  (
    .i0(\u2_Display/n6166 ),
    .i1(\u2_Display/n5016 [5]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6201 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11953  (
    .i0(\u2_Display/n6167 ),
    .i1(\u2_Display/n5016 [4]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6202 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11954  (
    .i0(\u2_Display/n6168 ),
    .i1(\u2_Display/n5016 [3]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6203 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11955  (
    .i0(\u2_Display/n6169 ),
    .i1(\u2_Display/n5016 [2]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6204 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11956  (
    .i0(\u2_Display/n6170 ),
    .i1(\u2_Display/n5016 [1]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6205 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11957  (
    .i0(\u2_Display/n6171 ),
    .i1(\u2_Display/n5016 [0]),
    .sel(\u2_Display/n6173 ),
    .o(\u2_Display/n6206 ));  // source/rtl/Display.v(163)
  not \u2_Display/u11958  (\u2_Display/n6208 , \u2_Display/n5049 );  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11991  (
    .i0(\u2_Display/n6175 ),
    .i1(\u2_Display/n5051 [31]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6210 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11992  (
    .i0(\u2_Display/n6176 ),
    .i1(\u2_Display/n5051 [30]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6211 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11993  (
    .i0(\u2_Display/n6177 ),
    .i1(\u2_Display/n5051 [29]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6212 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11994  (
    .i0(\u2_Display/n6178 ),
    .i1(\u2_Display/n5051 [28]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6213 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11995  (
    .i0(\u2_Display/n6179 ),
    .i1(\u2_Display/n5051 [27]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6214 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11996  (
    .i0(\u2_Display/n6180 ),
    .i1(\u2_Display/n5051 [26]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6215 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11997  (
    .i0(\u2_Display/n6181 ),
    .i1(\u2_Display/n5051 [25]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6216 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11998  (
    .i0(\u2_Display/n6182 ),
    .i1(\u2_Display/n5051 [24]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6217 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u11999  (
    .i0(\u2_Display/n6183 ),
    .i1(\u2_Display/n5051 [23]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6218 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12000  (
    .i0(\u2_Display/n6184 ),
    .i1(\u2_Display/n5051 [22]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6219 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12001  (
    .i0(\u2_Display/n6185 ),
    .i1(\u2_Display/n5051 [21]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6220 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12002  (
    .i0(\u2_Display/n6186 ),
    .i1(\u2_Display/n5051 [20]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6221 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12003  (
    .i0(\u2_Display/n6187 ),
    .i1(\u2_Display/n5051 [19]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6222 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12004  (
    .i0(\u2_Display/n6188 ),
    .i1(\u2_Display/n5051 [18]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6223 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12005  (
    .i0(\u2_Display/n6189 ),
    .i1(\u2_Display/n5051 [17]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6224 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12006  (
    .i0(\u2_Display/n6190 ),
    .i1(\u2_Display/n5051 [16]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6225 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12007  (
    .i0(\u2_Display/n6191 ),
    .i1(\u2_Display/n5051 [15]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6226 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12008  (
    .i0(\u2_Display/n6192 ),
    .i1(\u2_Display/n5051 [14]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6227 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12009  (
    .i0(\u2_Display/n6193 ),
    .i1(\u2_Display/n5051 [13]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6228 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12010  (
    .i0(\u2_Display/n6194 ),
    .i1(\u2_Display/n5051 [12]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6229 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12011  (
    .i0(\u2_Display/n6195 ),
    .i1(\u2_Display/n5051 [11]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6230 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12012  (
    .i0(\u2_Display/n6196 ),
    .i1(\u2_Display/n5051 [10]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6231 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12013  (
    .i0(\u2_Display/n6197 ),
    .i1(\u2_Display/n5051 [9]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6232 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12014  (
    .i0(\u2_Display/n6198 ),
    .i1(\u2_Display/n5051 [8]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6233 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12015  (
    .i0(\u2_Display/n6199 ),
    .i1(\u2_Display/n5051 [7]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6234 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12016  (
    .i0(\u2_Display/n6200 ),
    .i1(\u2_Display/n5051 [6]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6235 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12017  (
    .i0(\u2_Display/n6201 ),
    .i1(\u2_Display/n5051 [5]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6236 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12018  (
    .i0(\u2_Display/n6202 ),
    .i1(\u2_Display/n5051 [4]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6237 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12019  (
    .i0(\u2_Display/n6203 ),
    .i1(\u2_Display/n5051 [3]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6238 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12020  (
    .i0(\u2_Display/n6204 ),
    .i1(\u2_Display/n5051 [2]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6239 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12021  (
    .i0(\u2_Display/n6205 ),
    .i1(\u2_Display/n5051 [1]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6240 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12022  (
    .i0(\u2_Display/n6206 ),
    .i1(\u2_Display/n5051 [0]),
    .sel(\u2_Display/n6208 ),
    .o(\u2_Display/n6241 ));  // source/rtl/Display.v(163)
  not \u2_Display/u12023  (\u2_Display/n6243 , \u2_Display/n5084 );  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12056  (
    .i0(\u2_Display/n6210 ),
    .i1(\u2_Display/n5086 [31]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6245 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12057  (
    .i0(\u2_Display/n6211 ),
    .i1(\u2_Display/n5086 [30]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6246 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12058  (
    .i0(\u2_Display/n6212 ),
    .i1(\u2_Display/n5086 [29]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6247 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12059  (
    .i0(\u2_Display/n6213 ),
    .i1(\u2_Display/n5086 [28]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6248 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12060  (
    .i0(\u2_Display/n6214 ),
    .i1(\u2_Display/n5086 [27]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6249 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12061  (
    .i0(\u2_Display/n6215 ),
    .i1(\u2_Display/n5086 [26]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6250 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12062  (
    .i0(\u2_Display/n6216 ),
    .i1(\u2_Display/n5086 [25]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6251 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12063  (
    .i0(\u2_Display/n6217 ),
    .i1(\u2_Display/n5086 [24]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6252 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12064  (
    .i0(\u2_Display/n6218 ),
    .i1(\u2_Display/n5086 [23]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6253 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12065  (
    .i0(\u2_Display/n6219 ),
    .i1(\u2_Display/n5086 [22]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6254 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12066  (
    .i0(\u2_Display/n6220 ),
    .i1(\u2_Display/n5086 [21]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6255 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12067  (
    .i0(\u2_Display/n6221 ),
    .i1(\u2_Display/n5086 [20]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6256 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12068  (
    .i0(\u2_Display/n6222 ),
    .i1(\u2_Display/n5086 [19]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6257 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12069  (
    .i0(\u2_Display/n6223 ),
    .i1(\u2_Display/n5086 [18]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6258 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12070  (
    .i0(\u2_Display/n6224 ),
    .i1(\u2_Display/n5086 [17]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6259 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12071  (
    .i0(\u2_Display/n6225 ),
    .i1(\u2_Display/n5086 [16]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6260 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12072  (
    .i0(\u2_Display/n6226 ),
    .i1(\u2_Display/n5086 [15]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6261 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12073  (
    .i0(\u2_Display/n6227 ),
    .i1(\u2_Display/n5086 [14]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6262 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12074  (
    .i0(\u2_Display/n6228 ),
    .i1(\u2_Display/n5086 [13]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6263 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12075  (
    .i0(\u2_Display/n6229 ),
    .i1(\u2_Display/n5086 [12]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6264 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12076  (
    .i0(\u2_Display/n6230 ),
    .i1(\u2_Display/n5086 [11]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6265 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12077  (
    .i0(\u2_Display/n6231 ),
    .i1(\u2_Display/n5086 [10]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6266 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12078  (
    .i0(\u2_Display/n6232 ),
    .i1(\u2_Display/n5086 [9]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6267 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12079  (
    .i0(\u2_Display/n6233 ),
    .i1(\u2_Display/n5086 [8]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6268 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12080  (
    .i0(\u2_Display/n6234 ),
    .i1(\u2_Display/n5086 [7]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6269 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12081  (
    .i0(\u2_Display/n6235 ),
    .i1(\u2_Display/n5086 [6]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6270 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12082  (
    .i0(\u2_Display/n6236 ),
    .i1(\u2_Display/n5086 [5]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6271 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12083  (
    .i0(\u2_Display/n6237 ),
    .i1(\u2_Display/n5086 [4]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6272 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12084  (
    .i0(\u2_Display/n6238 ),
    .i1(\u2_Display/n5086 [3]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6273 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12085  (
    .i0(\u2_Display/n6239 ),
    .i1(\u2_Display/n5086 [2]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6274 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12086  (
    .i0(\u2_Display/n6240 ),
    .i1(\u2_Display/n5086 [1]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6275 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12087  (
    .i0(\u2_Display/n6241 ),
    .i1(\u2_Display/n5086 [0]),
    .sel(\u2_Display/n6243 ),
    .o(\u2_Display/n6276 ));  // source/rtl/Display.v(163)
  not \u2_Display/u12088  (\u2_Display/n6278 , \u2_Display/n5119 );  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12121  (
    .i0(\u2_Display/n6245 ),
    .i1(\u2_Display/n5121 [31]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6280 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12122  (
    .i0(\u2_Display/n6246 ),
    .i1(\u2_Display/n5121 [30]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6281 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12123  (
    .i0(\u2_Display/n6247 ),
    .i1(\u2_Display/n5121 [29]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6282 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12124  (
    .i0(\u2_Display/n6248 ),
    .i1(\u2_Display/n5121 [28]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6283 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12125  (
    .i0(\u2_Display/n6249 ),
    .i1(\u2_Display/n5121 [27]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6284 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12126  (
    .i0(\u2_Display/n6250 ),
    .i1(\u2_Display/n5121 [26]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6285 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12127  (
    .i0(\u2_Display/n6251 ),
    .i1(\u2_Display/n5121 [25]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6286 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12128  (
    .i0(\u2_Display/n6252 ),
    .i1(\u2_Display/n5121 [24]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6287 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12129  (
    .i0(\u2_Display/n6253 ),
    .i1(\u2_Display/n5121 [23]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6288 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12130  (
    .i0(\u2_Display/n6254 ),
    .i1(\u2_Display/n5121 [22]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6289 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12131  (
    .i0(\u2_Display/n6255 ),
    .i1(\u2_Display/n5121 [21]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6290 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12132  (
    .i0(\u2_Display/n6256 ),
    .i1(\u2_Display/n5121 [20]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6291 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12133  (
    .i0(\u2_Display/n6257 ),
    .i1(\u2_Display/n5121 [19]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6292 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12134  (
    .i0(\u2_Display/n6258 ),
    .i1(\u2_Display/n5121 [18]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6293 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12135  (
    .i0(\u2_Display/n6259 ),
    .i1(\u2_Display/n5121 [17]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6294 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12136  (
    .i0(\u2_Display/n6260 ),
    .i1(\u2_Display/n5121 [16]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6295 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12137  (
    .i0(\u2_Display/n6261 ),
    .i1(\u2_Display/n5121 [15]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6296 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12138  (
    .i0(\u2_Display/n6262 ),
    .i1(\u2_Display/n5121 [14]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6297 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12139  (
    .i0(\u2_Display/n6263 ),
    .i1(\u2_Display/n5121 [13]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6298 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12140  (
    .i0(\u2_Display/n6264 ),
    .i1(\u2_Display/n5121 [12]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6299 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12141  (
    .i0(\u2_Display/n6265 ),
    .i1(\u2_Display/n5121 [11]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6300 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12142  (
    .i0(\u2_Display/n6266 ),
    .i1(\u2_Display/n5121 [10]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6301 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12143  (
    .i0(\u2_Display/n6267 ),
    .i1(\u2_Display/n5121 [9]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6302 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12144  (
    .i0(\u2_Display/n6268 ),
    .i1(\u2_Display/n5121 [8]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6303 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12145  (
    .i0(\u2_Display/n6269 ),
    .i1(\u2_Display/n5121 [7]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6304 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12146  (
    .i0(\u2_Display/n6270 ),
    .i1(\u2_Display/n5121 [6]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6305 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12147  (
    .i0(\u2_Display/n6271 ),
    .i1(\u2_Display/n5121 [5]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6306 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12148  (
    .i0(\u2_Display/n6272 ),
    .i1(\u2_Display/n5121 [4]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6307 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12149  (
    .i0(\u2_Display/n6273 ),
    .i1(\u2_Display/n5121 [3]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6308 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1215  (
    .i0(\u2_Display/n630 ),
    .i1(\u2_Display/n664 [31]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n665 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u12150  (
    .i0(\u2_Display/n6274 ),
    .i1(\u2_Display/n5121 [2]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6309 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12151  (
    .i0(\u2_Display/n6275 ),
    .i1(\u2_Display/n5121 [1]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6310 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12152  (
    .i0(\u2_Display/n6276 ),
    .i1(\u2_Display/n5121 [0]),
    .sel(\u2_Display/n6278 ),
    .o(\u2_Display/n6311 ));  // source/rtl/Display.v(163)
  not \u2_Display/u12153  (\u2_Display/n6313 , \u2_Display/n5154 );  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1216  (
    .i0(\u2_Display/n631 ),
    .i1(\u2_Display/n664 [30]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n666 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1217  (
    .i0(\u2_Display/n632 ),
    .i1(\u2_Display/n664 [29]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n667 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1218  (
    .i0(\u2_Display/n633 ),
    .i1(\u2_Display/n664 [28]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n668 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u12186  (
    .i0(\u2_Display/n6280 ),
    .i1(\u2_Display/n5156 [31]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6315 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12187  (
    .i0(\u2_Display/n6281 ),
    .i1(\u2_Display/n5156 [30]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6316 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12188  (
    .i0(\u2_Display/n6282 ),
    .i1(\u2_Display/n5156 [29]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6317 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12189  (
    .i0(\u2_Display/n6283 ),
    .i1(\u2_Display/n5156 [28]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6318 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1219  (
    .i0(\u2_Display/n634 ),
    .i1(\u2_Display/n664 [27]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n669 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u12190  (
    .i0(\u2_Display/n6284 ),
    .i1(\u2_Display/n5156 [27]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6319 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12191  (
    .i0(\u2_Display/n6285 ),
    .i1(\u2_Display/n5156 [26]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6320 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12192  (
    .i0(\u2_Display/n6286 ),
    .i1(\u2_Display/n5156 [25]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6321 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12193  (
    .i0(\u2_Display/n6287 ),
    .i1(\u2_Display/n5156 [24]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6322 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12194  (
    .i0(\u2_Display/n6288 ),
    .i1(\u2_Display/n5156 [23]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6323 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12195  (
    .i0(\u2_Display/n6289 ),
    .i1(\u2_Display/n5156 [22]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6324 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12196  (
    .i0(\u2_Display/n6290 ),
    .i1(\u2_Display/n5156 [21]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6325 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12197  (
    .i0(\u2_Display/n6291 ),
    .i1(\u2_Display/n5156 [20]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6326 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12198  (
    .i0(\u2_Display/n6292 ),
    .i1(\u2_Display/n5156 [19]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6327 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12199  (
    .i0(\u2_Display/n6293 ),
    .i1(\u2_Display/n5156 [18]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6328 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1220  (
    .i0(\u2_Display/n635 ),
    .i1(\u2_Display/n664 [26]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n670 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u12200  (
    .i0(\u2_Display/n6294 ),
    .i1(\u2_Display/n5156 [17]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6329 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12201  (
    .i0(\u2_Display/n6295 ),
    .i1(\u2_Display/n5156 [16]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6330 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12202  (
    .i0(\u2_Display/n6296 ),
    .i1(\u2_Display/n5156 [15]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6331 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12203  (
    .i0(\u2_Display/n6297 ),
    .i1(\u2_Display/n5156 [14]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6332 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12204  (
    .i0(\u2_Display/n6298 ),
    .i1(\u2_Display/n5156 [13]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6333 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12205  (
    .i0(\u2_Display/n6299 ),
    .i1(\u2_Display/n5156 [12]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6334 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12206  (
    .i0(\u2_Display/n6300 ),
    .i1(\u2_Display/n5156 [11]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6335 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12207  (
    .i0(\u2_Display/n6301 ),
    .i1(\u2_Display/n5156 [10]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6336 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12208  (
    .i0(\u2_Display/n6302 ),
    .i1(\u2_Display/n5156 [9]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6337 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12209  (
    .i0(\u2_Display/n6303 ),
    .i1(\u2_Display/n5156 [8]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6338 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1221  (
    .i0(\u2_Display/n636 ),
    .i1(\u2_Display/n664 [25]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n671 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u12210  (
    .i0(\u2_Display/n6304 ),
    .i1(\u2_Display/n5156 [7]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6339 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12211  (
    .i0(\u2_Display/n6305 ),
    .i1(\u2_Display/n5156 [6]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6340 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12212  (
    .i0(\u2_Display/n6306 ),
    .i1(\u2_Display/n5156 [5]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6341 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12213  (
    .i0(\u2_Display/n6307 ),
    .i1(\u2_Display/n5156 [4]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6342 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12214  (
    .i0(\u2_Display/n6308 ),
    .i1(\u2_Display/n5156 [3]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6343 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12215  (
    .i0(\u2_Display/n6309 ),
    .i1(\u2_Display/n5156 [2]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6344 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12216  (
    .i0(\u2_Display/n6310 ),
    .i1(\u2_Display/n5156 [1]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6345 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12217  (
    .i0(\u2_Display/n6311 ),
    .i1(\u2_Display/n5156 [0]),
    .sel(\u2_Display/n6313 ),
    .o(\u2_Display/n6346 ));  // source/rtl/Display.v(163)
  not \u2_Display/u12218  (\u2_Display/n6348 , \u2_Display/n5189 );  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1222  (
    .i0(\u2_Display/n637 ),
    .i1(\u2_Display/n664 [24]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n672 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1223  (
    .i0(\u2_Display/n638 ),
    .i1(\u2_Display/n664 [23]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n673 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1224  (
    .i0(\u2_Display/n639 ),
    .i1(\u2_Display/n664 [22]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n674 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1225  (
    .i0(\u2_Display/n640 ),
    .i1(\u2_Display/n664 [21]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n675 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u12251  (
    .i0(\u2_Display/n6315 ),
    .i1(\u2_Display/n5191 [31]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n6350 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12252  (
    .i0(\u2_Display/n6316 ),
    .i1(\u2_Display/n5191 [30]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n6351 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12253  (
    .i0(\u2_Display/n6317 ),
    .i1(\u2_Display/n5191 [29]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n6352 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u12254  (
    .i0(\u2_Display/n6318 ),
    .i1(\u2_Display/n5191 [28]),
    .sel(\u2_Display/n6348 ),
    .o(\u2_Display/n6353 ));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1226  (
    .i0(\u2_Display/n641 ),
    .i1(\u2_Display/n664 [20]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n676 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1227  (
    .i0(\u2_Display/n642 ),
    .i1(\u2_Display/n664 [19]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n677 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1228  (
    .i0(\u2_Display/n643 ),
    .i1(\u2_Display/n664 [18]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n678 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1229  (
    .i0(\u2_Display/n644 ),
    .i1(\u2_Display/n664 [17]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n679 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1230  (
    .i0(\u2_Display/n645 ),
    .i1(\u2_Display/n664 [16]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n680 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1231  (
    .i0(\u2_Display/n646 ),
    .i1(\u2_Display/n664 [15]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n681 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1232  (
    .i0(\u2_Display/n647 ),
    .i1(\u2_Display/n664 [14]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n682 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1233  (
    .i0(\u2_Display/n648 ),
    .i1(\u2_Display/n664 [13]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n683 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1234  (
    .i0(\u2_Display/n649 ),
    .i1(\u2_Display/n664 [12]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n684 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1235  (
    .i0(\u2_Display/n650 ),
    .i1(\u2_Display/n664 [11]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n685 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1236  (
    .i0(\u2_Display/n651 ),
    .i1(\u2_Display/n664 [10]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n686 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1237  (
    .i0(\u2_Display/n652 ),
    .i1(\u2_Display/n664 [9]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n687 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1238  (
    .i0(\u2_Display/n653 ),
    .i1(\u2_Display/n664 [8]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n688 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1239  (
    .i0(\u2_Display/n654 ),
    .i1(\u2_Display/n664 [7]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n689 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1240  (
    .i0(\u2_Display/n655 ),
    .i1(\u2_Display/n664 [6]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n690 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1241  (
    .i0(\u2_Display/n656 ),
    .i1(\u2_Display/n664 [5]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n691 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1242  (
    .i0(\u2_Display/n657 ),
    .i1(\u2_Display/n664 [4]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n692 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1243  (
    .i0(\u2_Display/n658 ),
    .i1(\u2_Display/n664 [3]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n693 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1244  (
    .i0(\u2_Display/n659 ),
    .i1(\u2_Display/n664 [2]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n694 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1245  (
    .i0(\u2_Display/n660 ),
    .i1(\u2_Display/n664 [1]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n695 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1246  (
    .i0(\u2_Display/n661 ),
    .i1(\u2_Display/n664 [0]),
    .sel(\u2_Display/n663 ),
    .o(\u2_Display/n696 ));  // source/rtl/Display.v(230)
  not \u2_Display/u1247  (\u2_Display/n698 , \u2_Display/n697 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1280  (
    .i0(\u2_Display/n665 ),
    .i1(\u2_Display/n699 [31]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n700 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1281  (
    .i0(\u2_Display/n666 ),
    .i1(\u2_Display/n699 [30]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n701 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1282  (
    .i0(\u2_Display/n667 ),
    .i1(\u2_Display/n699 [29]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n702 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1283  (
    .i0(\u2_Display/n668 ),
    .i1(\u2_Display/n699 [28]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n703 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1284  (
    .i0(\u2_Display/n669 ),
    .i1(\u2_Display/n699 [27]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n704 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1285  (
    .i0(\u2_Display/n670 ),
    .i1(\u2_Display/n699 [26]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n705 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1286  (
    .i0(\u2_Display/n671 ),
    .i1(\u2_Display/n699 [25]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n706 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1287  (
    .i0(\u2_Display/n672 ),
    .i1(\u2_Display/n699 [24]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n707 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1288  (
    .i0(\u2_Display/n673 ),
    .i1(\u2_Display/n699 [23]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n708 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1289  (
    .i0(\u2_Display/n674 ),
    .i1(\u2_Display/n699 [22]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n709 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1290  (
    .i0(\u2_Display/n675 ),
    .i1(\u2_Display/n699 [21]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n710 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1291  (
    .i0(\u2_Display/n676 ),
    .i1(\u2_Display/n699 [20]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n711 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1292  (
    .i0(\u2_Display/n677 ),
    .i1(\u2_Display/n699 [19]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n712 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1293  (
    .i0(\u2_Display/n678 ),
    .i1(\u2_Display/n699 [18]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n713 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1294  (
    .i0(\u2_Display/n679 ),
    .i1(\u2_Display/n699 [17]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n714 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1295  (
    .i0(\u2_Display/n680 ),
    .i1(\u2_Display/n699 [16]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n715 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1296  (
    .i0(\u2_Display/n681 ),
    .i1(\u2_Display/n699 [15]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n716 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1297  (
    .i0(\u2_Display/n682 ),
    .i1(\u2_Display/n699 [14]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n717 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1298  (
    .i0(\u2_Display/n683 ),
    .i1(\u2_Display/n699 [13]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n718 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1299  (
    .i0(\u2_Display/n684 ),
    .i1(\u2_Display/n699 [12]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n719 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1300  (
    .i0(\u2_Display/n685 ),
    .i1(\u2_Display/n699 [11]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n720 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1301  (
    .i0(\u2_Display/n686 ),
    .i1(\u2_Display/n699 [10]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n721 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1302  (
    .i0(\u2_Display/n687 ),
    .i1(\u2_Display/n699 [9]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n722 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1303  (
    .i0(\u2_Display/n688 ),
    .i1(\u2_Display/n699 [8]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n723 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1304  (
    .i0(\u2_Display/n689 ),
    .i1(\u2_Display/n699 [7]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n724 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1305  (
    .i0(\u2_Display/n690 ),
    .i1(\u2_Display/n699 [6]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n725 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1306  (
    .i0(\u2_Display/n691 ),
    .i1(\u2_Display/n699 [5]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n726 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1307  (
    .i0(\u2_Display/n692 ),
    .i1(\u2_Display/n699 [4]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n727 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1308  (
    .i0(\u2_Display/n693 ),
    .i1(\u2_Display/n699 [3]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n728 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1309  (
    .i0(\u2_Display/n694 ),
    .i1(\u2_Display/n699 [2]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n729 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u13095  (
    .i0(\u2_Display/n5633 ),
    .i1(\u2_Display/n6804 [10]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n42 [10]));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u13096  (
    .i0(\u2_Display/n5634 ),
    .i1(\u2_Display/n6804 [9]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n42 [9]));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u13097  (
    .i0(\u2_Display/n5635 ),
    .i1(\u2_Display/n6804 [8]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n42 [8]));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u13098  (
    .i0(\u2_Display/n5636 ),
    .i1(\u2_Display/n6804 [7]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n42 [7]));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u13099  (
    .i0(\u2_Display/n5637 ),
    .i1(\u2_Display/n6804 [6]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n42 [6]));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1310  (
    .i0(\u2_Display/n695 ),
    .i1(\u2_Display/n699 [1]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n730 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u13100  (
    .i0(\u2_Display/n5638 ),
    .i1(\u2_Display/n6804 [5]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n42 [5]));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u13101  (
    .i0(\u2_Display/n5639 ),
    .i1(\u2_Display/n6804 [4]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n42 [4]));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u13102  (
    .i0(\u2_Display/n5640 ),
    .i1(\u2_Display/n6804 [3]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n42 [3]));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u13103  (
    .i0(\u2_Display/n5641 ),
    .i1(\u2_Display/n6804 [2]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n42 [2]));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u13104  (
    .i0(\u2_Display/n5642 ),
    .i1(\u2_Display/n6804 [1]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n42 [1]));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u13105  (
    .i0(\u2_Display/n5643 ),
    .i1(\u2_Display/n6804 [0]),
    .sel(\u2_Display/n5645 ),
    .o(\u2_Display/n42 [0]));  // source/rtl/Display.v(163)
  AL_MUX \u2_Display/u1311  (
    .i0(\u2_Display/n696 ),
    .i1(\u2_Display/n699 [0]),
    .sel(\u2_Display/n698 ),
    .o(\u2_Display/n731 ));  // source/rtl/Display.v(230)
  not \u2_Display/u1312  (\u2_Display/n733 , \u2_Display/n732 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1345  (
    .i0(\u2_Display/n700 ),
    .i1(\u2_Display/n734 [31]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n735 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1346  (
    .i0(\u2_Display/n701 ),
    .i1(\u2_Display/n734 [30]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n736 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1347  (
    .i0(\u2_Display/n702 ),
    .i1(\u2_Display/n734 [29]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n737 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1348  (
    .i0(\u2_Display/n703 ),
    .i1(\u2_Display/n734 [28]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n738 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1349  (
    .i0(\u2_Display/n704 ),
    .i1(\u2_Display/n734 [27]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n739 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1350  (
    .i0(\u2_Display/n705 ),
    .i1(\u2_Display/n734 [26]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n740 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1351  (
    .i0(\u2_Display/n706 ),
    .i1(\u2_Display/n734 [25]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n741 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1352  (
    .i0(\u2_Display/n707 ),
    .i1(\u2_Display/n734 [24]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n742 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1353  (
    .i0(\u2_Display/n708 ),
    .i1(\u2_Display/n734 [23]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n743 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1354  (
    .i0(\u2_Display/n709 ),
    .i1(\u2_Display/n734 [22]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n744 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1355  (
    .i0(\u2_Display/n710 ),
    .i1(\u2_Display/n734 [21]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n745 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1356  (
    .i0(\u2_Display/n711 ),
    .i1(\u2_Display/n734 [20]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n746 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1357  (
    .i0(\u2_Display/n712 ),
    .i1(\u2_Display/n734 [19]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n747 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1358  (
    .i0(\u2_Display/n713 ),
    .i1(\u2_Display/n734 [18]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n748 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1359  (
    .i0(\u2_Display/n714 ),
    .i1(\u2_Display/n734 [17]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n749 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1360  (
    .i0(\u2_Display/n715 ),
    .i1(\u2_Display/n734 [16]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n750 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1361  (
    .i0(\u2_Display/n716 ),
    .i1(\u2_Display/n734 [15]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n751 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1362  (
    .i0(\u2_Display/n717 ),
    .i1(\u2_Display/n734 [14]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n752 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1363  (
    .i0(\u2_Display/n718 ),
    .i1(\u2_Display/n734 [13]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n753 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1364  (
    .i0(\u2_Display/n719 ),
    .i1(\u2_Display/n734 [12]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n754 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1365  (
    .i0(\u2_Display/n720 ),
    .i1(\u2_Display/n734 [11]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n755 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1366  (
    .i0(\u2_Display/n721 ),
    .i1(\u2_Display/n734 [10]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n756 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1367  (
    .i0(\u2_Display/n722 ),
    .i1(\u2_Display/n734 [9]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n757 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1368  (
    .i0(\u2_Display/n723 ),
    .i1(\u2_Display/n734 [8]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n758 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1369  (
    .i0(\u2_Display/n724 ),
    .i1(\u2_Display/n734 [7]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n759 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1370  (
    .i0(\u2_Display/n725 ),
    .i1(\u2_Display/n734 [6]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n760 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1371  (
    .i0(\u2_Display/n726 ),
    .i1(\u2_Display/n734 [5]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n761 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1372  (
    .i0(\u2_Display/n727 ),
    .i1(\u2_Display/n734 [4]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n762 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1373  (
    .i0(\u2_Display/n728 ),
    .i1(\u2_Display/n734 [3]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n763 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1374  (
    .i0(\u2_Display/n729 ),
    .i1(\u2_Display/n734 [2]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n764 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1375  (
    .i0(\u2_Display/n730 ),
    .i1(\u2_Display/n734 [1]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n765 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1376  (
    .i0(\u2_Display/n731 ),
    .i1(\u2_Display/n734 [0]),
    .sel(\u2_Display/n733 ),
    .o(\u2_Display/n766 ));  // source/rtl/Display.v(230)
  not \u2_Display/u1377  (\u2_Display/n768 , \u2_Display/n767 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1410  (
    .i0(\u2_Display/n735 ),
    .i1(\u2_Display/n769 [31]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n770 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1411  (
    .i0(\u2_Display/n736 ),
    .i1(\u2_Display/n769 [30]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n771 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1412  (
    .i0(\u2_Display/n737 ),
    .i1(\u2_Display/n769 [29]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n772 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1413  (
    .i0(\u2_Display/n738 ),
    .i1(\u2_Display/n769 [28]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n773 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1414  (
    .i0(\u2_Display/n739 ),
    .i1(\u2_Display/n769 [27]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n774 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1415  (
    .i0(\u2_Display/n740 ),
    .i1(\u2_Display/n769 [26]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n775 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1416  (
    .i0(\u2_Display/n741 ),
    .i1(\u2_Display/n769 [25]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n776 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1417  (
    .i0(\u2_Display/n742 ),
    .i1(\u2_Display/n769 [24]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n777 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1418  (
    .i0(\u2_Display/n743 ),
    .i1(\u2_Display/n769 [23]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n778 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1419  (
    .i0(\u2_Display/n744 ),
    .i1(\u2_Display/n769 [22]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n779 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1420  (
    .i0(\u2_Display/n745 ),
    .i1(\u2_Display/n769 [21]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n780 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1421  (
    .i0(\u2_Display/n746 ),
    .i1(\u2_Display/n769 [20]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n781 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1422  (
    .i0(\u2_Display/n747 ),
    .i1(\u2_Display/n769 [19]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n782 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1423  (
    .i0(\u2_Display/n748 ),
    .i1(\u2_Display/n769 [18]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n783 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1424  (
    .i0(\u2_Display/n749 ),
    .i1(\u2_Display/n769 [17]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n784 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1425  (
    .i0(\u2_Display/n750 ),
    .i1(\u2_Display/n769 [16]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n785 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1426  (
    .i0(\u2_Display/n751 ),
    .i1(\u2_Display/n769 [15]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n786 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1427  (
    .i0(\u2_Display/n752 ),
    .i1(\u2_Display/n769 [14]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n787 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1428  (
    .i0(\u2_Display/n753 ),
    .i1(\u2_Display/n769 [13]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n788 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1429  (
    .i0(\u2_Display/n754 ),
    .i1(\u2_Display/n769 [12]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n789 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1430  (
    .i0(\u2_Display/n755 ),
    .i1(\u2_Display/n769 [11]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n790 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1431  (
    .i0(\u2_Display/n756 ),
    .i1(\u2_Display/n769 [10]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n791 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1432  (
    .i0(\u2_Display/n757 ),
    .i1(\u2_Display/n769 [9]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n792 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1433  (
    .i0(\u2_Display/n758 ),
    .i1(\u2_Display/n769 [8]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n793 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1434  (
    .i0(\u2_Display/n759 ),
    .i1(\u2_Display/n769 [7]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n794 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1435  (
    .i0(\u2_Display/n760 ),
    .i1(\u2_Display/n769 [6]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n795 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1436  (
    .i0(\u2_Display/n761 ),
    .i1(\u2_Display/n769 [5]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n796 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1437  (
    .i0(\u2_Display/n762 ),
    .i1(\u2_Display/n769 [4]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n797 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1438  (
    .i0(\u2_Display/n763 ),
    .i1(\u2_Display/n769 [3]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n798 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1439  (
    .i0(\u2_Display/n764 ),
    .i1(\u2_Display/n769 [2]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n799 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1440  (
    .i0(\u2_Display/n765 ),
    .i1(\u2_Display/n769 [1]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n800 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1441  (
    .i0(\u2_Display/n766 ),
    .i1(\u2_Display/n769 [0]),
    .sel(\u2_Display/n768 ),
    .o(\u2_Display/n801 ));  // source/rtl/Display.v(230)
  not \u2_Display/u1442  (\u2_Display/n803 , \u2_Display/n802 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1475  (
    .i0(\u2_Display/n770 ),
    .i1(\u2_Display/n804 [31]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n805 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1476  (
    .i0(\u2_Display/n771 ),
    .i1(\u2_Display/n804 [30]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n806 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1477  (
    .i0(\u2_Display/n772 ),
    .i1(\u2_Display/n804 [29]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n807 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1478  (
    .i0(\u2_Display/n773 ),
    .i1(\u2_Display/n804 [28]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n808 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1479  (
    .i0(\u2_Display/n774 ),
    .i1(\u2_Display/n804 [27]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n809 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1480  (
    .i0(\u2_Display/n775 ),
    .i1(\u2_Display/n804 [26]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n810 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1481  (
    .i0(\u2_Display/n776 ),
    .i1(\u2_Display/n804 [25]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n811 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1482  (
    .i0(\u2_Display/n777 ),
    .i1(\u2_Display/n804 [24]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n812 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1483  (
    .i0(\u2_Display/n778 ),
    .i1(\u2_Display/n804 [23]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n813 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1484  (
    .i0(\u2_Display/n779 ),
    .i1(\u2_Display/n804 [22]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n814 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1485  (
    .i0(\u2_Display/n780 ),
    .i1(\u2_Display/n804 [21]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n815 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1486  (
    .i0(\u2_Display/n781 ),
    .i1(\u2_Display/n804 [20]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n816 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1487  (
    .i0(\u2_Display/n782 ),
    .i1(\u2_Display/n804 [19]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n817 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1488  (
    .i0(\u2_Display/n783 ),
    .i1(\u2_Display/n804 [18]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n818 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1489  (
    .i0(\u2_Display/n784 ),
    .i1(\u2_Display/n804 [17]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n819 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1490  (
    .i0(\u2_Display/n785 ),
    .i1(\u2_Display/n804 [16]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n820 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1491  (
    .i0(\u2_Display/n786 ),
    .i1(\u2_Display/n804 [15]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n821 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1492  (
    .i0(\u2_Display/n787 ),
    .i1(\u2_Display/n804 [14]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n822 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1493  (
    .i0(\u2_Display/n788 ),
    .i1(\u2_Display/n804 [13]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n823 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1494  (
    .i0(\u2_Display/n789 ),
    .i1(\u2_Display/n804 [12]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n824 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1495  (
    .i0(\u2_Display/n790 ),
    .i1(\u2_Display/n804 [11]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n825 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1496  (
    .i0(\u2_Display/n791 ),
    .i1(\u2_Display/n804 [10]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n826 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1497  (
    .i0(\u2_Display/n792 ),
    .i1(\u2_Display/n804 [9]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n827 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1498  (
    .i0(\u2_Display/n793 ),
    .i1(\u2_Display/n804 [8]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n828 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1499  (
    .i0(\u2_Display/n794 ),
    .i1(\u2_Display/n804 [7]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n829 ));  // source/rtl/Display.v(230)
  and \u2_Display/u15  (\u2_Display/n98 , \u2_Display/n95 , \u2_Display/n97 );  // source/rtl/Display.v(181)
  AL_MUX \u2_Display/u1500  (
    .i0(\u2_Display/n795 ),
    .i1(\u2_Display/n804 [6]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n830 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1501  (
    .i0(\u2_Display/n796 ),
    .i1(\u2_Display/n804 [5]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n831 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1502  (
    .i0(\u2_Display/n797 ),
    .i1(\u2_Display/n804 [4]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n832 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1503  (
    .i0(\u2_Display/n798 ),
    .i1(\u2_Display/n804 [3]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n833 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1504  (
    .i0(\u2_Display/n799 ),
    .i1(\u2_Display/n804 [2]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n834 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1505  (
    .i0(\u2_Display/n800 ),
    .i1(\u2_Display/n804 [1]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n835 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1506  (
    .i0(\u2_Display/n801 ),
    .i1(\u2_Display/n804 [0]),
    .sel(\u2_Display/n803 ),
    .o(\u2_Display/n836 ));  // source/rtl/Display.v(230)
  not \u2_Display/u1507  (\u2_Display/n838 , \u2_Display/n837 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1540  (
    .i0(\u2_Display/n805 ),
    .i1(\u2_Display/n839 [31]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n840 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1541  (
    .i0(\u2_Display/n806 ),
    .i1(\u2_Display/n839 [30]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n841 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1542  (
    .i0(\u2_Display/n807 ),
    .i1(\u2_Display/n839 [29]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n842 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1543  (
    .i0(\u2_Display/n808 ),
    .i1(\u2_Display/n839 [28]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n843 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1544  (
    .i0(\u2_Display/n809 ),
    .i1(\u2_Display/n839 [27]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n844 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1545  (
    .i0(\u2_Display/n810 ),
    .i1(\u2_Display/n839 [26]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n845 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1546  (
    .i0(\u2_Display/n811 ),
    .i1(\u2_Display/n839 [25]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n846 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1547  (
    .i0(\u2_Display/n812 ),
    .i1(\u2_Display/n839 [24]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n847 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1548  (
    .i0(\u2_Display/n813 ),
    .i1(\u2_Display/n839 [23]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n848 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1549  (
    .i0(\u2_Display/n814 ),
    .i1(\u2_Display/n839 [22]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n849 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1550  (
    .i0(\u2_Display/n815 ),
    .i1(\u2_Display/n839 [21]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n850 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1551  (
    .i0(\u2_Display/n816 ),
    .i1(\u2_Display/n839 [20]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n851 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1552  (
    .i0(\u2_Display/n817 ),
    .i1(\u2_Display/n839 [19]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n852 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1553  (
    .i0(\u2_Display/n818 ),
    .i1(\u2_Display/n839 [18]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n853 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1554  (
    .i0(\u2_Display/n819 ),
    .i1(\u2_Display/n839 [17]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n854 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1555  (
    .i0(\u2_Display/n820 ),
    .i1(\u2_Display/n839 [16]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n855 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1556  (
    .i0(\u2_Display/n821 ),
    .i1(\u2_Display/n839 [15]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n856 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1557  (
    .i0(\u2_Display/n822 ),
    .i1(\u2_Display/n839 [14]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n857 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1558  (
    .i0(\u2_Display/n823 ),
    .i1(\u2_Display/n839 [13]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n858 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1559  (
    .i0(\u2_Display/n824 ),
    .i1(\u2_Display/n839 [12]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n859 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1560  (
    .i0(\u2_Display/n825 ),
    .i1(\u2_Display/n839 [11]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n860 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1561  (
    .i0(\u2_Display/n826 ),
    .i1(\u2_Display/n839 [10]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n861 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1562  (
    .i0(\u2_Display/n827 ),
    .i1(\u2_Display/n839 [9]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n862 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1563  (
    .i0(\u2_Display/n828 ),
    .i1(\u2_Display/n839 [8]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n863 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1564  (
    .i0(\u2_Display/n829 ),
    .i1(\u2_Display/n839 [7]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n864 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1565  (
    .i0(\u2_Display/n830 ),
    .i1(\u2_Display/n839 [6]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n865 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1566  (
    .i0(\u2_Display/n831 ),
    .i1(\u2_Display/n839 [5]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n866 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1567  (
    .i0(\u2_Display/n832 ),
    .i1(\u2_Display/n839 [4]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n867 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1568  (
    .i0(\u2_Display/n833 ),
    .i1(\u2_Display/n839 [3]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n868 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1569  (
    .i0(\u2_Display/n834 ),
    .i1(\u2_Display/n839 [2]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n869 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1570  (
    .i0(\u2_Display/n835 ),
    .i1(\u2_Display/n839 [1]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n870 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1571  (
    .i0(\u2_Display/n836 ),
    .i1(\u2_Display/n839 [0]),
    .sel(\u2_Display/n838 ),
    .o(\u2_Display/n871 ));  // source/rtl/Display.v(230)
  not \u2_Display/u1572  (\u2_Display/n873 , \u2_Display/n872 );  // source/rtl/Display.v(230)
  and \u2_Display/u16  (\u2_Display/n101 , \u2_Display/n98 , \u2_Display/n100 );  // source/rtl/Display.v(181)
  AL_MUX \u2_Display/u1605  (
    .i0(\u2_Display/n840 ),
    .i1(\u2_Display/n874 [31]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n875 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1606  (
    .i0(\u2_Display/n841 ),
    .i1(\u2_Display/n874 [30]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n876 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1607  (
    .i0(\u2_Display/n842 ),
    .i1(\u2_Display/n874 [29]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n877 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1608  (
    .i0(\u2_Display/n843 ),
    .i1(\u2_Display/n874 [28]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n878 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1609  (
    .i0(\u2_Display/n844 ),
    .i1(\u2_Display/n874 [27]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n879 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1610  (
    .i0(\u2_Display/n845 ),
    .i1(\u2_Display/n874 [26]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n880 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1611  (
    .i0(\u2_Display/n846 ),
    .i1(\u2_Display/n874 [25]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n881 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1612  (
    .i0(\u2_Display/n847 ),
    .i1(\u2_Display/n874 [24]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n882 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1613  (
    .i0(\u2_Display/n848 ),
    .i1(\u2_Display/n874 [23]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n883 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1614  (
    .i0(\u2_Display/n849 ),
    .i1(\u2_Display/n874 [22]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n884 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1615  (
    .i0(\u2_Display/n850 ),
    .i1(\u2_Display/n874 [21]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n885 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1616  (
    .i0(\u2_Display/n851 ),
    .i1(\u2_Display/n874 [20]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n886 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1617  (
    .i0(\u2_Display/n852 ),
    .i1(\u2_Display/n874 [19]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n887 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1618  (
    .i0(\u2_Display/n853 ),
    .i1(\u2_Display/n874 [18]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n888 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1619  (
    .i0(\u2_Display/n854 ),
    .i1(\u2_Display/n874 [17]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n889 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1620  (
    .i0(\u2_Display/n855 ),
    .i1(\u2_Display/n874 [16]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n890 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1621  (
    .i0(\u2_Display/n856 ),
    .i1(\u2_Display/n874 [15]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n891 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1622  (
    .i0(\u2_Display/n857 ),
    .i1(\u2_Display/n874 [14]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n892 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1623  (
    .i0(\u2_Display/n858 ),
    .i1(\u2_Display/n874 [13]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n893 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1624  (
    .i0(\u2_Display/n859 ),
    .i1(\u2_Display/n874 [12]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n894 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1625  (
    .i0(\u2_Display/n860 ),
    .i1(\u2_Display/n874 [11]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n895 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1626  (
    .i0(\u2_Display/n861 ),
    .i1(\u2_Display/n874 [10]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n896 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1627  (
    .i0(\u2_Display/n862 ),
    .i1(\u2_Display/n874 [9]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n897 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1628  (
    .i0(\u2_Display/n863 ),
    .i1(\u2_Display/n874 [8]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n898 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1629  (
    .i0(\u2_Display/n864 ),
    .i1(\u2_Display/n874 [7]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n899 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1630  (
    .i0(\u2_Display/n865 ),
    .i1(\u2_Display/n874 [6]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n900 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1631  (
    .i0(\u2_Display/n866 ),
    .i1(\u2_Display/n874 [5]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n901 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1632  (
    .i0(\u2_Display/n867 ),
    .i1(\u2_Display/n874 [4]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n902 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1633  (
    .i0(\u2_Display/n868 ),
    .i1(\u2_Display/n874 [3]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n903 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1634  (
    .i0(\u2_Display/n869 ),
    .i1(\u2_Display/n874 [2]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n904 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1635  (
    .i0(\u2_Display/n870 ),
    .i1(\u2_Display/n874 [1]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n905 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1636  (
    .i0(\u2_Display/n871 ),
    .i1(\u2_Display/n874 [0]),
    .sel(\u2_Display/n873 ),
    .o(\u2_Display/n906 ));  // source/rtl/Display.v(230)
  not \u2_Display/u1637  (\u2_Display/n908 , \u2_Display/n907 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1670  (
    .i0(\u2_Display/n875 ),
    .i1(\u2_Display/n909 [31]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n910 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1671  (
    .i0(\u2_Display/n876 ),
    .i1(\u2_Display/n909 [30]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n911 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1672  (
    .i0(\u2_Display/n877 ),
    .i1(\u2_Display/n909 [29]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n912 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1673  (
    .i0(\u2_Display/n878 ),
    .i1(\u2_Display/n909 [28]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n913 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1674  (
    .i0(\u2_Display/n879 ),
    .i1(\u2_Display/n909 [27]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n914 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1675  (
    .i0(\u2_Display/n880 ),
    .i1(\u2_Display/n909 [26]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n915 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1676  (
    .i0(\u2_Display/n881 ),
    .i1(\u2_Display/n909 [25]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n916 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1677  (
    .i0(\u2_Display/n882 ),
    .i1(\u2_Display/n909 [24]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n917 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1678  (
    .i0(\u2_Display/n883 ),
    .i1(\u2_Display/n909 [23]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n918 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1679  (
    .i0(\u2_Display/n884 ),
    .i1(\u2_Display/n909 [22]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n919 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1680  (
    .i0(\u2_Display/n885 ),
    .i1(\u2_Display/n909 [21]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n920 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1681  (
    .i0(\u2_Display/n886 ),
    .i1(\u2_Display/n909 [20]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n921 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1682  (
    .i0(\u2_Display/n887 ),
    .i1(\u2_Display/n909 [19]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n922 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1683  (
    .i0(\u2_Display/n888 ),
    .i1(\u2_Display/n909 [18]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n923 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1684  (
    .i0(\u2_Display/n889 ),
    .i1(\u2_Display/n909 [17]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n924 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1685  (
    .i0(\u2_Display/n890 ),
    .i1(\u2_Display/n909 [16]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n925 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1686  (
    .i0(\u2_Display/n891 ),
    .i1(\u2_Display/n909 [15]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n926 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1687  (
    .i0(\u2_Display/n892 ),
    .i1(\u2_Display/n909 [14]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n927 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1688  (
    .i0(\u2_Display/n893 ),
    .i1(\u2_Display/n909 [13]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n928 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1689  (
    .i0(\u2_Display/n894 ),
    .i1(\u2_Display/n909 [12]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n929 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1690  (
    .i0(\u2_Display/n895 ),
    .i1(\u2_Display/n909 [11]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n930 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1691  (
    .i0(\u2_Display/n896 ),
    .i1(\u2_Display/n909 [10]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n931 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1692  (
    .i0(\u2_Display/n897 ),
    .i1(\u2_Display/n909 [9]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n932 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1693  (
    .i0(\u2_Display/n898 ),
    .i1(\u2_Display/n909 [8]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n933 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1694  (
    .i0(\u2_Display/n899 ),
    .i1(\u2_Display/n909 [7]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n934 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1695  (
    .i0(\u2_Display/n900 ),
    .i1(\u2_Display/n909 [6]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n935 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1696  (
    .i0(\u2_Display/n901 ),
    .i1(\u2_Display/n909 [5]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n936 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1697  (
    .i0(\u2_Display/n902 ),
    .i1(\u2_Display/n909 [4]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n937 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1698  (
    .i0(\u2_Display/n903 ),
    .i1(\u2_Display/n909 [3]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n938 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1699  (
    .i0(\u2_Display/n904 ),
    .i1(\u2_Display/n909 [2]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n939 ));  // source/rtl/Display.v(230)
  and \u2_Display/u17  (\u2_Display/n104 , \u2_Display/n101 , \u2_Display/n103 );  // source/rtl/Display.v(181)
  AL_MUX \u2_Display/u1700  (
    .i0(\u2_Display/n905 ),
    .i1(\u2_Display/n909 [1]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n940 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1701  (
    .i0(\u2_Display/n906 ),
    .i1(\u2_Display/n909 [0]),
    .sel(\u2_Display/n908 ),
    .o(\u2_Display/n941 ));  // source/rtl/Display.v(230)
  not \u2_Display/u1702  (\u2_Display/n943 , \u2_Display/n942 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1735  (
    .i0(\u2_Display/n910 ),
    .i1(\u2_Display/n944 [31]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n945 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1736  (
    .i0(\u2_Display/n911 ),
    .i1(\u2_Display/n944 [30]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n946 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1737  (
    .i0(\u2_Display/n912 ),
    .i1(\u2_Display/n944 [29]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n947 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1738  (
    .i0(\u2_Display/n913 ),
    .i1(\u2_Display/n944 [28]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n948 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1739  (
    .i0(\u2_Display/n914 ),
    .i1(\u2_Display/n944 [27]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n949 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1740  (
    .i0(\u2_Display/n915 ),
    .i1(\u2_Display/n944 [26]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n950 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1741  (
    .i0(\u2_Display/n916 ),
    .i1(\u2_Display/n944 [25]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n951 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1742  (
    .i0(\u2_Display/n917 ),
    .i1(\u2_Display/n944 [24]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n952 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1743  (
    .i0(\u2_Display/n918 ),
    .i1(\u2_Display/n944 [23]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n953 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1744  (
    .i0(\u2_Display/n919 ),
    .i1(\u2_Display/n944 [22]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n954 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1745  (
    .i0(\u2_Display/n920 ),
    .i1(\u2_Display/n944 [21]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n955 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1746  (
    .i0(\u2_Display/n921 ),
    .i1(\u2_Display/n944 [20]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n956 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1747  (
    .i0(\u2_Display/n922 ),
    .i1(\u2_Display/n944 [19]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n957 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1748  (
    .i0(\u2_Display/n923 ),
    .i1(\u2_Display/n944 [18]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n958 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1749  (
    .i0(\u2_Display/n924 ),
    .i1(\u2_Display/n944 [17]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n959 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1750  (
    .i0(\u2_Display/n925 ),
    .i1(\u2_Display/n944 [16]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n960 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1751  (
    .i0(\u2_Display/n926 ),
    .i1(\u2_Display/n944 [15]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n961 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1752  (
    .i0(\u2_Display/n927 ),
    .i1(\u2_Display/n944 [14]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n962 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1753  (
    .i0(\u2_Display/n928 ),
    .i1(\u2_Display/n944 [13]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n963 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1754  (
    .i0(\u2_Display/n929 ),
    .i1(\u2_Display/n944 [12]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n964 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1755  (
    .i0(\u2_Display/n930 ),
    .i1(\u2_Display/n944 [11]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n965 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1756  (
    .i0(\u2_Display/n931 ),
    .i1(\u2_Display/n944 [10]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n966 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1757  (
    .i0(\u2_Display/n932 ),
    .i1(\u2_Display/n944 [9]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n967 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1758  (
    .i0(\u2_Display/n933 ),
    .i1(\u2_Display/n944 [8]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n968 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1759  (
    .i0(\u2_Display/n934 ),
    .i1(\u2_Display/n944 [7]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n969 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1760  (
    .i0(\u2_Display/n935 ),
    .i1(\u2_Display/n944 [6]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n970 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1761  (
    .i0(\u2_Display/n936 ),
    .i1(\u2_Display/n944 [5]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n971 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1762  (
    .i0(\u2_Display/n937 ),
    .i1(\u2_Display/n944 [4]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n972 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1763  (
    .i0(\u2_Display/n938 ),
    .i1(\u2_Display/n944 [3]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n973 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1764  (
    .i0(\u2_Display/n939 ),
    .i1(\u2_Display/n944 [2]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n974 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1765  (
    .i0(\u2_Display/n940 ),
    .i1(\u2_Display/n944 [1]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n975 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1766  (
    .i0(\u2_Display/n941 ),
    .i1(\u2_Display/n944 [0]),
    .sel(\u2_Display/n943 ),
    .o(\u2_Display/n976 ));  // source/rtl/Display.v(230)
  not \u2_Display/u1767  (\u2_Display/n978 , \u2_Display/n977 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1800  (
    .i0(\u2_Display/n945 ),
    .i1(\u2_Display/n979 [31]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n980 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1801  (
    .i0(\u2_Display/n946 ),
    .i1(\u2_Display/n979 [30]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n981 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1802  (
    .i0(\u2_Display/n947 ),
    .i1(\u2_Display/n979 [29]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n982 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1803  (
    .i0(\u2_Display/n948 ),
    .i1(\u2_Display/n979 [28]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n983 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1804  (
    .i0(\u2_Display/n949 ),
    .i1(\u2_Display/n979 [27]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n984 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1805  (
    .i0(\u2_Display/n950 ),
    .i1(\u2_Display/n979 [26]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n985 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1806  (
    .i0(\u2_Display/n951 ),
    .i1(\u2_Display/n979 [25]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n986 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1807  (
    .i0(\u2_Display/n952 ),
    .i1(\u2_Display/n979 [24]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n987 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1808  (
    .i0(\u2_Display/n953 ),
    .i1(\u2_Display/n979 [23]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n988 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1809  (
    .i0(\u2_Display/n954 ),
    .i1(\u2_Display/n979 [22]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n989 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1810  (
    .i0(\u2_Display/n955 ),
    .i1(\u2_Display/n979 [21]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n990 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1811  (
    .i0(\u2_Display/n956 ),
    .i1(\u2_Display/n979 [20]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n991 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1812  (
    .i0(\u2_Display/n957 ),
    .i1(\u2_Display/n979 [19]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n992 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1813  (
    .i0(\u2_Display/n958 ),
    .i1(\u2_Display/n979 [18]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n993 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1814  (
    .i0(\u2_Display/n959 ),
    .i1(\u2_Display/n979 [17]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n994 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1815  (
    .i0(\u2_Display/n960 ),
    .i1(\u2_Display/n979 [16]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n995 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1816  (
    .i0(\u2_Display/n961 ),
    .i1(\u2_Display/n979 [15]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n996 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1817  (
    .i0(\u2_Display/n962 ),
    .i1(\u2_Display/n979 [14]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n997 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1818  (
    .i0(\u2_Display/n963 ),
    .i1(\u2_Display/n979 [13]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n998 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1819  (
    .i0(\u2_Display/n964 ),
    .i1(\u2_Display/n979 [12]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n999 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1820  (
    .i0(\u2_Display/n965 ),
    .i1(\u2_Display/n979 [11]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n1000 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1821  (
    .i0(\u2_Display/n966 ),
    .i1(\u2_Display/n979 [10]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n1001 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1822  (
    .i0(\u2_Display/n967 ),
    .i1(\u2_Display/n979 [9]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n1002 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1823  (
    .i0(\u2_Display/n968 ),
    .i1(\u2_Display/n979 [8]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n1003 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1824  (
    .i0(\u2_Display/n969 ),
    .i1(\u2_Display/n979 [7]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n1004 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1825  (
    .i0(\u2_Display/n970 ),
    .i1(\u2_Display/n979 [6]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n1005 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1826  (
    .i0(\u2_Display/n971 ),
    .i1(\u2_Display/n979 [5]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n1006 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1827  (
    .i0(\u2_Display/n972 ),
    .i1(\u2_Display/n979 [4]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n1007 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1828  (
    .i0(\u2_Display/n973 ),
    .i1(\u2_Display/n979 [3]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n1008 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1829  (
    .i0(\u2_Display/n974 ),
    .i1(\u2_Display/n979 [2]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n1009 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1830  (
    .i0(\u2_Display/n975 ),
    .i1(\u2_Display/n979 [1]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n1010 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1831  (
    .i0(\u2_Display/n976 ),
    .i1(\u2_Display/n979 [0]),
    .sel(\u2_Display/n978 ),
    .o(\u2_Display/n1011 ));  // source/rtl/Display.v(230)
  not \u2_Display/u1832  (\u2_Display/n1013 , \u2_Display/n1012 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1865  (
    .i0(\u2_Display/n980 ),
    .i1(\u2_Display/n1014 [31]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1015 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1866  (
    .i0(\u2_Display/n981 ),
    .i1(\u2_Display/n1014 [30]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1016 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1867  (
    .i0(\u2_Display/n982 ),
    .i1(\u2_Display/n1014 [29]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1017 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1868  (
    .i0(\u2_Display/n983 ),
    .i1(\u2_Display/n1014 [28]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1018 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1869  (
    .i0(\u2_Display/n984 ),
    .i1(\u2_Display/n1014 [27]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1019 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1870  (
    .i0(\u2_Display/n985 ),
    .i1(\u2_Display/n1014 [26]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1020 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1871  (
    .i0(\u2_Display/n986 ),
    .i1(\u2_Display/n1014 [25]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1021 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1872  (
    .i0(\u2_Display/n987 ),
    .i1(\u2_Display/n1014 [24]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1022 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1873  (
    .i0(\u2_Display/n988 ),
    .i1(\u2_Display/n1014 [23]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1023 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1874  (
    .i0(\u2_Display/n989 ),
    .i1(\u2_Display/n1014 [22]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1024 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1875  (
    .i0(\u2_Display/n990 ),
    .i1(\u2_Display/n1014 [21]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1025 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1876  (
    .i0(\u2_Display/n991 ),
    .i1(\u2_Display/n1014 [20]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1026 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1877  (
    .i0(\u2_Display/n992 ),
    .i1(\u2_Display/n1014 [19]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1027 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1878  (
    .i0(\u2_Display/n993 ),
    .i1(\u2_Display/n1014 [18]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1028 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1879  (
    .i0(\u2_Display/n994 ),
    .i1(\u2_Display/n1014 [17]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1029 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1880  (
    .i0(\u2_Display/n995 ),
    .i1(\u2_Display/n1014 [16]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1030 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1881  (
    .i0(\u2_Display/n996 ),
    .i1(\u2_Display/n1014 [15]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1031 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1882  (
    .i0(\u2_Display/n997 ),
    .i1(\u2_Display/n1014 [14]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1032 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1883  (
    .i0(\u2_Display/n998 ),
    .i1(\u2_Display/n1014 [13]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1033 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1884  (
    .i0(\u2_Display/n999 ),
    .i1(\u2_Display/n1014 [12]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1034 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1885  (
    .i0(\u2_Display/n1000 ),
    .i1(\u2_Display/n1014 [11]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1035 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1886  (
    .i0(\u2_Display/n1001 ),
    .i1(\u2_Display/n1014 [10]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1036 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1887  (
    .i0(\u2_Display/n1002 ),
    .i1(\u2_Display/n1014 [9]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1037 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1888  (
    .i0(\u2_Display/n1003 ),
    .i1(\u2_Display/n1014 [8]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1038 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1889  (
    .i0(\u2_Display/n1004 ),
    .i1(\u2_Display/n1014 [7]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1039 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1890  (
    .i0(\u2_Display/n1005 ),
    .i1(\u2_Display/n1014 [6]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1040 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1891  (
    .i0(\u2_Display/n1006 ),
    .i1(\u2_Display/n1014 [5]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1041 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1892  (
    .i0(\u2_Display/n1007 ),
    .i1(\u2_Display/n1014 [4]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1042 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1893  (
    .i0(\u2_Display/n1008 ),
    .i1(\u2_Display/n1014 [3]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1043 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1894  (
    .i0(\u2_Display/n1009 ),
    .i1(\u2_Display/n1014 [2]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1044 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1895  (
    .i0(\u2_Display/n1010 ),
    .i1(\u2_Display/n1014 [1]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1045 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1896  (
    .i0(\u2_Display/n1011 ),
    .i1(\u2_Display/n1014 [0]),
    .sel(\u2_Display/n1013 ),
    .o(\u2_Display/n1046 ));  // source/rtl/Display.v(230)
  not \u2_Display/u1897  (\u2_Display/n1048 , \u2_Display/n1047 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1930  (
    .i0(\u2_Display/n1015 ),
    .i1(\u2_Display/n1049 [31]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1050 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1931  (
    .i0(\u2_Display/n1016 ),
    .i1(\u2_Display/n1049 [30]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1051 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1932  (
    .i0(\u2_Display/n1017 ),
    .i1(\u2_Display/n1049 [29]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1052 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1933  (
    .i0(\u2_Display/n1018 ),
    .i1(\u2_Display/n1049 [28]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1053 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1934  (
    .i0(\u2_Display/n1019 ),
    .i1(\u2_Display/n1049 [27]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1054 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1935  (
    .i0(\u2_Display/n1020 ),
    .i1(\u2_Display/n1049 [26]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1055 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1936  (
    .i0(\u2_Display/n1021 ),
    .i1(\u2_Display/n1049 [25]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1056 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1937  (
    .i0(\u2_Display/n1022 ),
    .i1(\u2_Display/n1049 [24]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1057 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1938  (
    .i0(\u2_Display/n1023 ),
    .i1(\u2_Display/n1049 [23]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1058 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1939  (
    .i0(\u2_Display/n1024 ),
    .i1(\u2_Display/n1049 [22]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1059 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1940  (
    .i0(\u2_Display/n1025 ),
    .i1(\u2_Display/n1049 [21]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1060 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1941  (
    .i0(\u2_Display/n1026 ),
    .i1(\u2_Display/n1049 [20]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1061 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1942  (
    .i0(\u2_Display/n1027 ),
    .i1(\u2_Display/n1049 [19]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1062 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1943  (
    .i0(\u2_Display/n1028 ),
    .i1(\u2_Display/n1049 [18]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1063 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1944  (
    .i0(\u2_Display/n1029 ),
    .i1(\u2_Display/n1049 [17]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1064 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1945  (
    .i0(\u2_Display/n1030 ),
    .i1(\u2_Display/n1049 [16]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1065 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1946  (
    .i0(\u2_Display/n1031 ),
    .i1(\u2_Display/n1049 [15]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1066 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1947  (
    .i0(\u2_Display/n1032 ),
    .i1(\u2_Display/n1049 [14]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1067 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1948  (
    .i0(\u2_Display/n1033 ),
    .i1(\u2_Display/n1049 [13]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1068 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1949  (
    .i0(\u2_Display/n1034 ),
    .i1(\u2_Display/n1049 [12]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1069 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1950  (
    .i0(\u2_Display/n1035 ),
    .i1(\u2_Display/n1049 [11]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1070 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1951  (
    .i0(\u2_Display/n1036 ),
    .i1(\u2_Display/n1049 [10]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1071 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1952  (
    .i0(\u2_Display/n1037 ),
    .i1(\u2_Display/n1049 [9]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1072 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1953  (
    .i0(\u2_Display/n1038 ),
    .i1(\u2_Display/n1049 [8]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1073 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1954  (
    .i0(\u2_Display/n1039 ),
    .i1(\u2_Display/n1049 [7]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1074 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1955  (
    .i0(\u2_Display/n1040 ),
    .i1(\u2_Display/n1049 [6]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1075 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1956  (
    .i0(\u2_Display/n1041 ),
    .i1(\u2_Display/n1049 [5]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1076 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1957  (
    .i0(\u2_Display/n1042 ),
    .i1(\u2_Display/n1049 [4]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1077 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1958  (
    .i0(\u2_Display/n1043 ),
    .i1(\u2_Display/n1049 [3]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1078 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1959  (
    .i0(\u2_Display/n1044 ),
    .i1(\u2_Display/n1049 [2]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1079 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1960  (
    .i0(\u2_Display/n1045 ),
    .i1(\u2_Display/n1049 [1]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1080 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1961  (
    .i0(\u2_Display/n1046 ),
    .i1(\u2_Display/n1049 [0]),
    .sel(\u2_Display/n1048 ),
    .o(\u2_Display/n1081 ));  // source/rtl/Display.v(230)
  not \u2_Display/u1962  (\u2_Display/n1083 , \u2_Display/n1082 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1995  (
    .i0(\u2_Display/n1050 ),
    .i1(\u2_Display/n1084 [31]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1085 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1996  (
    .i0(\u2_Display/n1051 ),
    .i1(\u2_Display/n1084 [30]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1086 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1997  (
    .i0(\u2_Display/n1052 ),
    .i1(\u2_Display/n1084 [29]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1087 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1998  (
    .i0(\u2_Display/n1053 ),
    .i1(\u2_Display/n1084 [28]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1088 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u1999  (
    .i0(\u2_Display/n1054 ),
    .i1(\u2_Display/n1084 [27]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1089 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2000  (
    .i0(\u2_Display/n1055 ),
    .i1(\u2_Display/n1084 [26]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1090 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2001  (
    .i0(\u2_Display/n1056 ),
    .i1(\u2_Display/n1084 [25]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1091 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2002  (
    .i0(\u2_Display/n1057 ),
    .i1(\u2_Display/n1084 [24]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1092 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2003  (
    .i0(\u2_Display/n1058 ),
    .i1(\u2_Display/n1084 [23]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1093 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2004  (
    .i0(\u2_Display/n1059 ),
    .i1(\u2_Display/n1084 [22]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1094 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2005  (
    .i0(\u2_Display/n1060 ),
    .i1(\u2_Display/n1084 [21]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1095 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2006  (
    .i0(\u2_Display/n1061 ),
    .i1(\u2_Display/n1084 [20]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1096 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2007  (
    .i0(\u2_Display/n1062 ),
    .i1(\u2_Display/n1084 [19]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1097 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2008  (
    .i0(\u2_Display/n1063 ),
    .i1(\u2_Display/n1084 [18]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1098 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2009  (
    .i0(\u2_Display/n1064 ),
    .i1(\u2_Display/n1084 [17]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1099 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2010  (
    .i0(\u2_Display/n1065 ),
    .i1(\u2_Display/n1084 [16]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1100 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2011  (
    .i0(\u2_Display/n1066 ),
    .i1(\u2_Display/n1084 [15]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1101 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2012  (
    .i0(\u2_Display/n1067 ),
    .i1(\u2_Display/n1084 [14]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1102 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2013  (
    .i0(\u2_Display/n1068 ),
    .i1(\u2_Display/n1084 [13]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1103 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2014  (
    .i0(\u2_Display/n1069 ),
    .i1(\u2_Display/n1084 [12]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1104 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2015  (
    .i0(\u2_Display/n1070 ),
    .i1(\u2_Display/n1084 [11]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1105 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2016  (
    .i0(\u2_Display/n1071 ),
    .i1(\u2_Display/n1084 [10]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1106 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2017  (
    .i0(\u2_Display/n1072 ),
    .i1(\u2_Display/n1084 [9]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1107 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2018  (
    .i0(\u2_Display/n1073 ),
    .i1(\u2_Display/n1084 [8]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1108 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2019  (
    .i0(\u2_Display/n1074 ),
    .i1(\u2_Display/n1084 [7]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1109 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2020  (
    .i0(\u2_Display/n1075 ),
    .i1(\u2_Display/n1084 [6]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1110 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2021  (
    .i0(\u2_Display/n1076 ),
    .i1(\u2_Display/n1084 [5]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1111 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2022  (
    .i0(\u2_Display/n1077 ),
    .i1(\u2_Display/n1084 [4]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1112 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2023  (
    .i0(\u2_Display/n1078 ),
    .i1(\u2_Display/n1084 [3]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1113 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2024  (
    .i0(\u2_Display/n1079 ),
    .i1(\u2_Display/n1084 [2]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1114 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2025  (
    .i0(\u2_Display/n1080 ),
    .i1(\u2_Display/n1084 [1]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1115 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2026  (
    .i0(\u2_Display/n1081 ),
    .i1(\u2_Display/n1084 [0]),
    .sel(\u2_Display/n1083 ),
    .o(\u2_Display/n1116 ));  // source/rtl/Display.v(230)
  not \u2_Display/u2027  (\u2_Display/n1118 , \u2_Display/n1117 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2060  (
    .i0(\u2_Display/n1085 ),
    .i1(\u2_Display/n1119 [31]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1120 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2061  (
    .i0(\u2_Display/n1086 ),
    .i1(\u2_Display/n1119 [30]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1121 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2062  (
    .i0(\u2_Display/n1087 ),
    .i1(\u2_Display/n1119 [29]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1122 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2063  (
    .i0(\u2_Display/n1088 ),
    .i1(\u2_Display/n1119 [28]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1123 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2064  (
    .i0(\u2_Display/n1089 ),
    .i1(\u2_Display/n1119 [27]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1124 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2065  (
    .i0(\u2_Display/n1090 ),
    .i1(\u2_Display/n1119 [26]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1125 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2066  (
    .i0(\u2_Display/n1091 ),
    .i1(\u2_Display/n1119 [25]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1126 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2067  (
    .i0(\u2_Display/n1092 ),
    .i1(\u2_Display/n1119 [24]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1127 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2068  (
    .i0(\u2_Display/n1093 ),
    .i1(\u2_Display/n1119 [23]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1128 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2069  (
    .i0(\u2_Display/n1094 ),
    .i1(\u2_Display/n1119 [22]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1129 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2070  (
    .i0(\u2_Display/n1095 ),
    .i1(\u2_Display/n1119 [21]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1130 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2071  (
    .i0(\u2_Display/n1096 ),
    .i1(\u2_Display/n1119 [20]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1131 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2072  (
    .i0(\u2_Display/n1097 ),
    .i1(\u2_Display/n1119 [19]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1132 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2073  (
    .i0(\u2_Display/n1098 ),
    .i1(\u2_Display/n1119 [18]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1133 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2074  (
    .i0(\u2_Display/n1099 ),
    .i1(\u2_Display/n1119 [17]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1134 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2075  (
    .i0(\u2_Display/n1100 ),
    .i1(\u2_Display/n1119 [16]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1135 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2076  (
    .i0(\u2_Display/n1101 ),
    .i1(\u2_Display/n1119 [15]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1136 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2077  (
    .i0(\u2_Display/n1102 ),
    .i1(\u2_Display/n1119 [14]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1137 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2078  (
    .i0(\u2_Display/n1103 ),
    .i1(\u2_Display/n1119 [13]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1138 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2079  (
    .i0(\u2_Display/n1104 ),
    .i1(\u2_Display/n1119 [12]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1139 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2080  (
    .i0(\u2_Display/n1105 ),
    .i1(\u2_Display/n1119 [11]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1140 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2081  (
    .i0(\u2_Display/n1106 ),
    .i1(\u2_Display/n1119 [10]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1141 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2082  (
    .i0(\u2_Display/n1107 ),
    .i1(\u2_Display/n1119 [9]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1142 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2083  (
    .i0(\u2_Display/n1108 ),
    .i1(\u2_Display/n1119 [8]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1143 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2084  (
    .i0(\u2_Display/n1109 ),
    .i1(\u2_Display/n1119 [7]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1144 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2085  (
    .i0(\u2_Display/n1110 ),
    .i1(\u2_Display/n1119 [6]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1145 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2086  (
    .i0(\u2_Display/n1111 ),
    .i1(\u2_Display/n1119 [5]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1146 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2087  (
    .i0(\u2_Display/n1112 ),
    .i1(\u2_Display/n1119 [4]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1147 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2088  (
    .i0(\u2_Display/n1113 ),
    .i1(\u2_Display/n1119 [3]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1148 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2089  (
    .i0(\u2_Display/n1114 ),
    .i1(\u2_Display/n1119 [2]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1149 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2090  (
    .i0(\u2_Display/n1115 ),
    .i1(\u2_Display/n1119 [1]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1150 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2091  (
    .i0(\u2_Display/n1116 ),
    .i1(\u2_Display/n1119 [0]),
    .sel(\u2_Display/n1118 ),
    .o(\u2_Display/n1151 ));  // source/rtl/Display.v(230)
  not \u2_Display/u2092  (\u2_Display/n1153 , \u2_Display/n1152 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2125  (
    .i0(\u2_Display/n1120 ),
    .i1(\u2_Display/n1154 [31]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1155 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2126  (
    .i0(\u2_Display/n1121 ),
    .i1(\u2_Display/n1154 [30]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1156 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2127  (
    .i0(\u2_Display/n1122 ),
    .i1(\u2_Display/n1154 [29]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1157 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2128  (
    .i0(\u2_Display/n1123 ),
    .i1(\u2_Display/n1154 [28]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1158 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2129  (
    .i0(\u2_Display/n1124 ),
    .i1(\u2_Display/n1154 [27]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1159 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2130  (
    .i0(\u2_Display/n1125 ),
    .i1(\u2_Display/n1154 [26]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1160 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2131  (
    .i0(\u2_Display/n1126 ),
    .i1(\u2_Display/n1154 [25]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1161 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2132  (
    .i0(\u2_Display/n1127 ),
    .i1(\u2_Display/n1154 [24]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1162 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2133  (
    .i0(\u2_Display/n1128 ),
    .i1(\u2_Display/n1154 [23]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1163 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2134  (
    .i0(\u2_Display/n1129 ),
    .i1(\u2_Display/n1154 [22]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1164 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2135  (
    .i0(\u2_Display/n1130 ),
    .i1(\u2_Display/n1154 [21]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1165 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2136  (
    .i0(\u2_Display/n1131 ),
    .i1(\u2_Display/n1154 [20]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1166 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2137  (
    .i0(\u2_Display/n1132 ),
    .i1(\u2_Display/n1154 [19]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1167 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2138  (
    .i0(\u2_Display/n1133 ),
    .i1(\u2_Display/n1154 [18]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1168 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2139  (
    .i0(\u2_Display/n1134 ),
    .i1(\u2_Display/n1154 [17]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1169 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2140  (
    .i0(\u2_Display/n1135 ),
    .i1(\u2_Display/n1154 [16]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1170 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2141  (
    .i0(\u2_Display/n1136 ),
    .i1(\u2_Display/n1154 [15]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1171 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2142  (
    .i0(\u2_Display/n1137 ),
    .i1(\u2_Display/n1154 [14]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1172 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2143  (
    .i0(\u2_Display/n1138 ),
    .i1(\u2_Display/n1154 [13]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1173 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2144  (
    .i0(\u2_Display/n1139 ),
    .i1(\u2_Display/n1154 [12]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1174 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2145  (
    .i0(\u2_Display/n1140 ),
    .i1(\u2_Display/n1154 [11]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1175 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2146  (
    .i0(\u2_Display/n1141 ),
    .i1(\u2_Display/n1154 [10]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1176 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2147  (
    .i0(\u2_Display/n1142 ),
    .i1(\u2_Display/n1154 [9]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1177 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2148  (
    .i0(\u2_Display/n1143 ),
    .i1(\u2_Display/n1154 [8]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1178 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2149  (
    .i0(\u2_Display/n1144 ),
    .i1(\u2_Display/n1154 [7]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1179 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2150  (
    .i0(\u2_Display/n1145 ),
    .i1(\u2_Display/n1154 [6]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1180 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2151  (
    .i0(\u2_Display/n1146 ),
    .i1(\u2_Display/n1154 [5]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1181 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2152  (
    .i0(\u2_Display/n1147 ),
    .i1(\u2_Display/n1154 [4]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1182 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2153  (
    .i0(\u2_Display/n1148 ),
    .i1(\u2_Display/n1154 [3]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1183 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2154  (
    .i0(\u2_Display/n1149 ),
    .i1(\u2_Display/n1154 [2]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1184 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2155  (
    .i0(\u2_Display/n1150 ),
    .i1(\u2_Display/n1154 [1]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1185 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2156  (
    .i0(\u2_Display/n1151 ),
    .i1(\u2_Display/n1154 [0]),
    .sel(\u2_Display/n1153 ),
    .o(\u2_Display/n1186 ));  // source/rtl/Display.v(230)
  not \u2_Display/u2157  (\u2_Display/n1188 , \u2_Display/n1187 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2190  (
    .i0(\u2_Display/n1177 ),
    .i1(\u2_Display/n1189 [9]),
    .sel(\u2_Display/n1188 ),
    .o(\u2_Display/n196 [9]));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2191  (
    .i0(\u2_Display/n1178 ),
    .i1(\u2_Display/n1189 [8]),
    .sel(\u2_Display/n1188 ),
    .o(\u2_Display/n196 [8]));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2192  (
    .i0(\u2_Display/n1179 ),
    .i1(\u2_Display/n1189 [7]),
    .sel(\u2_Display/n1188 ),
    .o(\u2_Display/n196 [7]));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2193  (
    .i0(\u2_Display/n1180 ),
    .i1(\u2_Display/n1189 [6]),
    .sel(\u2_Display/n1188 ),
    .o(\u2_Display/n196 [6]));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2194  (
    .i0(\u2_Display/n1181 ),
    .i1(\u2_Display/n1189 [5]),
    .sel(\u2_Display/n1188 ),
    .o(\u2_Display/n196 [5]));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2195  (
    .i0(\u2_Display/n1182 ),
    .i1(\u2_Display/n1189 [4]),
    .sel(\u2_Display/n1188 ),
    .o(\u2_Display/n196 [4]));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2196  (
    .i0(\u2_Display/n1183 ),
    .i1(\u2_Display/n1189 [3]),
    .sel(\u2_Display/n1188 ),
    .o(\u2_Display/n196 [3]));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2197  (
    .i0(\u2_Display/n1184 ),
    .i1(\u2_Display/n1189 [2]),
    .sel(\u2_Display/n1188 ),
    .o(\u2_Display/n196 [2]));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2198  (
    .i0(\u2_Display/n1185 ),
    .i1(\u2_Display/n1189 [1]),
    .sel(\u2_Display/n1188 ),
    .o(\u2_Display/n196 [1]));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u2199  (
    .i0(\u2_Display/n1186 ),
    .i1(\u2_Display/n1189 [0]),
    .sel(\u2_Display/n1188 ),
    .o(\u2_Display/n196 [0]));  // source/rtl/Display.v(230)
  and \u2_Display/u22  (\u2_Display/n139 , \u2_Display/n136 , \u2_Display/n138 );  // source/rtl/Display.v(197)
  and \u2_Display/u23  (\u2_Display/n142 , \u2_Display/n139 , \u2_Display/n141 );  // source/rtl/Display.v(197)
  and \u2_Display/u24  (\u2_Display/n145 , \u2_Display/n142 , \u2_Display/n144 );  // source/rtl/Display.v(197)
  not \u2_Display/u2906  (\u2_Display/n1541 , \u2_Display/n1540 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2939  (
    .i0(\u2_Display/counta [31]),
    .i1(\u2_Display/n1542 [31]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1543 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2940  (
    .i0(\u2_Display/counta [30]),
    .i1(\u2_Display/n1542 [30]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1544 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2941  (
    .i0(\u2_Display/counta [29]),
    .i1(\u2_Display/n1542 [29]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1545 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2942  (
    .i0(\u2_Display/counta [28]),
    .i1(\u2_Display/n1542 [28]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1546 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2943  (
    .i0(\u2_Display/counta [27]),
    .i1(\u2_Display/n1542 [27]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1547 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2944  (
    .i0(\u2_Display/counta [26]),
    .i1(\u2_Display/n1542 [26]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1548 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2945  (
    .i0(\u2_Display/counta [25]),
    .i1(\u2_Display/n1542 [25]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1549 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2946  (
    .i0(\u2_Display/counta [24]),
    .i1(\u2_Display/n1542 [24]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1550 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2947  (
    .i0(\u2_Display/counta [23]),
    .i1(\u2_Display/n1542 [23]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1551 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2948  (
    .i0(\u2_Display/counta [22]),
    .i1(\u2_Display/n1542 [22]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1552 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2949  (
    .i0(\u2_Display/counta [21]),
    .i1(\u2_Display/n1542 [21]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1553 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2950  (
    .i0(\u2_Display/counta [20]),
    .i1(\u2_Display/n1542 [20]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1554 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2951  (
    .i0(\u2_Display/counta [19]),
    .i1(\u2_Display/n1542 [19]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1555 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2952  (
    .i0(\u2_Display/counta [18]),
    .i1(\u2_Display/n1542 [18]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1556 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2953  (
    .i0(\u2_Display/counta [17]),
    .i1(\u2_Display/n1542 [17]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1557 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2954  (
    .i0(\u2_Display/counta [16]),
    .i1(\u2_Display/n1542 [16]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1558 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2955  (
    .i0(\u2_Display/counta [15]),
    .i1(\u2_Display/n1542 [15]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1559 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2956  (
    .i0(\u2_Display/counta [14]),
    .i1(\u2_Display/n1542 [14]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1560 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2957  (
    .i0(\u2_Display/counta [13]),
    .i1(\u2_Display/n1542 [13]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1561 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2958  (
    .i0(\u2_Display/counta [12]),
    .i1(\u2_Display/n1542 [12]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1562 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2959  (
    .i0(\u2_Display/counta [11]),
    .i1(\u2_Display/n1542 [11]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1563 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2960  (
    .i0(\u2_Display/counta [10]),
    .i1(\u2_Display/n1542 [10]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1564 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2961  (
    .i0(\u2_Display/counta [9]),
    .i1(\u2_Display/n1542 [9]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1565 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2962  (
    .i0(\u2_Display/counta [8]),
    .i1(\u2_Display/n1542 [8]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1566 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2963  (
    .i0(\u2_Display/counta [7]),
    .i1(\u2_Display/n1542 [7]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1567 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2964  (
    .i0(\u2_Display/counta [6]),
    .i1(\u2_Display/n1542 [6]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1568 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2965  (
    .i0(\u2_Display/counta [5]),
    .i1(\u2_Display/n1542 [5]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1569 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2966  (
    .i0(\u2_Display/counta [4]),
    .i1(\u2_Display/n1542 [4]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1570 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2967  (
    .i0(\u2_Display/counta [3]),
    .i1(\u2_Display/n1542 [3]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1571 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2968  (
    .i0(\u2_Display/counta [2]),
    .i1(\u2_Display/n1542 [2]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1572 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2969  (
    .i0(\u2_Display/counta [1]),
    .i1(\u2_Display/n1542 [1]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1573 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u2970  (
    .i0(\u2_Display/counta [0]),
    .i1(\u2_Display/n1542 [0]),
    .sel(\u2_Display/n1541 ),
    .o(\u2_Display/n1574 ));  // source/rtl/Display.v(213)
  not \u2_Display/u2971  (\u2_Display/n1576 , \u2_Display/n1575 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3004  (
    .i0(\u2_Display/n1543 ),
    .i1(\u2_Display/n1577 [31]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1578 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3005  (
    .i0(\u2_Display/n1544 ),
    .i1(\u2_Display/n1577 [30]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1579 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3006  (
    .i0(\u2_Display/n1545 ),
    .i1(\u2_Display/n1577 [29]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1580 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3007  (
    .i0(\u2_Display/n1546 ),
    .i1(\u2_Display/n1577 [28]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1581 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3008  (
    .i0(\u2_Display/n1547 ),
    .i1(\u2_Display/n1577 [27]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1582 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3009  (
    .i0(\u2_Display/n1548 ),
    .i1(\u2_Display/n1577 [26]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1583 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3010  (
    .i0(\u2_Display/n1549 ),
    .i1(\u2_Display/n1577 [25]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1584 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3011  (
    .i0(\u2_Display/n1550 ),
    .i1(\u2_Display/n1577 [24]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1585 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3012  (
    .i0(\u2_Display/n1551 ),
    .i1(\u2_Display/n1577 [23]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1586 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3013  (
    .i0(\u2_Display/n1552 ),
    .i1(\u2_Display/n1577 [22]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1587 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3014  (
    .i0(\u2_Display/n1553 ),
    .i1(\u2_Display/n1577 [21]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1588 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3015  (
    .i0(\u2_Display/n1554 ),
    .i1(\u2_Display/n1577 [20]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1589 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3016  (
    .i0(\u2_Display/n1555 ),
    .i1(\u2_Display/n1577 [19]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1590 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3017  (
    .i0(\u2_Display/n1556 ),
    .i1(\u2_Display/n1577 [18]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1591 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3018  (
    .i0(\u2_Display/n1557 ),
    .i1(\u2_Display/n1577 [17]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1592 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3019  (
    .i0(\u2_Display/n1558 ),
    .i1(\u2_Display/n1577 [16]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1593 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3020  (
    .i0(\u2_Display/n1559 ),
    .i1(\u2_Display/n1577 [15]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1594 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3021  (
    .i0(\u2_Display/n1560 ),
    .i1(\u2_Display/n1577 [14]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1595 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3022  (
    .i0(\u2_Display/n1561 ),
    .i1(\u2_Display/n1577 [13]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1596 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3023  (
    .i0(\u2_Display/n1562 ),
    .i1(\u2_Display/n1577 [12]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1597 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3024  (
    .i0(\u2_Display/n1563 ),
    .i1(\u2_Display/n1577 [11]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1598 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3025  (
    .i0(\u2_Display/n1564 ),
    .i1(\u2_Display/n1577 [10]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1599 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3026  (
    .i0(\u2_Display/n1565 ),
    .i1(\u2_Display/n1577 [9]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1600 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3027  (
    .i0(\u2_Display/n1566 ),
    .i1(\u2_Display/n1577 [8]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1601 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3028  (
    .i0(\u2_Display/n1567 ),
    .i1(\u2_Display/n1577 [7]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1602 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3029  (
    .i0(\u2_Display/n1568 ),
    .i1(\u2_Display/n1577 [6]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1603 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3030  (
    .i0(\u2_Display/n1569 ),
    .i1(\u2_Display/n1577 [5]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1604 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3031  (
    .i0(\u2_Display/n1570 ),
    .i1(\u2_Display/n1577 [4]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1605 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3032  (
    .i0(\u2_Display/n1571 ),
    .i1(\u2_Display/n1577 [3]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1606 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3033  (
    .i0(\u2_Display/n1572 ),
    .i1(\u2_Display/n1577 [2]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1607 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3034  (
    .i0(\u2_Display/n1573 ),
    .i1(\u2_Display/n1577 [1]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1608 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3035  (
    .i0(\u2_Display/n1574 ),
    .i1(\u2_Display/n1577 [0]),
    .sel(\u2_Display/n1576 ),
    .o(\u2_Display/n1609 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3036  (\u2_Display/n1611 , \u2_Display/n1610 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3069  (
    .i0(\u2_Display/n1578 ),
    .i1(\u2_Display/n1612 [31]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1613 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3070  (
    .i0(\u2_Display/n1579 ),
    .i1(\u2_Display/n1612 [30]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1614 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3071  (
    .i0(\u2_Display/n1580 ),
    .i1(\u2_Display/n1612 [29]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1615 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3072  (
    .i0(\u2_Display/n1581 ),
    .i1(\u2_Display/n1612 [28]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1616 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3073  (
    .i0(\u2_Display/n1582 ),
    .i1(\u2_Display/n1612 [27]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1617 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3074  (
    .i0(\u2_Display/n1583 ),
    .i1(\u2_Display/n1612 [26]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1618 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3075  (
    .i0(\u2_Display/n1584 ),
    .i1(\u2_Display/n1612 [25]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1619 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3076  (
    .i0(\u2_Display/n1585 ),
    .i1(\u2_Display/n1612 [24]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1620 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3077  (
    .i0(\u2_Display/n1586 ),
    .i1(\u2_Display/n1612 [23]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1621 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3078  (
    .i0(\u2_Display/n1587 ),
    .i1(\u2_Display/n1612 [22]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1622 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3079  (
    .i0(\u2_Display/n1588 ),
    .i1(\u2_Display/n1612 [21]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1623 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3080  (
    .i0(\u2_Display/n1589 ),
    .i1(\u2_Display/n1612 [20]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1624 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3081  (
    .i0(\u2_Display/n1590 ),
    .i1(\u2_Display/n1612 [19]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1625 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3082  (
    .i0(\u2_Display/n1591 ),
    .i1(\u2_Display/n1612 [18]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1626 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3083  (
    .i0(\u2_Display/n1592 ),
    .i1(\u2_Display/n1612 [17]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1627 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3084  (
    .i0(\u2_Display/n1593 ),
    .i1(\u2_Display/n1612 [16]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1628 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3085  (
    .i0(\u2_Display/n1594 ),
    .i1(\u2_Display/n1612 [15]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1629 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3086  (
    .i0(\u2_Display/n1595 ),
    .i1(\u2_Display/n1612 [14]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1630 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3087  (
    .i0(\u2_Display/n1596 ),
    .i1(\u2_Display/n1612 [13]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1631 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3088  (
    .i0(\u2_Display/n1597 ),
    .i1(\u2_Display/n1612 [12]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1632 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3089  (
    .i0(\u2_Display/n1598 ),
    .i1(\u2_Display/n1612 [11]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1633 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3090  (
    .i0(\u2_Display/n1599 ),
    .i1(\u2_Display/n1612 [10]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1634 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3091  (
    .i0(\u2_Display/n1600 ),
    .i1(\u2_Display/n1612 [9]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1635 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3092  (
    .i0(\u2_Display/n1601 ),
    .i1(\u2_Display/n1612 [8]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1636 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3093  (
    .i0(\u2_Display/n1602 ),
    .i1(\u2_Display/n1612 [7]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1637 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3094  (
    .i0(\u2_Display/n1603 ),
    .i1(\u2_Display/n1612 [6]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1638 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3095  (
    .i0(\u2_Display/n1604 ),
    .i1(\u2_Display/n1612 [5]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1639 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3096  (
    .i0(\u2_Display/n1605 ),
    .i1(\u2_Display/n1612 [4]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1640 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3097  (
    .i0(\u2_Display/n1606 ),
    .i1(\u2_Display/n1612 [3]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1641 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3098  (
    .i0(\u2_Display/n1607 ),
    .i1(\u2_Display/n1612 [2]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1642 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3099  (
    .i0(\u2_Display/n1608 ),
    .i1(\u2_Display/n1612 [1]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1643 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3100  (
    .i0(\u2_Display/n1609 ),
    .i1(\u2_Display/n1612 [0]),
    .sel(\u2_Display/n1611 ),
    .o(\u2_Display/n1644 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3101  (\u2_Display/n1646 , \u2_Display/n1645 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3134  (
    .i0(\u2_Display/n1613 ),
    .i1(\u2_Display/n1647 [31]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1648 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3135  (
    .i0(\u2_Display/n1614 ),
    .i1(\u2_Display/n1647 [30]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1649 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3136  (
    .i0(\u2_Display/n1615 ),
    .i1(\u2_Display/n1647 [29]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1650 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3137  (
    .i0(\u2_Display/n1616 ),
    .i1(\u2_Display/n1647 [28]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1651 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3138  (
    .i0(\u2_Display/n1617 ),
    .i1(\u2_Display/n1647 [27]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1652 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3139  (
    .i0(\u2_Display/n1618 ),
    .i1(\u2_Display/n1647 [26]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1653 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3140  (
    .i0(\u2_Display/n1619 ),
    .i1(\u2_Display/n1647 [25]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1654 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3141  (
    .i0(\u2_Display/n1620 ),
    .i1(\u2_Display/n1647 [24]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1655 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3142  (
    .i0(\u2_Display/n1621 ),
    .i1(\u2_Display/n1647 [23]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1656 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3143  (
    .i0(\u2_Display/n1622 ),
    .i1(\u2_Display/n1647 [22]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1657 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3144  (
    .i0(\u2_Display/n1623 ),
    .i1(\u2_Display/n1647 [21]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1658 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3145  (
    .i0(\u2_Display/n1624 ),
    .i1(\u2_Display/n1647 [20]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1659 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3146  (
    .i0(\u2_Display/n1625 ),
    .i1(\u2_Display/n1647 [19]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1660 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3147  (
    .i0(\u2_Display/n1626 ),
    .i1(\u2_Display/n1647 [18]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1661 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3148  (
    .i0(\u2_Display/n1627 ),
    .i1(\u2_Display/n1647 [17]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1662 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3149  (
    .i0(\u2_Display/n1628 ),
    .i1(\u2_Display/n1647 [16]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1663 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3150  (
    .i0(\u2_Display/n1629 ),
    .i1(\u2_Display/n1647 [15]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1664 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3151  (
    .i0(\u2_Display/n1630 ),
    .i1(\u2_Display/n1647 [14]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1665 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3152  (
    .i0(\u2_Display/n1631 ),
    .i1(\u2_Display/n1647 [13]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1666 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3153  (
    .i0(\u2_Display/n1632 ),
    .i1(\u2_Display/n1647 [12]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1667 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3154  (
    .i0(\u2_Display/n1633 ),
    .i1(\u2_Display/n1647 [11]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1668 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3155  (
    .i0(\u2_Display/n1634 ),
    .i1(\u2_Display/n1647 [10]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1669 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3156  (
    .i0(\u2_Display/n1635 ),
    .i1(\u2_Display/n1647 [9]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1670 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3157  (
    .i0(\u2_Display/n1636 ),
    .i1(\u2_Display/n1647 [8]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1671 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3158  (
    .i0(\u2_Display/n1637 ),
    .i1(\u2_Display/n1647 [7]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1672 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3159  (
    .i0(\u2_Display/n1638 ),
    .i1(\u2_Display/n1647 [6]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1673 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3160  (
    .i0(\u2_Display/n1639 ),
    .i1(\u2_Display/n1647 [5]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1674 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3161  (
    .i0(\u2_Display/n1640 ),
    .i1(\u2_Display/n1647 [4]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1675 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3162  (
    .i0(\u2_Display/n1641 ),
    .i1(\u2_Display/n1647 [3]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1676 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3163  (
    .i0(\u2_Display/n1642 ),
    .i1(\u2_Display/n1647 [2]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1677 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3164  (
    .i0(\u2_Display/n1643 ),
    .i1(\u2_Display/n1647 [1]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1678 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3165  (
    .i0(\u2_Display/n1644 ),
    .i1(\u2_Display/n1647 [0]),
    .sel(\u2_Display/n1646 ),
    .o(\u2_Display/n1679 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3166  (\u2_Display/n1681 , \u2_Display/n1680 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3199  (
    .i0(\u2_Display/n1648 ),
    .i1(\u2_Display/n1682 [31]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1683 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3200  (
    .i0(\u2_Display/n1649 ),
    .i1(\u2_Display/n1682 [30]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1684 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3201  (
    .i0(\u2_Display/n1650 ),
    .i1(\u2_Display/n1682 [29]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1685 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3202  (
    .i0(\u2_Display/n1651 ),
    .i1(\u2_Display/n1682 [28]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1686 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3203  (
    .i0(\u2_Display/n1652 ),
    .i1(\u2_Display/n1682 [27]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1687 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3204  (
    .i0(\u2_Display/n1653 ),
    .i1(\u2_Display/n1682 [26]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1688 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3205  (
    .i0(\u2_Display/n1654 ),
    .i1(\u2_Display/n1682 [25]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1689 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3206  (
    .i0(\u2_Display/n1655 ),
    .i1(\u2_Display/n1682 [24]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1690 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3207  (
    .i0(\u2_Display/n1656 ),
    .i1(\u2_Display/n1682 [23]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1691 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3208  (
    .i0(\u2_Display/n1657 ),
    .i1(\u2_Display/n1682 [22]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1692 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3209  (
    .i0(\u2_Display/n1658 ),
    .i1(\u2_Display/n1682 [21]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1693 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3210  (
    .i0(\u2_Display/n1659 ),
    .i1(\u2_Display/n1682 [20]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1694 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3211  (
    .i0(\u2_Display/n1660 ),
    .i1(\u2_Display/n1682 [19]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1695 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3212  (
    .i0(\u2_Display/n1661 ),
    .i1(\u2_Display/n1682 [18]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1696 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3213  (
    .i0(\u2_Display/n1662 ),
    .i1(\u2_Display/n1682 [17]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1697 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3214  (
    .i0(\u2_Display/n1663 ),
    .i1(\u2_Display/n1682 [16]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1698 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3215  (
    .i0(\u2_Display/n1664 ),
    .i1(\u2_Display/n1682 [15]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1699 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3216  (
    .i0(\u2_Display/n1665 ),
    .i1(\u2_Display/n1682 [14]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1700 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3217  (
    .i0(\u2_Display/n1666 ),
    .i1(\u2_Display/n1682 [13]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1701 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3218  (
    .i0(\u2_Display/n1667 ),
    .i1(\u2_Display/n1682 [12]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1702 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3219  (
    .i0(\u2_Display/n1668 ),
    .i1(\u2_Display/n1682 [11]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1703 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3220  (
    .i0(\u2_Display/n1669 ),
    .i1(\u2_Display/n1682 [10]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1704 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3221  (
    .i0(\u2_Display/n1670 ),
    .i1(\u2_Display/n1682 [9]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1705 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3222  (
    .i0(\u2_Display/n1671 ),
    .i1(\u2_Display/n1682 [8]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1706 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3223  (
    .i0(\u2_Display/n1672 ),
    .i1(\u2_Display/n1682 [7]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1707 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3224  (
    .i0(\u2_Display/n1673 ),
    .i1(\u2_Display/n1682 [6]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1708 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3225  (
    .i0(\u2_Display/n1674 ),
    .i1(\u2_Display/n1682 [5]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1709 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3226  (
    .i0(\u2_Display/n1675 ),
    .i1(\u2_Display/n1682 [4]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1710 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3227  (
    .i0(\u2_Display/n1676 ),
    .i1(\u2_Display/n1682 [3]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1711 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3228  (
    .i0(\u2_Display/n1677 ),
    .i1(\u2_Display/n1682 [2]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1712 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3229  (
    .i0(\u2_Display/n1678 ),
    .i1(\u2_Display/n1682 [1]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1713 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3230  (
    .i0(\u2_Display/n1679 ),
    .i1(\u2_Display/n1682 [0]),
    .sel(\u2_Display/n1681 ),
    .o(\u2_Display/n1714 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3231  (\u2_Display/n1716 , \u2_Display/n1715 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3264  (
    .i0(\u2_Display/n1683 ),
    .i1(\u2_Display/n1717 [31]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1718 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3265  (
    .i0(\u2_Display/n1684 ),
    .i1(\u2_Display/n1717 [30]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1719 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3266  (
    .i0(\u2_Display/n1685 ),
    .i1(\u2_Display/n1717 [29]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1720 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3267  (
    .i0(\u2_Display/n1686 ),
    .i1(\u2_Display/n1717 [28]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1721 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3268  (
    .i0(\u2_Display/n1687 ),
    .i1(\u2_Display/n1717 [27]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1722 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3269  (
    .i0(\u2_Display/n1688 ),
    .i1(\u2_Display/n1717 [26]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1723 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3270  (
    .i0(\u2_Display/n1689 ),
    .i1(\u2_Display/n1717 [25]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1724 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3271  (
    .i0(\u2_Display/n1690 ),
    .i1(\u2_Display/n1717 [24]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1725 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3272  (
    .i0(\u2_Display/n1691 ),
    .i1(\u2_Display/n1717 [23]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1726 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3273  (
    .i0(\u2_Display/n1692 ),
    .i1(\u2_Display/n1717 [22]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1727 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3274  (
    .i0(\u2_Display/n1693 ),
    .i1(\u2_Display/n1717 [21]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1728 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3275  (
    .i0(\u2_Display/n1694 ),
    .i1(\u2_Display/n1717 [20]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1729 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3276  (
    .i0(\u2_Display/n1695 ),
    .i1(\u2_Display/n1717 [19]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1730 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3277  (
    .i0(\u2_Display/n1696 ),
    .i1(\u2_Display/n1717 [18]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1731 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3278  (
    .i0(\u2_Display/n1697 ),
    .i1(\u2_Display/n1717 [17]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1732 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3279  (
    .i0(\u2_Display/n1698 ),
    .i1(\u2_Display/n1717 [16]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1733 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3280  (
    .i0(\u2_Display/n1699 ),
    .i1(\u2_Display/n1717 [15]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1734 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3281  (
    .i0(\u2_Display/n1700 ),
    .i1(\u2_Display/n1717 [14]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1735 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3282  (
    .i0(\u2_Display/n1701 ),
    .i1(\u2_Display/n1717 [13]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1736 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3283  (
    .i0(\u2_Display/n1702 ),
    .i1(\u2_Display/n1717 [12]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1737 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3284  (
    .i0(\u2_Display/n1703 ),
    .i1(\u2_Display/n1717 [11]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1738 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3285  (
    .i0(\u2_Display/n1704 ),
    .i1(\u2_Display/n1717 [10]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1739 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3286  (
    .i0(\u2_Display/n1705 ),
    .i1(\u2_Display/n1717 [9]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1740 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3287  (
    .i0(\u2_Display/n1706 ),
    .i1(\u2_Display/n1717 [8]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1741 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3288  (
    .i0(\u2_Display/n1707 ),
    .i1(\u2_Display/n1717 [7]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1742 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3289  (
    .i0(\u2_Display/n1708 ),
    .i1(\u2_Display/n1717 [6]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1743 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3290  (
    .i0(\u2_Display/n1709 ),
    .i1(\u2_Display/n1717 [5]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1744 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3291  (
    .i0(\u2_Display/n1710 ),
    .i1(\u2_Display/n1717 [4]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1745 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3292  (
    .i0(\u2_Display/n1711 ),
    .i1(\u2_Display/n1717 [3]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1746 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3293  (
    .i0(\u2_Display/n1712 ),
    .i1(\u2_Display/n1717 [2]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1747 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3294  (
    .i0(\u2_Display/n1713 ),
    .i1(\u2_Display/n1717 [1]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1748 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3295  (
    .i0(\u2_Display/n1714 ),
    .i1(\u2_Display/n1717 [0]),
    .sel(\u2_Display/n1716 ),
    .o(\u2_Display/n1749 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3296  (\u2_Display/n1751 , \u2_Display/n1750 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3329  (
    .i0(\u2_Display/n1718 ),
    .i1(\u2_Display/n1752 [31]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1753 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3330  (
    .i0(\u2_Display/n1719 ),
    .i1(\u2_Display/n1752 [30]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1754 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3331  (
    .i0(\u2_Display/n1720 ),
    .i1(\u2_Display/n1752 [29]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1755 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3332  (
    .i0(\u2_Display/n1721 ),
    .i1(\u2_Display/n1752 [28]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1756 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3333  (
    .i0(\u2_Display/n1722 ),
    .i1(\u2_Display/n1752 [27]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1757 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3334  (
    .i0(\u2_Display/n1723 ),
    .i1(\u2_Display/n1752 [26]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1758 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3335  (
    .i0(\u2_Display/n1724 ),
    .i1(\u2_Display/n1752 [25]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1759 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3336  (
    .i0(\u2_Display/n1725 ),
    .i1(\u2_Display/n1752 [24]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1760 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3337  (
    .i0(\u2_Display/n1726 ),
    .i1(\u2_Display/n1752 [23]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1761 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3338  (
    .i0(\u2_Display/n1727 ),
    .i1(\u2_Display/n1752 [22]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1762 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3339  (
    .i0(\u2_Display/n1728 ),
    .i1(\u2_Display/n1752 [21]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1763 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3340  (
    .i0(\u2_Display/n1729 ),
    .i1(\u2_Display/n1752 [20]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1764 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3341  (
    .i0(\u2_Display/n1730 ),
    .i1(\u2_Display/n1752 [19]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1765 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3342  (
    .i0(\u2_Display/n1731 ),
    .i1(\u2_Display/n1752 [18]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1766 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3343  (
    .i0(\u2_Display/n1732 ),
    .i1(\u2_Display/n1752 [17]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1767 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3344  (
    .i0(\u2_Display/n1733 ),
    .i1(\u2_Display/n1752 [16]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1768 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3345  (
    .i0(\u2_Display/n1734 ),
    .i1(\u2_Display/n1752 [15]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1769 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3346  (
    .i0(\u2_Display/n1735 ),
    .i1(\u2_Display/n1752 [14]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1770 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3347  (
    .i0(\u2_Display/n1736 ),
    .i1(\u2_Display/n1752 [13]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1771 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3348  (
    .i0(\u2_Display/n1737 ),
    .i1(\u2_Display/n1752 [12]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1772 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3349  (
    .i0(\u2_Display/n1738 ),
    .i1(\u2_Display/n1752 [11]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1773 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3350  (
    .i0(\u2_Display/n1739 ),
    .i1(\u2_Display/n1752 [10]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1774 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3351  (
    .i0(\u2_Display/n1740 ),
    .i1(\u2_Display/n1752 [9]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1775 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3352  (
    .i0(\u2_Display/n1741 ),
    .i1(\u2_Display/n1752 [8]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1776 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3353  (
    .i0(\u2_Display/n1742 ),
    .i1(\u2_Display/n1752 [7]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1777 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3354  (
    .i0(\u2_Display/n1743 ),
    .i1(\u2_Display/n1752 [6]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1778 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3355  (
    .i0(\u2_Display/n1744 ),
    .i1(\u2_Display/n1752 [5]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1779 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3356  (
    .i0(\u2_Display/n1745 ),
    .i1(\u2_Display/n1752 [4]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1780 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3357  (
    .i0(\u2_Display/n1746 ),
    .i1(\u2_Display/n1752 [3]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1781 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3358  (
    .i0(\u2_Display/n1747 ),
    .i1(\u2_Display/n1752 [2]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1782 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3359  (
    .i0(\u2_Display/n1748 ),
    .i1(\u2_Display/n1752 [1]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1783 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3360  (
    .i0(\u2_Display/n1749 ),
    .i1(\u2_Display/n1752 [0]),
    .sel(\u2_Display/n1751 ),
    .o(\u2_Display/n1784 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3361  (\u2_Display/n1786 , \u2_Display/n1785 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3394  (
    .i0(\u2_Display/n1753 ),
    .i1(\u2_Display/n1787 [31]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1788 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3395  (
    .i0(\u2_Display/n1754 ),
    .i1(\u2_Display/n1787 [30]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1789 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3396  (
    .i0(\u2_Display/n1755 ),
    .i1(\u2_Display/n1787 [29]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1790 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3397  (
    .i0(\u2_Display/n1756 ),
    .i1(\u2_Display/n1787 [28]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1791 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3398  (
    .i0(\u2_Display/n1757 ),
    .i1(\u2_Display/n1787 [27]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1792 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3399  (
    .i0(\u2_Display/n1758 ),
    .i1(\u2_Display/n1787 [26]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1793 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3400  (
    .i0(\u2_Display/n1759 ),
    .i1(\u2_Display/n1787 [25]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1794 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3401  (
    .i0(\u2_Display/n1760 ),
    .i1(\u2_Display/n1787 [24]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1795 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3402  (
    .i0(\u2_Display/n1761 ),
    .i1(\u2_Display/n1787 [23]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1796 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3403  (
    .i0(\u2_Display/n1762 ),
    .i1(\u2_Display/n1787 [22]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1797 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3404  (
    .i0(\u2_Display/n1763 ),
    .i1(\u2_Display/n1787 [21]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1798 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3405  (
    .i0(\u2_Display/n1764 ),
    .i1(\u2_Display/n1787 [20]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1799 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3406  (
    .i0(\u2_Display/n1765 ),
    .i1(\u2_Display/n1787 [19]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1800 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3407  (
    .i0(\u2_Display/n1766 ),
    .i1(\u2_Display/n1787 [18]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1801 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3408  (
    .i0(\u2_Display/n1767 ),
    .i1(\u2_Display/n1787 [17]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1802 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3409  (
    .i0(\u2_Display/n1768 ),
    .i1(\u2_Display/n1787 [16]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1803 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3410  (
    .i0(\u2_Display/n1769 ),
    .i1(\u2_Display/n1787 [15]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1804 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3411  (
    .i0(\u2_Display/n1770 ),
    .i1(\u2_Display/n1787 [14]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1805 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3412  (
    .i0(\u2_Display/n1771 ),
    .i1(\u2_Display/n1787 [13]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1806 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3413  (
    .i0(\u2_Display/n1772 ),
    .i1(\u2_Display/n1787 [12]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1807 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3414  (
    .i0(\u2_Display/n1773 ),
    .i1(\u2_Display/n1787 [11]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1808 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3415  (
    .i0(\u2_Display/n1774 ),
    .i1(\u2_Display/n1787 [10]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1809 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3416  (
    .i0(\u2_Display/n1775 ),
    .i1(\u2_Display/n1787 [9]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1810 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3417  (
    .i0(\u2_Display/n1776 ),
    .i1(\u2_Display/n1787 [8]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1811 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3418  (
    .i0(\u2_Display/n1777 ),
    .i1(\u2_Display/n1787 [7]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1812 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3419  (
    .i0(\u2_Display/n1778 ),
    .i1(\u2_Display/n1787 [6]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1813 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3420  (
    .i0(\u2_Display/n1779 ),
    .i1(\u2_Display/n1787 [5]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1814 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3421  (
    .i0(\u2_Display/n1780 ),
    .i1(\u2_Display/n1787 [4]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1815 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3422  (
    .i0(\u2_Display/n1781 ),
    .i1(\u2_Display/n1787 [3]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1816 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3423  (
    .i0(\u2_Display/n1782 ),
    .i1(\u2_Display/n1787 [2]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1817 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3424  (
    .i0(\u2_Display/n1783 ),
    .i1(\u2_Display/n1787 [1]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1818 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3425  (
    .i0(\u2_Display/n1784 ),
    .i1(\u2_Display/n1787 [0]),
    .sel(\u2_Display/n1786 ),
    .o(\u2_Display/n1819 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3426  (\u2_Display/n1821 , \u2_Display/n1820 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3459  (
    .i0(\u2_Display/n1788 ),
    .i1(\u2_Display/n1822 [31]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1823 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3460  (
    .i0(\u2_Display/n1789 ),
    .i1(\u2_Display/n1822 [30]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1824 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3461  (
    .i0(\u2_Display/n1790 ),
    .i1(\u2_Display/n1822 [29]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1825 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3462  (
    .i0(\u2_Display/n1791 ),
    .i1(\u2_Display/n1822 [28]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1826 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3463  (
    .i0(\u2_Display/n1792 ),
    .i1(\u2_Display/n1822 [27]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1827 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3464  (
    .i0(\u2_Display/n1793 ),
    .i1(\u2_Display/n1822 [26]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1828 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3465  (
    .i0(\u2_Display/n1794 ),
    .i1(\u2_Display/n1822 [25]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1829 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3466  (
    .i0(\u2_Display/n1795 ),
    .i1(\u2_Display/n1822 [24]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1830 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3467  (
    .i0(\u2_Display/n1796 ),
    .i1(\u2_Display/n1822 [23]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1831 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3468  (
    .i0(\u2_Display/n1797 ),
    .i1(\u2_Display/n1822 [22]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1832 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3469  (
    .i0(\u2_Display/n1798 ),
    .i1(\u2_Display/n1822 [21]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1833 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3470  (
    .i0(\u2_Display/n1799 ),
    .i1(\u2_Display/n1822 [20]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1834 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3471  (
    .i0(\u2_Display/n1800 ),
    .i1(\u2_Display/n1822 [19]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1835 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3472  (
    .i0(\u2_Display/n1801 ),
    .i1(\u2_Display/n1822 [18]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1836 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3473  (
    .i0(\u2_Display/n1802 ),
    .i1(\u2_Display/n1822 [17]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1837 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3474  (
    .i0(\u2_Display/n1803 ),
    .i1(\u2_Display/n1822 [16]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1838 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3475  (
    .i0(\u2_Display/n1804 ),
    .i1(\u2_Display/n1822 [15]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1839 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3476  (
    .i0(\u2_Display/n1805 ),
    .i1(\u2_Display/n1822 [14]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1840 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3477  (
    .i0(\u2_Display/n1806 ),
    .i1(\u2_Display/n1822 [13]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1841 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3478  (
    .i0(\u2_Display/n1807 ),
    .i1(\u2_Display/n1822 [12]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1842 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3479  (
    .i0(\u2_Display/n1808 ),
    .i1(\u2_Display/n1822 [11]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1843 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3480  (
    .i0(\u2_Display/n1809 ),
    .i1(\u2_Display/n1822 [10]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1844 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3481  (
    .i0(\u2_Display/n1810 ),
    .i1(\u2_Display/n1822 [9]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1845 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3482  (
    .i0(\u2_Display/n1811 ),
    .i1(\u2_Display/n1822 [8]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1846 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3483  (
    .i0(\u2_Display/n1812 ),
    .i1(\u2_Display/n1822 [7]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1847 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3484  (
    .i0(\u2_Display/n1813 ),
    .i1(\u2_Display/n1822 [6]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1848 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3485  (
    .i0(\u2_Display/n1814 ),
    .i1(\u2_Display/n1822 [5]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1849 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3486  (
    .i0(\u2_Display/n1815 ),
    .i1(\u2_Display/n1822 [4]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1850 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3487  (
    .i0(\u2_Display/n1816 ),
    .i1(\u2_Display/n1822 [3]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1851 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3488  (
    .i0(\u2_Display/n1817 ),
    .i1(\u2_Display/n1822 [2]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1852 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3489  (
    .i0(\u2_Display/n1818 ),
    .i1(\u2_Display/n1822 [1]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1853 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3490  (
    .i0(\u2_Display/n1819 ),
    .i1(\u2_Display/n1822 [0]),
    .sel(\u2_Display/n1821 ),
    .o(\u2_Display/n1854 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3491  (\u2_Display/n1856 , \u2_Display/n1855 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3524  (
    .i0(\u2_Display/n1823 ),
    .i1(\u2_Display/n1857 [31]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1858 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3525  (
    .i0(\u2_Display/n1824 ),
    .i1(\u2_Display/n1857 [30]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1859 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3526  (
    .i0(\u2_Display/n1825 ),
    .i1(\u2_Display/n1857 [29]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1860 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3527  (
    .i0(\u2_Display/n1826 ),
    .i1(\u2_Display/n1857 [28]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1861 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3528  (
    .i0(\u2_Display/n1827 ),
    .i1(\u2_Display/n1857 [27]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1862 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3529  (
    .i0(\u2_Display/n1828 ),
    .i1(\u2_Display/n1857 [26]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1863 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3530  (
    .i0(\u2_Display/n1829 ),
    .i1(\u2_Display/n1857 [25]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1864 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3531  (
    .i0(\u2_Display/n1830 ),
    .i1(\u2_Display/n1857 [24]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1865 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3532  (
    .i0(\u2_Display/n1831 ),
    .i1(\u2_Display/n1857 [23]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1866 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3533  (
    .i0(\u2_Display/n1832 ),
    .i1(\u2_Display/n1857 [22]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1867 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3534  (
    .i0(\u2_Display/n1833 ),
    .i1(\u2_Display/n1857 [21]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1868 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3535  (
    .i0(\u2_Display/n1834 ),
    .i1(\u2_Display/n1857 [20]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1869 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3536  (
    .i0(\u2_Display/n1835 ),
    .i1(\u2_Display/n1857 [19]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1870 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3537  (
    .i0(\u2_Display/n1836 ),
    .i1(\u2_Display/n1857 [18]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1871 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3538  (
    .i0(\u2_Display/n1837 ),
    .i1(\u2_Display/n1857 [17]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1872 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3539  (
    .i0(\u2_Display/n1838 ),
    .i1(\u2_Display/n1857 [16]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1873 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3540  (
    .i0(\u2_Display/n1839 ),
    .i1(\u2_Display/n1857 [15]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1874 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3541  (
    .i0(\u2_Display/n1840 ),
    .i1(\u2_Display/n1857 [14]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1875 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3542  (
    .i0(\u2_Display/n1841 ),
    .i1(\u2_Display/n1857 [13]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1876 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3543  (
    .i0(\u2_Display/n1842 ),
    .i1(\u2_Display/n1857 [12]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1877 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3544  (
    .i0(\u2_Display/n1843 ),
    .i1(\u2_Display/n1857 [11]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1878 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3545  (
    .i0(\u2_Display/n1844 ),
    .i1(\u2_Display/n1857 [10]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1879 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3546  (
    .i0(\u2_Display/n1845 ),
    .i1(\u2_Display/n1857 [9]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1880 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3547  (
    .i0(\u2_Display/n1846 ),
    .i1(\u2_Display/n1857 [8]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1881 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3548  (
    .i0(\u2_Display/n1847 ),
    .i1(\u2_Display/n1857 [7]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1882 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3549  (
    .i0(\u2_Display/n1848 ),
    .i1(\u2_Display/n1857 [6]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1883 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3550  (
    .i0(\u2_Display/n1849 ),
    .i1(\u2_Display/n1857 [5]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1884 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3551  (
    .i0(\u2_Display/n1850 ),
    .i1(\u2_Display/n1857 [4]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1885 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3552  (
    .i0(\u2_Display/n1851 ),
    .i1(\u2_Display/n1857 [3]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1886 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3553  (
    .i0(\u2_Display/n1852 ),
    .i1(\u2_Display/n1857 [2]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1887 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3554  (
    .i0(\u2_Display/n1853 ),
    .i1(\u2_Display/n1857 [1]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1888 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3555  (
    .i0(\u2_Display/n1854 ),
    .i1(\u2_Display/n1857 [0]),
    .sel(\u2_Display/n1856 ),
    .o(\u2_Display/n1889 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3556  (\u2_Display/n1891 , \u2_Display/n1890 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3589  (
    .i0(\u2_Display/n1858 ),
    .i1(\u2_Display/n1892 [31]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1893 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3590  (
    .i0(\u2_Display/n1859 ),
    .i1(\u2_Display/n1892 [30]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1894 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3591  (
    .i0(\u2_Display/n1860 ),
    .i1(\u2_Display/n1892 [29]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1895 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3592  (
    .i0(\u2_Display/n1861 ),
    .i1(\u2_Display/n1892 [28]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1896 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3593  (
    .i0(\u2_Display/n1862 ),
    .i1(\u2_Display/n1892 [27]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1897 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3594  (
    .i0(\u2_Display/n1863 ),
    .i1(\u2_Display/n1892 [26]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1898 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3595  (
    .i0(\u2_Display/n1864 ),
    .i1(\u2_Display/n1892 [25]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1899 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3596  (
    .i0(\u2_Display/n1865 ),
    .i1(\u2_Display/n1892 [24]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1900 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3597  (
    .i0(\u2_Display/n1866 ),
    .i1(\u2_Display/n1892 [23]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1901 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3598  (
    .i0(\u2_Display/n1867 ),
    .i1(\u2_Display/n1892 [22]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1902 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3599  (
    .i0(\u2_Display/n1868 ),
    .i1(\u2_Display/n1892 [21]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1903 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3600  (
    .i0(\u2_Display/n1869 ),
    .i1(\u2_Display/n1892 [20]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1904 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3601  (
    .i0(\u2_Display/n1870 ),
    .i1(\u2_Display/n1892 [19]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1905 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3602  (
    .i0(\u2_Display/n1871 ),
    .i1(\u2_Display/n1892 [18]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1906 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3603  (
    .i0(\u2_Display/n1872 ),
    .i1(\u2_Display/n1892 [17]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1907 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3604  (
    .i0(\u2_Display/n1873 ),
    .i1(\u2_Display/n1892 [16]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1908 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3605  (
    .i0(\u2_Display/n1874 ),
    .i1(\u2_Display/n1892 [15]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1909 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3606  (
    .i0(\u2_Display/n1875 ),
    .i1(\u2_Display/n1892 [14]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1910 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3607  (
    .i0(\u2_Display/n1876 ),
    .i1(\u2_Display/n1892 [13]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1911 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3608  (
    .i0(\u2_Display/n1877 ),
    .i1(\u2_Display/n1892 [12]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1912 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3609  (
    .i0(\u2_Display/n1878 ),
    .i1(\u2_Display/n1892 [11]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1913 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3610  (
    .i0(\u2_Display/n1879 ),
    .i1(\u2_Display/n1892 [10]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1914 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3611  (
    .i0(\u2_Display/n1880 ),
    .i1(\u2_Display/n1892 [9]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1915 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3612  (
    .i0(\u2_Display/n1881 ),
    .i1(\u2_Display/n1892 [8]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1916 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3613  (
    .i0(\u2_Display/n1882 ),
    .i1(\u2_Display/n1892 [7]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1917 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3614  (
    .i0(\u2_Display/n1883 ),
    .i1(\u2_Display/n1892 [6]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1918 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3615  (
    .i0(\u2_Display/n1884 ),
    .i1(\u2_Display/n1892 [5]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1919 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3616  (
    .i0(\u2_Display/n1885 ),
    .i1(\u2_Display/n1892 [4]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1920 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3617  (
    .i0(\u2_Display/n1886 ),
    .i1(\u2_Display/n1892 [3]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1921 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3618  (
    .i0(\u2_Display/n1887 ),
    .i1(\u2_Display/n1892 [2]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1922 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3619  (
    .i0(\u2_Display/n1888 ),
    .i1(\u2_Display/n1892 [1]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1923 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3620  (
    .i0(\u2_Display/n1889 ),
    .i1(\u2_Display/n1892 [0]),
    .sel(\u2_Display/n1891 ),
    .o(\u2_Display/n1924 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3621  (\u2_Display/n1926 , \u2_Display/n1925 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3654  (
    .i0(\u2_Display/n1893 ),
    .i1(\u2_Display/n1927 [31]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1928 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3655  (
    .i0(\u2_Display/n1894 ),
    .i1(\u2_Display/n1927 [30]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1929 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3656  (
    .i0(\u2_Display/n1895 ),
    .i1(\u2_Display/n1927 [29]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1930 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3657  (
    .i0(\u2_Display/n1896 ),
    .i1(\u2_Display/n1927 [28]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1931 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3658  (
    .i0(\u2_Display/n1897 ),
    .i1(\u2_Display/n1927 [27]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1932 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3659  (
    .i0(\u2_Display/n1898 ),
    .i1(\u2_Display/n1927 [26]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1933 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3660  (
    .i0(\u2_Display/n1899 ),
    .i1(\u2_Display/n1927 [25]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1934 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3661  (
    .i0(\u2_Display/n1900 ),
    .i1(\u2_Display/n1927 [24]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1935 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3662  (
    .i0(\u2_Display/n1901 ),
    .i1(\u2_Display/n1927 [23]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1936 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3663  (
    .i0(\u2_Display/n1902 ),
    .i1(\u2_Display/n1927 [22]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1937 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3664  (
    .i0(\u2_Display/n1903 ),
    .i1(\u2_Display/n1927 [21]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1938 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3665  (
    .i0(\u2_Display/n1904 ),
    .i1(\u2_Display/n1927 [20]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1939 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3666  (
    .i0(\u2_Display/n1905 ),
    .i1(\u2_Display/n1927 [19]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1940 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3667  (
    .i0(\u2_Display/n1906 ),
    .i1(\u2_Display/n1927 [18]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1941 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3668  (
    .i0(\u2_Display/n1907 ),
    .i1(\u2_Display/n1927 [17]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1942 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3669  (
    .i0(\u2_Display/n1908 ),
    .i1(\u2_Display/n1927 [16]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1943 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3670  (
    .i0(\u2_Display/n1909 ),
    .i1(\u2_Display/n1927 [15]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1944 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3671  (
    .i0(\u2_Display/n1910 ),
    .i1(\u2_Display/n1927 [14]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1945 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3672  (
    .i0(\u2_Display/n1911 ),
    .i1(\u2_Display/n1927 [13]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1946 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3673  (
    .i0(\u2_Display/n1912 ),
    .i1(\u2_Display/n1927 [12]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1947 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3674  (
    .i0(\u2_Display/n1913 ),
    .i1(\u2_Display/n1927 [11]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1948 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3675  (
    .i0(\u2_Display/n1914 ),
    .i1(\u2_Display/n1927 [10]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1949 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3676  (
    .i0(\u2_Display/n1915 ),
    .i1(\u2_Display/n1927 [9]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1950 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3677  (
    .i0(\u2_Display/n1916 ),
    .i1(\u2_Display/n1927 [8]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1951 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3678  (
    .i0(\u2_Display/n1917 ),
    .i1(\u2_Display/n1927 [7]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1952 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3679  (
    .i0(\u2_Display/n1918 ),
    .i1(\u2_Display/n1927 [6]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1953 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3680  (
    .i0(\u2_Display/n1919 ),
    .i1(\u2_Display/n1927 [5]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1954 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3681  (
    .i0(\u2_Display/n1920 ),
    .i1(\u2_Display/n1927 [4]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1955 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3682  (
    .i0(\u2_Display/n1921 ),
    .i1(\u2_Display/n1927 [3]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1956 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3683  (
    .i0(\u2_Display/n1922 ),
    .i1(\u2_Display/n1927 [2]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1957 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3684  (
    .i0(\u2_Display/n1923 ),
    .i1(\u2_Display/n1927 [1]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1958 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3685  (
    .i0(\u2_Display/n1924 ),
    .i1(\u2_Display/n1927 [0]),
    .sel(\u2_Display/n1926 ),
    .o(\u2_Display/n1959 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3686  (\u2_Display/n1961 , \u2_Display/n1960 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3719  (
    .i0(\u2_Display/n1928 ),
    .i1(\u2_Display/n1962 [31]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1963 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3720  (
    .i0(\u2_Display/n1929 ),
    .i1(\u2_Display/n1962 [30]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1964 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3721  (
    .i0(\u2_Display/n1930 ),
    .i1(\u2_Display/n1962 [29]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1965 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3722  (
    .i0(\u2_Display/n1931 ),
    .i1(\u2_Display/n1962 [28]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1966 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3723  (
    .i0(\u2_Display/n1932 ),
    .i1(\u2_Display/n1962 [27]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1967 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3724  (
    .i0(\u2_Display/n1933 ),
    .i1(\u2_Display/n1962 [26]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1968 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3725  (
    .i0(\u2_Display/n1934 ),
    .i1(\u2_Display/n1962 [25]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1969 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3726  (
    .i0(\u2_Display/n1935 ),
    .i1(\u2_Display/n1962 [24]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1970 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3727  (
    .i0(\u2_Display/n1936 ),
    .i1(\u2_Display/n1962 [23]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1971 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3728  (
    .i0(\u2_Display/n1937 ),
    .i1(\u2_Display/n1962 [22]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1972 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3729  (
    .i0(\u2_Display/n1938 ),
    .i1(\u2_Display/n1962 [21]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1973 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3730  (
    .i0(\u2_Display/n1939 ),
    .i1(\u2_Display/n1962 [20]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1974 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3731  (
    .i0(\u2_Display/n1940 ),
    .i1(\u2_Display/n1962 [19]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1975 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3732  (
    .i0(\u2_Display/n1941 ),
    .i1(\u2_Display/n1962 [18]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1976 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3733  (
    .i0(\u2_Display/n1942 ),
    .i1(\u2_Display/n1962 [17]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1977 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3734  (
    .i0(\u2_Display/n1943 ),
    .i1(\u2_Display/n1962 [16]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1978 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3735  (
    .i0(\u2_Display/n1944 ),
    .i1(\u2_Display/n1962 [15]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1979 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3736  (
    .i0(\u2_Display/n1945 ),
    .i1(\u2_Display/n1962 [14]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1980 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3737  (
    .i0(\u2_Display/n1946 ),
    .i1(\u2_Display/n1962 [13]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1981 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3738  (
    .i0(\u2_Display/n1947 ),
    .i1(\u2_Display/n1962 [12]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1982 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3739  (
    .i0(\u2_Display/n1948 ),
    .i1(\u2_Display/n1962 [11]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1983 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3740  (
    .i0(\u2_Display/n1949 ),
    .i1(\u2_Display/n1962 [10]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1984 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3741  (
    .i0(\u2_Display/n1950 ),
    .i1(\u2_Display/n1962 [9]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1985 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3742  (
    .i0(\u2_Display/n1951 ),
    .i1(\u2_Display/n1962 [8]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1986 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3743  (
    .i0(\u2_Display/n1952 ),
    .i1(\u2_Display/n1962 [7]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1987 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3744  (
    .i0(\u2_Display/n1953 ),
    .i1(\u2_Display/n1962 [6]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1988 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3745  (
    .i0(\u2_Display/n1954 ),
    .i1(\u2_Display/n1962 [5]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1989 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3746  (
    .i0(\u2_Display/n1955 ),
    .i1(\u2_Display/n1962 [4]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1990 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3747  (
    .i0(\u2_Display/n1956 ),
    .i1(\u2_Display/n1962 [3]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1991 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3748  (
    .i0(\u2_Display/n1957 ),
    .i1(\u2_Display/n1962 [2]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1992 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3749  (
    .i0(\u2_Display/n1958 ),
    .i1(\u2_Display/n1962 [1]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1993 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3750  (
    .i0(\u2_Display/n1959 ),
    .i1(\u2_Display/n1962 [0]),
    .sel(\u2_Display/n1961 ),
    .o(\u2_Display/n1994 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3751  (\u2_Display/n1996 , \u2_Display/n1995 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3784  (
    .i0(\u2_Display/n1963 ),
    .i1(\u2_Display/n1997 [31]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n1998 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3785  (
    .i0(\u2_Display/n1964 ),
    .i1(\u2_Display/n1997 [30]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n1999 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3786  (
    .i0(\u2_Display/n1965 ),
    .i1(\u2_Display/n1997 [29]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2000 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3787  (
    .i0(\u2_Display/n1966 ),
    .i1(\u2_Display/n1997 [28]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2001 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3788  (
    .i0(\u2_Display/n1967 ),
    .i1(\u2_Display/n1997 [27]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2002 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3789  (
    .i0(\u2_Display/n1968 ),
    .i1(\u2_Display/n1997 [26]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2003 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3790  (
    .i0(\u2_Display/n1969 ),
    .i1(\u2_Display/n1997 [25]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2004 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3791  (
    .i0(\u2_Display/n1970 ),
    .i1(\u2_Display/n1997 [24]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2005 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3792  (
    .i0(\u2_Display/n1971 ),
    .i1(\u2_Display/n1997 [23]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2006 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3793  (
    .i0(\u2_Display/n1972 ),
    .i1(\u2_Display/n1997 [22]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2007 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3794  (
    .i0(\u2_Display/n1973 ),
    .i1(\u2_Display/n1997 [21]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2008 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3795  (
    .i0(\u2_Display/n1974 ),
    .i1(\u2_Display/n1997 [20]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2009 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3796  (
    .i0(\u2_Display/n1975 ),
    .i1(\u2_Display/n1997 [19]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2010 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3797  (
    .i0(\u2_Display/n1976 ),
    .i1(\u2_Display/n1997 [18]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2011 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3798  (
    .i0(\u2_Display/n1977 ),
    .i1(\u2_Display/n1997 [17]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2012 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3799  (
    .i0(\u2_Display/n1978 ),
    .i1(\u2_Display/n1997 [16]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2013 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3800  (
    .i0(\u2_Display/n1979 ),
    .i1(\u2_Display/n1997 [15]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2014 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3801  (
    .i0(\u2_Display/n1980 ),
    .i1(\u2_Display/n1997 [14]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2015 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3802  (
    .i0(\u2_Display/n1981 ),
    .i1(\u2_Display/n1997 [13]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2016 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3803  (
    .i0(\u2_Display/n1982 ),
    .i1(\u2_Display/n1997 [12]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2017 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3804  (
    .i0(\u2_Display/n1983 ),
    .i1(\u2_Display/n1997 [11]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2018 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3805  (
    .i0(\u2_Display/n1984 ),
    .i1(\u2_Display/n1997 [10]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2019 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3806  (
    .i0(\u2_Display/n1985 ),
    .i1(\u2_Display/n1997 [9]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2020 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3807  (
    .i0(\u2_Display/n1986 ),
    .i1(\u2_Display/n1997 [8]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2021 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3808  (
    .i0(\u2_Display/n1987 ),
    .i1(\u2_Display/n1997 [7]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2022 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3809  (
    .i0(\u2_Display/n1988 ),
    .i1(\u2_Display/n1997 [6]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2023 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3810  (
    .i0(\u2_Display/n1989 ),
    .i1(\u2_Display/n1997 [5]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2024 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3811  (
    .i0(\u2_Display/n1990 ),
    .i1(\u2_Display/n1997 [4]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2025 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3812  (
    .i0(\u2_Display/n1991 ),
    .i1(\u2_Display/n1997 [3]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2026 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3813  (
    .i0(\u2_Display/n1992 ),
    .i1(\u2_Display/n1997 [2]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2027 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3814  (
    .i0(\u2_Display/n1993 ),
    .i1(\u2_Display/n1997 [1]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2028 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3815  (
    .i0(\u2_Display/n1994 ),
    .i1(\u2_Display/n1997 [0]),
    .sel(\u2_Display/n1996 ),
    .o(\u2_Display/n2029 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3816  (\u2_Display/n2031 , \u2_Display/n2030 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3849  (
    .i0(\u2_Display/n1998 ),
    .i1(\u2_Display/n2032 [31]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2033 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3850  (
    .i0(\u2_Display/n1999 ),
    .i1(\u2_Display/n2032 [30]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2034 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3851  (
    .i0(\u2_Display/n2000 ),
    .i1(\u2_Display/n2032 [29]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2035 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3852  (
    .i0(\u2_Display/n2001 ),
    .i1(\u2_Display/n2032 [28]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2036 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3853  (
    .i0(\u2_Display/n2002 ),
    .i1(\u2_Display/n2032 [27]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2037 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3854  (
    .i0(\u2_Display/n2003 ),
    .i1(\u2_Display/n2032 [26]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2038 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3855  (
    .i0(\u2_Display/n2004 ),
    .i1(\u2_Display/n2032 [25]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2039 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3856  (
    .i0(\u2_Display/n2005 ),
    .i1(\u2_Display/n2032 [24]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2040 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3857  (
    .i0(\u2_Display/n2006 ),
    .i1(\u2_Display/n2032 [23]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2041 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3858  (
    .i0(\u2_Display/n2007 ),
    .i1(\u2_Display/n2032 [22]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2042 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3859  (
    .i0(\u2_Display/n2008 ),
    .i1(\u2_Display/n2032 [21]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2043 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3860  (
    .i0(\u2_Display/n2009 ),
    .i1(\u2_Display/n2032 [20]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2044 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3861  (
    .i0(\u2_Display/n2010 ),
    .i1(\u2_Display/n2032 [19]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2045 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3862  (
    .i0(\u2_Display/n2011 ),
    .i1(\u2_Display/n2032 [18]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2046 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3863  (
    .i0(\u2_Display/n2012 ),
    .i1(\u2_Display/n2032 [17]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2047 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3864  (
    .i0(\u2_Display/n2013 ),
    .i1(\u2_Display/n2032 [16]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2048 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3865  (
    .i0(\u2_Display/n2014 ),
    .i1(\u2_Display/n2032 [15]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2049 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3866  (
    .i0(\u2_Display/n2015 ),
    .i1(\u2_Display/n2032 [14]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2050 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3867  (
    .i0(\u2_Display/n2016 ),
    .i1(\u2_Display/n2032 [13]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2051 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3868  (
    .i0(\u2_Display/n2017 ),
    .i1(\u2_Display/n2032 [12]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2052 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3869  (
    .i0(\u2_Display/n2018 ),
    .i1(\u2_Display/n2032 [11]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2053 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3870  (
    .i0(\u2_Display/n2019 ),
    .i1(\u2_Display/n2032 [10]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2054 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3871  (
    .i0(\u2_Display/n2020 ),
    .i1(\u2_Display/n2032 [9]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2055 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3872  (
    .i0(\u2_Display/n2021 ),
    .i1(\u2_Display/n2032 [8]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2056 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3873  (
    .i0(\u2_Display/n2022 ),
    .i1(\u2_Display/n2032 [7]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2057 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3874  (
    .i0(\u2_Display/n2023 ),
    .i1(\u2_Display/n2032 [6]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2058 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3875  (
    .i0(\u2_Display/n2024 ),
    .i1(\u2_Display/n2032 [5]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2059 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3876  (
    .i0(\u2_Display/n2025 ),
    .i1(\u2_Display/n2032 [4]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2060 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3877  (
    .i0(\u2_Display/n2026 ),
    .i1(\u2_Display/n2032 [3]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2061 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3878  (
    .i0(\u2_Display/n2027 ),
    .i1(\u2_Display/n2032 [2]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2062 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3879  (
    .i0(\u2_Display/n2028 ),
    .i1(\u2_Display/n2032 [1]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2063 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3880  (
    .i0(\u2_Display/n2029 ),
    .i1(\u2_Display/n2032 [0]),
    .sel(\u2_Display/n2031 ),
    .o(\u2_Display/n2064 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3881  (\u2_Display/n2066 , \u2_Display/n2065 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3914  (
    .i0(\u2_Display/n2033 ),
    .i1(\u2_Display/n2067 [31]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2068 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3915  (
    .i0(\u2_Display/n2034 ),
    .i1(\u2_Display/n2067 [30]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2069 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3916  (
    .i0(\u2_Display/n2035 ),
    .i1(\u2_Display/n2067 [29]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2070 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3917  (
    .i0(\u2_Display/n2036 ),
    .i1(\u2_Display/n2067 [28]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2071 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3918  (
    .i0(\u2_Display/n2037 ),
    .i1(\u2_Display/n2067 [27]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2072 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3919  (
    .i0(\u2_Display/n2038 ),
    .i1(\u2_Display/n2067 [26]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2073 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3920  (
    .i0(\u2_Display/n2039 ),
    .i1(\u2_Display/n2067 [25]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2074 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3921  (
    .i0(\u2_Display/n2040 ),
    .i1(\u2_Display/n2067 [24]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2075 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3922  (
    .i0(\u2_Display/n2041 ),
    .i1(\u2_Display/n2067 [23]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2076 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3923  (
    .i0(\u2_Display/n2042 ),
    .i1(\u2_Display/n2067 [22]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2077 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3924  (
    .i0(\u2_Display/n2043 ),
    .i1(\u2_Display/n2067 [21]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2078 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3925  (
    .i0(\u2_Display/n2044 ),
    .i1(\u2_Display/n2067 [20]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2079 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3926  (
    .i0(\u2_Display/n2045 ),
    .i1(\u2_Display/n2067 [19]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2080 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3927  (
    .i0(\u2_Display/n2046 ),
    .i1(\u2_Display/n2067 [18]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2081 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3928  (
    .i0(\u2_Display/n2047 ),
    .i1(\u2_Display/n2067 [17]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2082 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3929  (
    .i0(\u2_Display/n2048 ),
    .i1(\u2_Display/n2067 [16]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2083 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3930  (
    .i0(\u2_Display/n2049 ),
    .i1(\u2_Display/n2067 [15]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2084 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3931  (
    .i0(\u2_Display/n2050 ),
    .i1(\u2_Display/n2067 [14]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2085 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3932  (
    .i0(\u2_Display/n2051 ),
    .i1(\u2_Display/n2067 [13]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2086 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3933  (
    .i0(\u2_Display/n2052 ),
    .i1(\u2_Display/n2067 [12]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2087 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3934  (
    .i0(\u2_Display/n2053 ),
    .i1(\u2_Display/n2067 [11]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2088 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3935  (
    .i0(\u2_Display/n2054 ),
    .i1(\u2_Display/n2067 [10]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2089 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3936  (
    .i0(\u2_Display/n2055 ),
    .i1(\u2_Display/n2067 [9]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2090 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3937  (
    .i0(\u2_Display/n2056 ),
    .i1(\u2_Display/n2067 [8]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2091 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3938  (
    .i0(\u2_Display/n2057 ),
    .i1(\u2_Display/n2067 [7]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2092 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3939  (
    .i0(\u2_Display/n2058 ),
    .i1(\u2_Display/n2067 [6]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2093 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3940  (
    .i0(\u2_Display/n2059 ),
    .i1(\u2_Display/n2067 [5]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2094 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3941  (
    .i0(\u2_Display/n2060 ),
    .i1(\u2_Display/n2067 [4]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2095 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3942  (
    .i0(\u2_Display/n2061 ),
    .i1(\u2_Display/n2067 [3]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2096 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3943  (
    .i0(\u2_Display/n2062 ),
    .i1(\u2_Display/n2067 [2]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2097 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3944  (
    .i0(\u2_Display/n2063 ),
    .i1(\u2_Display/n2067 [1]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2098 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3945  (
    .i0(\u2_Display/n2064 ),
    .i1(\u2_Display/n2067 [0]),
    .sel(\u2_Display/n2066 ),
    .o(\u2_Display/n2099 ));  // source/rtl/Display.v(213)
  not \u2_Display/u3946  (\u2_Display/n2101 , \u2_Display/n2100 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3979  (
    .i0(\u2_Display/n2068 ),
    .i1(\u2_Display/n2102 [31]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2103 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3980  (
    .i0(\u2_Display/n2069 ),
    .i1(\u2_Display/n2102 [30]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2104 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3981  (
    .i0(\u2_Display/n2070 ),
    .i1(\u2_Display/n2102 [29]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2105 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3982  (
    .i0(\u2_Display/n2071 ),
    .i1(\u2_Display/n2102 [28]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2106 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3983  (
    .i0(\u2_Display/n2072 ),
    .i1(\u2_Display/n2102 [27]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2107 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3984  (
    .i0(\u2_Display/n2073 ),
    .i1(\u2_Display/n2102 [26]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2108 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3985  (
    .i0(\u2_Display/n2074 ),
    .i1(\u2_Display/n2102 [25]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2109 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3986  (
    .i0(\u2_Display/n2075 ),
    .i1(\u2_Display/n2102 [24]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2110 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3987  (
    .i0(\u2_Display/n2076 ),
    .i1(\u2_Display/n2102 [23]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2111 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3988  (
    .i0(\u2_Display/n2077 ),
    .i1(\u2_Display/n2102 [22]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2112 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3989  (
    .i0(\u2_Display/n2078 ),
    .i1(\u2_Display/n2102 [21]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2113 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3990  (
    .i0(\u2_Display/n2079 ),
    .i1(\u2_Display/n2102 [20]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2114 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3991  (
    .i0(\u2_Display/n2080 ),
    .i1(\u2_Display/n2102 [19]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2115 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3992  (
    .i0(\u2_Display/n2081 ),
    .i1(\u2_Display/n2102 [18]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2116 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3993  (
    .i0(\u2_Display/n2082 ),
    .i1(\u2_Display/n2102 [17]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2117 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3994  (
    .i0(\u2_Display/n2083 ),
    .i1(\u2_Display/n2102 [16]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2118 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3995  (
    .i0(\u2_Display/n2084 ),
    .i1(\u2_Display/n2102 [15]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2119 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3996  (
    .i0(\u2_Display/n2085 ),
    .i1(\u2_Display/n2102 [14]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2120 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3997  (
    .i0(\u2_Display/n2086 ),
    .i1(\u2_Display/n2102 [13]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2121 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3998  (
    .i0(\u2_Display/n2087 ),
    .i1(\u2_Display/n2102 [12]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2122 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u3999  (
    .i0(\u2_Display/n2088 ),
    .i1(\u2_Display/n2102 [11]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2123 ));  // source/rtl/Display.v(213)
  not \u2_Display/u4  (\u2_Display/n36 , \u2_Display/clk1s );  // source/rtl/Display.v(54)
  AL_MUX \u2_Display/u4000  (
    .i0(\u2_Display/n2089 ),
    .i1(\u2_Display/n2102 [10]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2124 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4001  (
    .i0(\u2_Display/n2090 ),
    .i1(\u2_Display/n2102 [9]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2125 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4002  (
    .i0(\u2_Display/n2091 ),
    .i1(\u2_Display/n2102 [8]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2126 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4003  (
    .i0(\u2_Display/n2092 ),
    .i1(\u2_Display/n2102 [7]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2127 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4004  (
    .i0(\u2_Display/n2093 ),
    .i1(\u2_Display/n2102 [6]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2128 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4005  (
    .i0(\u2_Display/n2094 ),
    .i1(\u2_Display/n2102 [5]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2129 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4006  (
    .i0(\u2_Display/n2095 ),
    .i1(\u2_Display/n2102 [4]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2130 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4007  (
    .i0(\u2_Display/n2096 ),
    .i1(\u2_Display/n2102 [3]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2131 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4008  (
    .i0(\u2_Display/n2097 ),
    .i1(\u2_Display/n2102 [2]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2132 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4009  (
    .i0(\u2_Display/n2098 ),
    .i1(\u2_Display/n2102 [1]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2133 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4010  (
    .i0(\u2_Display/n2099 ),
    .i1(\u2_Display/n2102 [0]),
    .sel(\u2_Display/n2101 ),
    .o(\u2_Display/n2134 ));  // source/rtl/Display.v(213)
  not \u2_Display/u4011  (\u2_Display/n2136 , \u2_Display/n2135 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4044  (
    .i0(\u2_Display/n2103 ),
    .i1(\u2_Display/n2137 [31]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2138 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4045  (
    .i0(\u2_Display/n2104 ),
    .i1(\u2_Display/n2137 [30]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2139 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4046  (
    .i0(\u2_Display/n2105 ),
    .i1(\u2_Display/n2137 [29]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2140 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4047  (
    .i0(\u2_Display/n2106 ),
    .i1(\u2_Display/n2137 [28]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2141 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4048  (
    .i0(\u2_Display/n2107 ),
    .i1(\u2_Display/n2137 [27]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2142 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4049  (
    .i0(\u2_Display/n2108 ),
    .i1(\u2_Display/n2137 [26]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2143 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4050  (
    .i0(\u2_Display/n2109 ),
    .i1(\u2_Display/n2137 [25]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2144 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4051  (
    .i0(\u2_Display/n2110 ),
    .i1(\u2_Display/n2137 [24]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2145 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4052  (
    .i0(\u2_Display/n2111 ),
    .i1(\u2_Display/n2137 [23]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2146 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4053  (
    .i0(\u2_Display/n2112 ),
    .i1(\u2_Display/n2137 [22]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2147 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4054  (
    .i0(\u2_Display/n2113 ),
    .i1(\u2_Display/n2137 [21]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2148 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4055  (
    .i0(\u2_Display/n2114 ),
    .i1(\u2_Display/n2137 [20]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2149 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4056  (
    .i0(\u2_Display/n2115 ),
    .i1(\u2_Display/n2137 [19]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2150 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4057  (
    .i0(\u2_Display/n2116 ),
    .i1(\u2_Display/n2137 [18]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2151 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4058  (
    .i0(\u2_Display/n2117 ),
    .i1(\u2_Display/n2137 [17]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2152 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4059  (
    .i0(\u2_Display/n2118 ),
    .i1(\u2_Display/n2137 [16]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2153 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4060  (
    .i0(\u2_Display/n2119 ),
    .i1(\u2_Display/n2137 [15]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2154 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4061  (
    .i0(\u2_Display/n2120 ),
    .i1(\u2_Display/n2137 [14]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2155 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4062  (
    .i0(\u2_Display/n2121 ),
    .i1(\u2_Display/n2137 [13]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2156 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4063  (
    .i0(\u2_Display/n2122 ),
    .i1(\u2_Display/n2137 [12]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2157 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4064  (
    .i0(\u2_Display/n2123 ),
    .i1(\u2_Display/n2137 [11]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2158 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4065  (
    .i0(\u2_Display/n2124 ),
    .i1(\u2_Display/n2137 [10]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2159 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4066  (
    .i0(\u2_Display/n2125 ),
    .i1(\u2_Display/n2137 [9]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2160 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4067  (
    .i0(\u2_Display/n2126 ),
    .i1(\u2_Display/n2137 [8]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2161 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4068  (
    .i0(\u2_Display/n2127 ),
    .i1(\u2_Display/n2137 [7]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2162 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4069  (
    .i0(\u2_Display/n2128 ),
    .i1(\u2_Display/n2137 [6]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2163 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4070  (
    .i0(\u2_Display/n2129 ),
    .i1(\u2_Display/n2137 [5]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2164 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4071  (
    .i0(\u2_Display/n2130 ),
    .i1(\u2_Display/n2137 [4]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2165 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4072  (
    .i0(\u2_Display/n2131 ),
    .i1(\u2_Display/n2137 [3]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2166 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4073  (
    .i0(\u2_Display/n2132 ),
    .i1(\u2_Display/n2137 [2]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2167 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4074  (
    .i0(\u2_Display/n2133 ),
    .i1(\u2_Display/n2137 [1]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2168 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4075  (
    .i0(\u2_Display/n2134 ),
    .i1(\u2_Display/n2137 [0]),
    .sel(\u2_Display/n2136 ),
    .o(\u2_Display/n2169 ));  // source/rtl/Display.v(213)
  not \u2_Display/u4076  (\u2_Display/n2171 , \u2_Display/n2170 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4109  (
    .i0(\u2_Display/n2138 ),
    .i1(\u2_Display/n2172 [31]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2173 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4110  (
    .i0(\u2_Display/n2139 ),
    .i1(\u2_Display/n2172 [30]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2174 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4111  (
    .i0(\u2_Display/n2140 ),
    .i1(\u2_Display/n2172 [29]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2175 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4112  (
    .i0(\u2_Display/n2141 ),
    .i1(\u2_Display/n2172 [28]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2176 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4113  (
    .i0(\u2_Display/n2142 ),
    .i1(\u2_Display/n2172 [27]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2177 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4114  (
    .i0(\u2_Display/n2143 ),
    .i1(\u2_Display/n2172 [26]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2178 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4115  (
    .i0(\u2_Display/n2144 ),
    .i1(\u2_Display/n2172 [25]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2179 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4116  (
    .i0(\u2_Display/n2145 ),
    .i1(\u2_Display/n2172 [24]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2180 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4117  (
    .i0(\u2_Display/n2146 ),
    .i1(\u2_Display/n2172 [23]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2181 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4118  (
    .i0(\u2_Display/n2147 ),
    .i1(\u2_Display/n2172 [22]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2182 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4119  (
    .i0(\u2_Display/n2148 ),
    .i1(\u2_Display/n2172 [21]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2183 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4120  (
    .i0(\u2_Display/n2149 ),
    .i1(\u2_Display/n2172 [20]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2184 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4121  (
    .i0(\u2_Display/n2150 ),
    .i1(\u2_Display/n2172 [19]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2185 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4122  (
    .i0(\u2_Display/n2151 ),
    .i1(\u2_Display/n2172 [18]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2186 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4123  (
    .i0(\u2_Display/n2152 ),
    .i1(\u2_Display/n2172 [17]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2187 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4124  (
    .i0(\u2_Display/n2153 ),
    .i1(\u2_Display/n2172 [16]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2188 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4125  (
    .i0(\u2_Display/n2154 ),
    .i1(\u2_Display/n2172 [15]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2189 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4126  (
    .i0(\u2_Display/n2155 ),
    .i1(\u2_Display/n2172 [14]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2190 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4127  (
    .i0(\u2_Display/n2156 ),
    .i1(\u2_Display/n2172 [13]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2191 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4128  (
    .i0(\u2_Display/n2157 ),
    .i1(\u2_Display/n2172 [12]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2192 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4129  (
    .i0(\u2_Display/n2158 ),
    .i1(\u2_Display/n2172 [11]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2193 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4130  (
    .i0(\u2_Display/n2159 ),
    .i1(\u2_Display/n2172 [10]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2194 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4131  (
    .i0(\u2_Display/n2160 ),
    .i1(\u2_Display/n2172 [9]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2195 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4132  (
    .i0(\u2_Display/n2161 ),
    .i1(\u2_Display/n2172 [8]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2196 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4133  (
    .i0(\u2_Display/n2162 ),
    .i1(\u2_Display/n2172 [7]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2197 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4134  (
    .i0(\u2_Display/n2163 ),
    .i1(\u2_Display/n2172 [6]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2198 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4135  (
    .i0(\u2_Display/n2164 ),
    .i1(\u2_Display/n2172 [5]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2199 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4136  (
    .i0(\u2_Display/n2165 ),
    .i1(\u2_Display/n2172 [4]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2200 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4137  (
    .i0(\u2_Display/n2166 ),
    .i1(\u2_Display/n2172 [3]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2201 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4138  (
    .i0(\u2_Display/n2167 ),
    .i1(\u2_Display/n2172 [2]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2202 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4139  (
    .i0(\u2_Display/n2168 ),
    .i1(\u2_Display/n2172 [1]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2203 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4140  (
    .i0(\u2_Display/n2169 ),
    .i1(\u2_Display/n2172 [0]),
    .sel(\u2_Display/n2171 ),
    .o(\u2_Display/n2204 ));  // source/rtl/Display.v(213)
  not \u2_Display/u4141  (\u2_Display/n2206 , \u2_Display/n2205 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4174  (
    .i0(\u2_Display/n2173 ),
    .i1(\u2_Display/n2207 [31]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2208 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4175  (
    .i0(\u2_Display/n2174 ),
    .i1(\u2_Display/n2207 [30]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2209 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4176  (
    .i0(\u2_Display/n2175 ),
    .i1(\u2_Display/n2207 [29]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2210 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4177  (
    .i0(\u2_Display/n2176 ),
    .i1(\u2_Display/n2207 [28]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2211 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4178  (
    .i0(\u2_Display/n2177 ),
    .i1(\u2_Display/n2207 [27]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2212 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4179  (
    .i0(\u2_Display/n2178 ),
    .i1(\u2_Display/n2207 [26]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2213 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4180  (
    .i0(\u2_Display/n2179 ),
    .i1(\u2_Display/n2207 [25]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2214 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4181  (
    .i0(\u2_Display/n2180 ),
    .i1(\u2_Display/n2207 [24]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2215 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4182  (
    .i0(\u2_Display/n2181 ),
    .i1(\u2_Display/n2207 [23]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2216 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4183  (
    .i0(\u2_Display/n2182 ),
    .i1(\u2_Display/n2207 [22]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2217 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4184  (
    .i0(\u2_Display/n2183 ),
    .i1(\u2_Display/n2207 [21]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2218 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4185  (
    .i0(\u2_Display/n2184 ),
    .i1(\u2_Display/n2207 [20]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2219 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4186  (
    .i0(\u2_Display/n2185 ),
    .i1(\u2_Display/n2207 [19]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2220 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4187  (
    .i0(\u2_Display/n2186 ),
    .i1(\u2_Display/n2207 [18]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2221 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4188  (
    .i0(\u2_Display/n2187 ),
    .i1(\u2_Display/n2207 [17]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2222 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4189  (
    .i0(\u2_Display/n2188 ),
    .i1(\u2_Display/n2207 [16]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2223 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4190  (
    .i0(\u2_Display/n2189 ),
    .i1(\u2_Display/n2207 [15]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2224 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4191  (
    .i0(\u2_Display/n2190 ),
    .i1(\u2_Display/n2207 [14]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2225 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4192  (
    .i0(\u2_Display/n2191 ),
    .i1(\u2_Display/n2207 [13]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2226 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4193  (
    .i0(\u2_Display/n2192 ),
    .i1(\u2_Display/n2207 [12]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2227 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4194  (
    .i0(\u2_Display/n2193 ),
    .i1(\u2_Display/n2207 [11]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2228 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4195  (
    .i0(\u2_Display/n2194 ),
    .i1(\u2_Display/n2207 [10]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2229 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4196  (
    .i0(\u2_Display/n2195 ),
    .i1(\u2_Display/n2207 [9]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2230 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4197  (
    .i0(\u2_Display/n2196 ),
    .i1(\u2_Display/n2207 [8]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2231 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4198  (
    .i0(\u2_Display/n2197 ),
    .i1(\u2_Display/n2207 [7]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2232 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4199  (
    .i0(\u2_Display/n2198 ),
    .i1(\u2_Display/n2207 [6]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2233 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4200  (
    .i0(\u2_Display/n2199 ),
    .i1(\u2_Display/n2207 [5]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2234 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4201  (
    .i0(\u2_Display/n2200 ),
    .i1(\u2_Display/n2207 [4]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2235 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4202  (
    .i0(\u2_Display/n2201 ),
    .i1(\u2_Display/n2207 [3]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2236 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4203  (
    .i0(\u2_Display/n2202 ),
    .i1(\u2_Display/n2207 [2]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2237 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4204  (
    .i0(\u2_Display/n2203 ),
    .i1(\u2_Display/n2207 [1]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2238 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4205  (
    .i0(\u2_Display/n2204 ),
    .i1(\u2_Display/n2207 [0]),
    .sel(\u2_Display/n2206 ),
    .o(\u2_Display/n2239 ));  // source/rtl/Display.v(213)
  not \u2_Display/u4206  (\u2_Display/n2241 , \u2_Display/n2240 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4239  (
    .i0(\u2_Display/n2208 ),
    .i1(\u2_Display/n2242 [31]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2243 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4240  (
    .i0(\u2_Display/n2209 ),
    .i1(\u2_Display/n2242 [30]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2244 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4241  (
    .i0(\u2_Display/n2210 ),
    .i1(\u2_Display/n2242 [29]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2245 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4242  (
    .i0(\u2_Display/n2211 ),
    .i1(\u2_Display/n2242 [28]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2246 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4243  (
    .i0(\u2_Display/n2212 ),
    .i1(\u2_Display/n2242 [27]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2247 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4244  (
    .i0(\u2_Display/n2213 ),
    .i1(\u2_Display/n2242 [26]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2248 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4245  (
    .i0(\u2_Display/n2214 ),
    .i1(\u2_Display/n2242 [25]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2249 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4246  (
    .i0(\u2_Display/n2215 ),
    .i1(\u2_Display/n2242 [24]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2250 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4247  (
    .i0(\u2_Display/n2216 ),
    .i1(\u2_Display/n2242 [23]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2251 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4248  (
    .i0(\u2_Display/n2217 ),
    .i1(\u2_Display/n2242 [22]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2252 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4249  (
    .i0(\u2_Display/n2218 ),
    .i1(\u2_Display/n2242 [21]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2253 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4250  (
    .i0(\u2_Display/n2219 ),
    .i1(\u2_Display/n2242 [20]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2254 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4251  (
    .i0(\u2_Display/n2220 ),
    .i1(\u2_Display/n2242 [19]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2255 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4252  (
    .i0(\u2_Display/n2221 ),
    .i1(\u2_Display/n2242 [18]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2256 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4253  (
    .i0(\u2_Display/n2222 ),
    .i1(\u2_Display/n2242 [17]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2257 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4254  (
    .i0(\u2_Display/n2223 ),
    .i1(\u2_Display/n2242 [16]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2258 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4255  (
    .i0(\u2_Display/n2224 ),
    .i1(\u2_Display/n2242 [15]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2259 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4256  (
    .i0(\u2_Display/n2225 ),
    .i1(\u2_Display/n2242 [14]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2260 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4257  (
    .i0(\u2_Display/n2226 ),
    .i1(\u2_Display/n2242 [13]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2261 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4258  (
    .i0(\u2_Display/n2227 ),
    .i1(\u2_Display/n2242 [12]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2262 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4259  (
    .i0(\u2_Display/n2228 ),
    .i1(\u2_Display/n2242 [11]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2263 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4260  (
    .i0(\u2_Display/n2229 ),
    .i1(\u2_Display/n2242 [10]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2264 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4261  (
    .i0(\u2_Display/n2230 ),
    .i1(\u2_Display/n2242 [9]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2265 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4262  (
    .i0(\u2_Display/n2231 ),
    .i1(\u2_Display/n2242 [8]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2266 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4263  (
    .i0(\u2_Display/n2232 ),
    .i1(\u2_Display/n2242 [7]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2267 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4264  (
    .i0(\u2_Display/n2233 ),
    .i1(\u2_Display/n2242 [6]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2268 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4265  (
    .i0(\u2_Display/n2234 ),
    .i1(\u2_Display/n2242 [5]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2269 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4266  (
    .i0(\u2_Display/n2235 ),
    .i1(\u2_Display/n2242 [4]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2270 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4267  (
    .i0(\u2_Display/n2236 ),
    .i1(\u2_Display/n2242 [3]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2271 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4268  (
    .i0(\u2_Display/n2237 ),
    .i1(\u2_Display/n2242 [2]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2272 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4269  (
    .i0(\u2_Display/n2238 ),
    .i1(\u2_Display/n2242 [1]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2273 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4270  (
    .i0(\u2_Display/n2239 ),
    .i1(\u2_Display/n2242 [0]),
    .sel(\u2_Display/n2241 ),
    .o(\u2_Display/n2274 ));  // source/rtl/Display.v(213)
  not \u2_Display/u4271  (\u2_Display/n2276 , \u2_Display/n2275 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4304  (
    .i0(\u2_Display/n2243 ),
    .i1(\u2_Display/n2277 [31]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2278 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4305  (
    .i0(\u2_Display/n2244 ),
    .i1(\u2_Display/n2277 [30]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2279 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4306  (
    .i0(\u2_Display/n2245 ),
    .i1(\u2_Display/n2277 [29]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2280 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4307  (
    .i0(\u2_Display/n2246 ),
    .i1(\u2_Display/n2277 [28]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2281 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4308  (
    .i0(\u2_Display/n2247 ),
    .i1(\u2_Display/n2277 [27]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2282 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4309  (
    .i0(\u2_Display/n2248 ),
    .i1(\u2_Display/n2277 [26]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2283 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4310  (
    .i0(\u2_Display/n2249 ),
    .i1(\u2_Display/n2277 [25]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2284 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4311  (
    .i0(\u2_Display/n2250 ),
    .i1(\u2_Display/n2277 [24]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2285 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4312  (
    .i0(\u2_Display/n2251 ),
    .i1(\u2_Display/n2277 [23]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2286 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4313  (
    .i0(\u2_Display/n2252 ),
    .i1(\u2_Display/n2277 [22]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2287 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4314  (
    .i0(\u2_Display/n2253 ),
    .i1(\u2_Display/n2277 [21]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2288 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4315  (
    .i0(\u2_Display/n2254 ),
    .i1(\u2_Display/n2277 [20]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2289 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4316  (
    .i0(\u2_Display/n2255 ),
    .i1(\u2_Display/n2277 [19]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2290 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4317  (
    .i0(\u2_Display/n2256 ),
    .i1(\u2_Display/n2277 [18]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2291 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4318  (
    .i0(\u2_Display/n2257 ),
    .i1(\u2_Display/n2277 [17]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2292 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4319  (
    .i0(\u2_Display/n2258 ),
    .i1(\u2_Display/n2277 [16]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2293 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4320  (
    .i0(\u2_Display/n2259 ),
    .i1(\u2_Display/n2277 [15]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2294 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4321  (
    .i0(\u2_Display/n2260 ),
    .i1(\u2_Display/n2277 [14]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2295 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4322  (
    .i0(\u2_Display/n2261 ),
    .i1(\u2_Display/n2277 [13]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2296 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4323  (
    .i0(\u2_Display/n2262 ),
    .i1(\u2_Display/n2277 [12]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2297 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4324  (
    .i0(\u2_Display/n2263 ),
    .i1(\u2_Display/n2277 [11]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2298 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4325  (
    .i0(\u2_Display/n2264 ),
    .i1(\u2_Display/n2277 [10]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2299 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4326  (
    .i0(\u2_Display/n2265 ),
    .i1(\u2_Display/n2277 [9]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2300 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4327  (
    .i0(\u2_Display/n2266 ),
    .i1(\u2_Display/n2277 [8]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2301 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4328  (
    .i0(\u2_Display/n2267 ),
    .i1(\u2_Display/n2277 [7]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2302 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4329  (
    .i0(\u2_Display/n2268 ),
    .i1(\u2_Display/n2277 [6]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2303 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4330  (
    .i0(\u2_Display/n2269 ),
    .i1(\u2_Display/n2277 [5]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2304 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4331  (
    .i0(\u2_Display/n2270 ),
    .i1(\u2_Display/n2277 [4]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2305 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4332  (
    .i0(\u2_Display/n2271 ),
    .i1(\u2_Display/n2277 [3]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2306 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4333  (
    .i0(\u2_Display/n2272 ),
    .i1(\u2_Display/n2277 [2]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2307 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4334  (
    .i0(\u2_Display/n2273 ),
    .i1(\u2_Display/n2277 [1]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2308 ));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4335  (
    .i0(\u2_Display/n2274 ),
    .i1(\u2_Display/n2277 [0]),
    .sel(\u2_Display/n2276 ),
    .o(\u2_Display/n2309 ));  // source/rtl/Display.v(213)
  not \u2_Display/u4336  (\u2_Display/n2311 , \u2_Display/n2310 );  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4369  (
    .i0(\u2_Display/n2300 ),
    .i1(\u2_Display/n2312 [9]),
    .sel(\u2_Display/n2311 ),
    .o(\u2_Display/n147 [9]));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4370  (
    .i0(\u2_Display/n2301 ),
    .i1(\u2_Display/n2312 [8]),
    .sel(\u2_Display/n2311 ),
    .o(\u2_Display/n147 [8]));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4371  (
    .i0(\u2_Display/n2302 ),
    .i1(\u2_Display/n2312 [7]),
    .sel(\u2_Display/n2311 ),
    .o(\u2_Display/n147 [7]));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4372  (
    .i0(\u2_Display/n2303 ),
    .i1(\u2_Display/n2312 [6]),
    .sel(\u2_Display/n2311 ),
    .o(\u2_Display/n147 [6]));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4373  (
    .i0(\u2_Display/n2304 ),
    .i1(\u2_Display/n2312 [5]),
    .sel(\u2_Display/n2311 ),
    .o(\u2_Display/n147 [5]));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4374  (
    .i0(\u2_Display/n2305 ),
    .i1(\u2_Display/n2312 [4]),
    .sel(\u2_Display/n2311 ),
    .o(\u2_Display/n147 [4]));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4375  (
    .i0(\u2_Display/n2306 ),
    .i1(\u2_Display/n2312 [3]),
    .sel(\u2_Display/n2311 ),
    .o(\u2_Display/n147 [3]));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4376  (
    .i0(\u2_Display/n2307 ),
    .i1(\u2_Display/n2312 [2]),
    .sel(\u2_Display/n2311 ),
    .o(\u2_Display/n147 [2]));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4377  (
    .i0(\u2_Display/n2308 ),
    .i1(\u2_Display/n2312 [1]),
    .sel(\u2_Display/n2311 ),
    .o(\u2_Display/n147 [1]));  // source/rtl/Display.v(213)
  AL_MUX \u2_Display/u4378  (
    .i0(\u2_Display/n2309 ),
    .i1(\u2_Display/n2312 [0]),
    .sel(\u2_Display/n2311 ),
    .o(\u2_Display/n147 [0]));  // source/rtl/Display.v(213)
  not \u2_Display/u5085  (\u2_Display/n2664 , \u2_Display/n2663 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5118  (
    .i0(\u2_Display/counta [31]),
    .i1(\u2_Display/n2665 [31]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2666 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5119  (
    .i0(\u2_Display/counta [30]),
    .i1(\u2_Display/n2665 [30]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2667 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5120  (
    .i0(\u2_Display/counta [29]),
    .i1(\u2_Display/n2665 [29]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2668 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5121  (
    .i0(\u2_Display/counta [28]),
    .i1(\u2_Display/n2665 [28]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2669 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5122  (
    .i0(\u2_Display/counta [27]),
    .i1(\u2_Display/n2665 [27]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2670 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5123  (
    .i0(\u2_Display/counta [26]),
    .i1(\u2_Display/n2665 [26]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2671 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5124  (
    .i0(\u2_Display/counta [25]),
    .i1(\u2_Display/n2665 [25]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2672 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5125  (
    .i0(\u2_Display/counta [24]),
    .i1(\u2_Display/n2665 [24]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2673 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5126  (
    .i0(\u2_Display/counta [23]),
    .i1(\u2_Display/n2665 [23]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2674 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5127  (
    .i0(\u2_Display/counta [22]),
    .i1(\u2_Display/n2665 [22]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2675 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5128  (
    .i0(\u2_Display/counta [21]),
    .i1(\u2_Display/n2665 [21]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2676 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5129  (
    .i0(\u2_Display/counta [20]),
    .i1(\u2_Display/n2665 [20]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2677 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5130  (
    .i0(\u2_Display/counta [19]),
    .i1(\u2_Display/n2665 [19]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2678 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5131  (
    .i0(\u2_Display/counta [18]),
    .i1(\u2_Display/n2665 [18]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2679 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5132  (
    .i0(\u2_Display/counta [17]),
    .i1(\u2_Display/n2665 [17]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2680 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5133  (
    .i0(\u2_Display/counta [16]),
    .i1(\u2_Display/n2665 [16]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2681 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5134  (
    .i0(\u2_Display/counta [15]),
    .i1(\u2_Display/n2665 [15]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2682 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5135  (
    .i0(\u2_Display/counta [14]),
    .i1(\u2_Display/n2665 [14]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2683 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5136  (
    .i0(\u2_Display/counta [13]),
    .i1(\u2_Display/n2665 [13]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2684 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5137  (
    .i0(\u2_Display/counta [12]),
    .i1(\u2_Display/n2665 [12]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2685 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5138  (
    .i0(\u2_Display/counta [11]),
    .i1(\u2_Display/n2665 [11]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2686 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5139  (
    .i0(\u2_Display/counta [10]),
    .i1(\u2_Display/n2665 [10]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2687 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5140  (
    .i0(\u2_Display/counta [9]),
    .i1(\u2_Display/n2665 [9]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2688 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5141  (
    .i0(\u2_Display/counta [8]),
    .i1(\u2_Display/n2665 [8]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2689 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5142  (
    .i0(\u2_Display/counta [7]),
    .i1(\u2_Display/n2665 [7]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2690 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5143  (
    .i0(\u2_Display/counta [6]),
    .i1(\u2_Display/n2665 [6]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2691 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5144  (
    .i0(\u2_Display/counta [5]),
    .i1(\u2_Display/n2665 [5]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2692 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5145  (
    .i0(\u2_Display/counta [4]),
    .i1(\u2_Display/n2665 [4]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2693 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5146  (
    .i0(\u2_Display/counta [3]),
    .i1(\u2_Display/n2665 [3]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2694 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5147  (
    .i0(\u2_Display/counta [2]),
    .i1(\u2_Display/n2665 [2]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2695 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5148  (
    .i0(\u2_Display/counta [1]),
    .i1(\u2_Display/n2665 [1]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2696 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5149  (
    .i0(\u2_Display/counta [0]),
    .i1(\u2_Display/n2665 [0]),
    .sel(\u2_Display/n2664 ),
    .o(\u2_Display/n2697 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5150  (\u2_Display/n2699 , \u2_Display/n2698 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5183  (
    .i0(\u2_Display/n2666 ),
    .i1(\u2_Display/n2700 [31]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2701 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5184  (
    .i0(\u2_Display/n2667 ),
    .i1(\u2_Display/n2700 [30]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2702 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5185  (
    .i0(\u2_Display/n2668 ),
    .i1(\u2_Display/n2700 [29]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2703 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5186  (
    .i0(\u2_Display/n2669 ),
    .i1(\u2_Display/n2700 [28]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2704 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5187  (
    .i0(\u2_Display/n2670 ),
    .i1(\u2_Display/n2700 [27]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2705 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5188  (
    .i0(\u2_Display/n2671 ),
    .i1(\u2_Display/n2700 [26]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2706 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5189  (
    .i0(\u2_Display/n2672 ),
    .i1(\u2_Display/n2700 [25]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2707 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5190  (
    .i0(\u2_Display/n2673 ),
    .i1(\u2_Display/n2700 [24]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2708 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5191  (
    .i0(\u2_Display/n2674 ),
    .i1(\u2_Display/n2700 [23]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2709 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5192  (
    .i0(\u2_Display/n2675 ),
    .i1(\u2_Display/n2700 [22]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2710 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5193  (
    .i0(\u2_Display/n2676 ),
    .i1(\u2_Display/n2700 [21]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2711 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5194  (
    .i0(\u2_Display/n2677 ),
    .i1(\u2_Display/n2700 [20]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2712 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5195  (
    .i0(\u2_Display/n2678 ),
    .i1(\u2_Display/n2700 [19]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2713 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5196  (
    .i0(\u2_Display/n2679 ),
    .i1(\u2_Display/n2700 [18]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2714 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5197  (
    .i0(\u2_Display/n2680 ),
    .i1(\u2_Display/n2700 [17]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2715 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5198  (
    .i0(\u2_Display/n2681 ),
    .i1(\u2_Display/n2700 [16]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2716 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5199  (
    .i0(\u2_Display/n2682 ),
    .i1(\u2_Display/n2700 [15]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2717 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5200  (
    .i0(\u2_Display/n2683 ),
    .i1(\u2_Display/n2700 [14]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2718 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5201  (
    .i0(\u2_Display/n2684 ),
    .i1(\u2_Display/n2700 [13]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2719 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5202  (
    .i0(\u2_Display/n2685 ),
    .i1(\u2_Display/n2700 [12]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2720 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5203  (
    .i0(\u2_Display/n2686 ),
    .i1(\u2_Display/n2700 [11]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2721 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5204  (
    .i0(\u2_Display/n2687 ),
    .i1(\u2_Display/n2700 [10]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2722 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5205  (
    .i0(\u2_Display/n2688 ),
    .i1(\u2_Display/n2700 [9]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2723 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5206  (
    .i0(\u2_Display/n2689 ),
    .i1(\u2_Display/n2700 [8]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2724 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5207  (
    .i0(\u2_Display/n2690 ),
    .i1(\u2_Display/n2700 [7]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2725 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5208  (
    .i0(\u2_Display/n2691 ),
    .i1(\u2_Display/n2700 [6]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2726 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5209  (
    .i0(\u2_Display/n2692 ),
    .i1(\u2_Display/n2700 [5]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2727 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5210  (
    .i0(\u2_Display/n2693 ),
    .i1(\u2_Display/n2700 [4]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2728 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5211  (
    .i0(\u2_Display/n2694 ),
    .i1(\u2_Display/n2700 [3]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2729 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5212  (
    .i0(\u2_Display/n2695 ),
    .i1(\u2_Display/n2700 [2]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2730 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5213  (
    .i0(\u2_Display/n2696 ),
    .i1(\u2_Display/n2700 [1]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2731 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5214  (
    .i0(\u2_Display/n2697 ),
    .i1(\u2_Display/n2700 [0]),
    .sel(\u2_Display/n2699 ),
    .o(\u2_Display/n2732 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5215  (\u2_Display/n2734 , \u2_Display/n2733 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5248  (
    .i0(\u2_Display/n2701 ),
    .i1(\u2_Display/n2735 [31]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2736 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5249  (
    .i0(\u2_Display/n2702 ),
    .i1(\u2_Display/n2735 [30]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2737 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5250  (
    .i0(\u2_Display/n2703 ),
    .i1(\u2_Display/n2735 [29]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2738 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5251  (
    .i0(\u2_Display/n2704 ),
    .i1(\u2_Display/n2735 [28]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2739 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5252  (
    .i0(\u2_Display/n2705 ),
    .i1(\u2_Display/n2735 [27]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2740 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5253  (
    .i0(\u2_Display/n2706 ),
    .i1(\u2_Display/n2735 [26]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2741 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5254  (
    .i0(\u2_Display/n2707 ),
    .i1(\u2_Display/n2735 [25]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2742 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5255  (
    .i0(\u2_Display/n2708 ),
    .i1(\u2_Display/n2735 [24]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2743 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5256  (
    .i0(\u2_Display/n2709 ),
    .i1(\u2_Display/n2735 [23]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2744 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5257  (
    .i0(\u2_Display/n2710 ),
    .i1(\u2_Display/n2735 [22]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2745 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5258  (
    .i0(\u2_Display/n2711 ),
    .i1(\u2_Display/n2735 [21]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2746 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5259  (
    .i0(\u2_Display/n2712 ),
    .i1(\u2_Display/n2735 [20]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2747 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5260  (
    .i0(\u2_Display/n2713 ),
    .i1(\u2_Display/n2735 [19]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2748 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5261  (
    .i0(\u2_Display/n2714 ),
    .i1(\u2_Display/n2735 [18]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2749 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5262  (
    .i0(\u2_Display/n2715 ),
    .i1(\u2_Display/n2735 [17]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2750 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5263  (
    .i0(\u2_Display/n2716 ),
    .i1(\u2_Display/n2735 [16]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2751 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5264  (
    .i0(\u2_Display/n2717 ),
    .i1(\u2_Display/n2735 [15]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2752 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5265  (
    .i0(\u2_Display/n2718 ),
    .i1(\u2_Display/n2735 [14]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2753 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5266  (
    .i0(\u2_Display/n2719 ),
    .i1(\u2_Display/n2735 [13]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2754 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5267  (
    .i0(\u2_Display/n2720 ),
    .i1(\u2_Display/n2735 [12]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2755 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5268  (
    .i0(\u2_Display/n2721 ),
    .i1(\u2_Display/n2735 [11]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2756 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5269  (
    .i0(\u2_Display/n2722 ),
    .i1(\u2_Display/n2735 [10]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2757 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5270  (
    .i0(\u2_Display/n2723 ),
    .i1(\u2_Display/n2735 [9]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2758 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5271  (
    .i0(\u2_Display/n2724 ),
    .i1(\u2_Display/n2735 [8]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2759 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5272  (
    .i0(\u2_Display/n2725 ),
    .i1(\u2_Display/n2735 [7]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2760 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5273  (
    .i0(\u2_Display/n2726 ),
    .i1(\u2_Display/n2735 [6]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2761 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5274  (
    .i0(\u2_Display/n2727 ),
    .i1(\u2_Display/n2735 [5]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2762 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5275  (
    .i0(\u2_Display/n2728 ),
    .i1(\u2_Display/n2735 [4]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2763 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5276  (
    .i0(\u2_Display/n2729 ),
    .i1(\u2_Display/n2735 [3]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2764 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5277  (
    .i0(\u2_Display/n2730 ),
    .i1(\u2_Display/n2735 [2]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2765 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5278  (
    .i0(\u2_Display/n2731 ),
    .i1(\u2_Display/n2735 [1]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2766 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5279  (
    .i0(\u2_Display/n2732 ),
    .i1(\u2_Display/n2735 [0]),
    .sel(\u2_Display/n2734 ),
    .o(\u2_Display/n2767 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5280  (\u2_Display/n2769 , \u2_Display/n2768 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5313  (
    .i0(\u2_Display/n2736 ),
    .i1(\u2_Display/n2770 [31]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2771 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5314  (
    .i0(\u2_Display/n2737 ),
    .i1(\u2_Display/n2770 [30]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2772 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5315  (
    .i0(\u2_Display/n2738 ),
    .i1(\u2_Display/n2770 [29]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2773 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5316  (
    .i0(\u2_Display/n2739 ),
    .i1(\u2_Display/n2770 [28]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2774 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5317  (
    .i0(\u2_Display/n2740 ),
    .i1(\u2_Display/n2770 [27]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2775 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5318  (
    .i0(\u2_Display/n2741 ),
    .i1(\u2_Display/n2770 [26]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2776 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5319  (
    .i0(\u2_Display/n2742 ),
    .i1(\u2_Display/n2770 [25]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2777 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5320  (
    .i0(\u2_Display/n2743 ),
    .i1(\u2_Display/n2770 [24]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2778 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5321  (
    .i0(\u2_Display/n2744 ),
    .i1(\u2_Display/n2770 [23]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2779 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5322  (
    .i0(\u2_Display/n2745 ),
    .i1(\u2_Display/n2770 [22]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2780 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5323  (
    .i0(\u2_Display/n2746 ),
    .i1(\u2_Display/n2770 [21]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2781 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5324  (
    .i0(\u2_Display/n2747 ),
    .i1(\u2_Display/n2770 [20]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2782 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5325  (
    .i0(\u2_Display/n2748 ),
    .i1(\u2_Display/n2770 [19]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2783 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5326  (
    .i0(\u2_Display/n2749 ),
    .i1(\u2_Display/n2770 [18]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2784 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5327  (
    .i0(\u2_Display/n2750 ),
    .i1(\u2_Display/n2770 [17]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2785 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5328  (
    .i0(\u2_Display/n2751 ),
    .i1(\u2_Display/n2770 [16]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2786 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5329  (
    .i0(\u2_Display/n2752 ),
    .i1(\u2_Display/n2770 [15]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2787 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5330  (
    .i0(\u2_Display/n2753 ),
    .i1(\u2_Display/n2770 [14]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2788 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5331  (
    .i0(\u2_Display/n2754 ),
    .i1(\u2_Display/n2770 [13]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2789 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5332  (
    .i0(\u2_Display/n2755 ),
    .i1(\u2_Display/n2770 [12]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2790 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5333  (
    .i0(\u2_Display/n2756 ),
    .i1(\u2_Display/n2770 [11]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2791 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5334  (
    .i0(\u2_Display/n2757 ),
    .i1(\u2_Display/n2770 [10]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2792 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5335  (
    .i0(\u2_Display/n2758 ),
    .i1(\u2_Display/n2770 [9]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2793 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5336  (
    .i0(\u2_Display/n2759 ),
    .i1(\u2_Display/n2770 [8]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2794 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5337  (
    .i0(\u2_Display/n2760 ),
    .i1(\u2_Display/n2770 [7]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2795 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5338  (
    .i0(\u2_Display/n2761 ),
    .i1(\u2_Display/n2770 [6]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2796 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5339  (
    .i0(\u2_Display/n2762 ),
    .i1(\u2_Display/n2770 [5]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2797 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5340  (
    .i0(\u2_Display/n2763 ),
    .i1(\u2_Display/n2770 [4]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2798 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5341  (
    .i0(\u2_Display/n2764 ),
    .i1(\u2_Display/n2770 [3]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2799 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5342  (
    .i0(\u2_Display/n2765 ),
    .i1(\u2_Display/n2770 [2]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2800 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5343  (
    .i0(\u2_Display/n2766 ),
    .i1(\u2_Display/n2770 [1]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2801 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5344  (
    .i0(\u2_Display/n2767 ),
    .i1(\u2_Display/n2770 [0]),
    .sel(\u2_Display/n2769 ),
    .o(\u2_Display/n2802 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5345  (\u2_Display/n2804 , \u2_Display/n2803 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5378  (
    .i0(\u2_Display/n2771 ),
    .i1(\u2_Display/n2805 [31]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2806 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5379  (
    .i0(\u2_Display/n2772 ),
    .i1(\u2_Display/n2805 [30]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2807 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5380  (
    .i0(\u2_Display/n2773 ),
    .i1(\u2_Display/n2805 [29]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2808 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5381  (
    .i0(\u2_Display/n2774 ),
    .i1(\u2_Display/n2805 [28]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2809 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5382  (
    .i0(\u2_Display/n2775 ),
    .i1(\u2_Display/n2805 [27]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2810 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5383  (
    .i0(\u2_Display/n2776 ),
    .i1(\u2_Display/n2805 [26]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2811 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5384  (
    .i0(\u2_Display/n2777 ),
    .i1(\u2_Display/n2805 [25]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2812 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5385  (
    .i0(\u2_Display/n2778 ),
    .i1(\u2_Display/n2805 [24]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2813 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5386  (
    .i0(\u2_Display/n2779 ),
    .i1(\u2_Display/n2805 [23]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2814 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5387  (
    .i0(\u2_Display/n2780 ),
    .i1(\u2_Display/n2805 [22]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2815 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5388  (
    .i0(\u2_Display/n2781 ),
    .i1(\u2_Display/n2805 [21]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2816 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5389  (
    .i0(\u2_Display/n2782 ),
    .i1(\u2_Display/n2805 [20]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2817 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5390  (
    .i0(\u2_Display/n2783 ),
    .i1(\u2_Display/n2805 [19]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2818 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5391  (
    .i0(\u2_Display/n2784 ),
    .i1(\u2_Display/n2805 [18]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2819 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5392  (
    .i0(\u2_Display/n2785 ),
    .i1(\u2_Display/n2805 [17]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2820 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5393  (
    .i0(\u2_Display/n2786 ),
    .i1(\u2_Display/n2805 [16]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2821 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5394  (
    .i0(\u2_Display/n2787 ),
    .i1(\u2_Display/n2805 [15]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2822 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5395  (
    .i0(\u2_Display/n2788 ),
    .i1(\u2_Display/n2805 [14]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2823 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5396  (
    .i0(\u2_Display/n2789 ),
    .i1(\u2_Display/n2805 [13]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2824 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5397  (
    .i0(\u2_Display/n2790 ),
    .i1(\u2_Display/n2805 [12]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2825 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5398  (
    .i0(\u2_Display/n2791 ),
    .i1(\u2_Display/n2805 [11]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2826 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5399  (
    .i0(\u2_Display/n2792 ),
    .i1(\u2_Display/n2805 [10]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2827 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5400  (
    .i0(\u2_Display/n2793 ),
    .i1(\u2_Display/n2805 [9]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2828 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5401  (
    .i0(\u2_Display/n2794 ),
    .i1(\u2_Display/n2805 [8]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2829 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5402  (
    .i0(\u2_Display/n2795 ),
    .i1(\u2_Display/n2805 [7]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2830 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5403  (
    .i0(\u2_Display/n2796 ),
    .i1(\u2_Display/n2805 [6]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2831 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5404  (
    .i0(\u2_Display/n2797 ),
    .i1(\u2_Display/n2805 [5]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2832 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5405  (
    .i0(\u2_Display/n2798 ),
    .i1(\u2_Display/n2805 [4]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2833 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5406  (
    .i0(\u2_Display/n2799 ),
    .i1(\u2_Display/n2805 [3]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2834 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5407  (
    .i0(\u2_Display/n2800 ),
    .i1(\u2_Display/n2805 [2]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2835 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5408  (
    .i0(\u2_Display/n2801 ),
    .i1(\u2_Display/n2805 [1]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2836 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5409  (
    .i0(\u2_Display/n2802 ),
    .i1(\u2_Display/n2805 [0]),
    .sel(\u2_Display/n2804 ),
    .o(\u2_Display/n2837 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5410  (\u2_Display/n2839 , \u2_Display/n2838 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5443  (
    .i0(\u2_Display/n2806 ),
    .i1(\u2_Display/n2840 [31]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2841 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5444  (
    .i0(\u2_Display/n2807 ),
    .i1(\u2_Display/n2840 [30]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2842 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5445  (
    .i0(\u2_Display/n2808 ),
    .i1(\u2_Display/n2840 [29]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2843 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5446  (
    .i0(\u2_Display/n2809 ),
    .i1(\u2_Display/n2840 [28]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2844 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5447  (
    .i0(\u2_Display/n2810 ),
    .i1(\u2_Display/n2840 [27]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2845 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5448  (
    .i0(\u2_Display/n2811 ),
    .i1(\u2_Display/n2840 [26]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2846 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5449  (
    .i0(\u2_Display/n2812 ),
    .i1(\u2_Display/n2840 [25]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2847 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5450  (
    .i0(\u2_Display/n2813 ),
    .i1(\u2_Display/n2840 [24]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2848 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5451  (
    .i0(\u2_Display/n2814 ),
    .i1(\u2_Display/n2840 [23]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2849 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5452  (
    .i0(\u2_Display/n2815 ),
    .i1(\u2_Display/n2840 [22]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2850 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5453  (
    .i0(\u2_Display/n2816 ),
    .i1(\u2_Display/n2840 [21]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2851 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5454  (
    .i0(\u2_Display/n2817 ),
    .i1(\u2_Display/n2840 [20]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2852 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5455  (
    .i0(\u2_Display/n2818 ),
    .i1(\u2_Display/n2840 [19]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2853 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5456  (
    .i0(\u2_Display/n2819 ),
    .i1(\u2_Display/n2840 [18]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2854 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5457  (
    .i0(\u2_Display/n2820 ),
    .i1(\u2_Display/n2840 [17]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2855 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5458  (
    .i0(\u2_Display/n2821 ),
    .i1(\u2_Display/n2840 [16]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2856 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5459  (
    .i0(\u2_Display/n2822 ),
    .i1(\u2_Display/n2840 [15]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2857 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5460  (
    .i0(\u2_Display/n2823 ),
    .i1(\u2_Display/n2840 [14]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2858 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5461  (
    .i0(\u2_Display/n2824 ),
    .i1(\u2_Display/n2840 [13]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2859 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5462  (
    .i0(\u2_Display/n2825 ),
    .i1(\u2_Display/n2840 [12]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2860 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5463  (
    .i0(\u2_Display/n2826 ),
    .i1(\u2_Display/n2840 [11]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2861 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5464  (
    .i0(\u2_Display/n2827 ),
    .i1(\u2_Display/n2840 [10]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2862 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5465  (
    .i0(\u2_Display/n2828 ),
    .i1(\u2_Display/n2840 [9]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2863 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5466  (
    .i0(\u2_Display/n2829 ),
    .i1(\u2_Display/n2840 [8]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2864 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5467  (
    .i0(\u2_Display/n2830 ),
    .i1(\u2_Display/n2840 [7]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2865 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5468  (
    .i0(\u2_Display/n2831 ),
    .i1(\u2_Display/n2840 [6]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2866 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5469  (
    .i0(\u2_Display/n2832 ),
    .i1(\u2_Display/n2840 [5]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2867 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5470  (
    .i0(\u2_Display/n2833 ),
    .i1(\u2_Display/n2840 [4]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2868 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5471  (
    .i0(\u2_Display/n2834 ),
    .i1(\u2_Display/n2840 [3]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2869 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5472  (
    .i0(\u2_Display/n2835 ),
    .i1(\u2_Display/n2840 [2]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2870 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5473  (
    .i0(\u2_Display/n2836 ),
    .i1(\u2_Display/n2840 [1]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2871 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5474  (
    .i0(\u2_Display/n2837 ),
    .i1(\u2_Display/n2840 [0]),
    .sel(\u2_Display/n2839 ),
    .o(\u2_Display/n2872 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5475  (\u2_Display/n2874 , \u2_Display/n2873 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5508  (
    .i0(\u2_Display/n2841 ),
    .i1(\u2_Display/n2875 [31]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2876 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5509  (
    .i0(\u2_Display/n2842 ),
    .i1(\u2_Display/n2875 [30]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2877 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5510  (
    .i0(\u2_Display/n2843 ),
    .i1(\u2_Display/n2875 [29]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2878 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5511  (
    .i0(\u2_Display/n2844 ),
    .i1(\u2_Display/n2875 [28]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2879 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5512  (
    .i0(\u2_Display/n2845 ),
    .i1(\u2_Display/n2875 [27]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2880 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5513  (
    .i0(\u2_Display/n2846 ),
    .i1(\u2_Display/n2875 [26]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2881 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5514  (
    .i0(\u2_Display/n2847 ),
    .i1(\u2_Display/n2875 [25]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2882 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5515  (
    .i0(\u2_Display/n2848 ),
    .i1(\u2_Display/n2875 [24]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2883 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5516  (
    .i0(\u2_Display/n2849 ),
    .i1(\u2_Display/n2875 [23]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2884 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5517  (
    .i0(\u2_Display/n2850 ),
    .i1(\u2_Display/n2875 [22]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2885 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5518  (
    .i0(\u2_Display/n2851 ),
    .i1(\u2_Display/n2875 [21]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2886 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5519  (
    .i0(\u2_Display/n2852 ),
    .i1(\u2_Display/n2875 [20]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2887 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5520  (
    .i0(\u2_Display/n2853 ),
    .i1(\u2_Display/n2875 [19]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2888 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5521  (
    .i0(\u2_Display/n2854 ),
    .i1(\u2_Display/n2875 [18]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2889 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5522  (
    .i0(\u2_Display/n2855 ),
    .i1(\u2_Display/n2875 [17]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2890 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5523  (
    .i0(\u2_Display/n2856 ),
    .i1(\u2_Display/n2875 [16]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2891 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5524  (
    .i0(\u2_Display/n2857 ),
    .i1(\u2_Display/n2875 [15]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2892 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5525  (
    .i0(\u2_Display/n2858 ),
    .i1(\u2_Display/n2875 [14]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2893 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5526  (
    .i0(\u2_Display/n2859 ),
    .i1(\u2_Display/n2875 [13]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2894 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5527  (
    .i0(\u2_Display/n2860 ),
    .i1(\u2_Display/n2875 [12]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2895 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5528  (
    .i0(\u2_Display/n2861 ),
    .i1(\u2_Display/n2875 [11]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2896 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5529  (
    .i0(\u2_Display/n2862 ),
    .i1(\u2_Display/n2875 [10]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2897 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5530  (
    .i0(\u2_Display/n2863 ),
    .i1(\u2_Display/n2875 [9]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2898 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5531  (
    .i0(\u2_Display/n2864 ),
    .i1(\u2_Display/n2875 [8]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2899 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5532  (
    .i0(\u2_Display/n2865 ),
    .i1(\u2_Display/n2875 [7]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2900 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5533  (
    .i0(\u2_Display/n2866 ),
    .i1(\u2_Display/n2875 [6]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2901 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5534  (
    .i0(\u2_Display/n2867 ),
    .i1(\u2_Display/n2875 [5]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2902 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5535  (
    .i0(\u2_Display/n2868 ),
    .i1(\u2_Display/n2875 [4]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2903 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5536  (
    .i0(\u2_Display/n2869 ),
    .i1(\u2_Display/n2875 [3]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2904 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5537  (
    .i0(\u2_Display/n2870 ),
    .i1(\u2_Display/n2875 [2]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2905 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5538  (
    .i0(\u2_Display/n2871 ),
    .i1(\u2_Display/n2875 [1]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2906 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5539  (
    .i0(\u2_Display/n2872 ),
    .i1(\u2_Display/n2875 [0]),
    .sel(\u2_Display/n2874 ),
    .o(\u2_Display/n2907 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5540  (\u2_Display/n2909 , \u2_Display/n2908 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5573  (
    .i0(\u2_Display/n2876 ),
    .i1(\u2_Display/n2910 [31]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2911 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5574  (
    .i0(\u2_Display/n2877 ),
    .i1(\u2_Display/n2910 [30]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2912 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5575  (
    .i0(\u2_Display/n2878 ),
    .i1(\u2_Display/n2910 [29]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2913 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5576  (
    .i0(\u2_Display/n2879 ),
    .i1(\u2_Display/n2910 [28]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2914 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5577  (
    .i0(\u2_Display/n2880 ),
    .i1(\u2_Display/n2910 [27]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2915 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5578  (
    .i0(\u2_Display/n2881 ),
    .i1(\u2_Display/n2910 [26]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2916 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5579  (
    .i0(\u2_Display/n2882 ),
    .i1(\u2_Display/n2910 [25]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2917 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5580  (
    .i0(\u2_Display/n2883 ),
    .i1(\u2_Display/n2910 [24]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2918 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5581  (
    .i0(\u2_Display/n2884 ),
    .i1(\u2_Display/n2910 [23]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2919 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5582  (
    .i0(\u2_Display/n2885 ),
    .i1(\u2_Display/n2910 [22]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2920 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5583  (
    .i0(\u2_Display/n2886 ),
    .i1(\u2_Display/n2910 [21]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2921 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5584  (
    .i0(\u2_Display/n2887 ),
    .i1(\u2_Display/n2910 [20]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2922 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5585  (
    .i0(\u2_Display/n2888 ),
    .i1(\u2_Display/n2910 [19]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2923 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5586  (
    .i0(\u2_Display/n2889 ),
    .i1(\u2_Display/n2910 [18]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2924 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5587  (
    .i0(\u2_Display/n2890 ),
    .i1(\u2_Display/n2910 [17]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2925 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5588  (
    .i0(\u2_Display/n2891 ),
    .i1(\u2_Display/n2910 [16]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2926 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5589  (
    .i0(\u2_Display/n2892 ),
    .i1(\u2_Display/n2910 [15]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2927 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5590  (
    .i0(\u2_Display/n2893 ),
    .i1(\u2_Display/n2910 [14]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2928 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5591  (
    .i0(\u2_Display/n2894 ),
    .i1(\u2_Display/n2910 [13]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2929 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5592  (
    .i0(\u2_Display/n2895 ),
    .i1(\u2_Display/n2910 [12]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2930 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5593  (
    .i0(\u2_Display/n2896 ),
    .i1(\u2_Display/n2910 [11]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2931 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5594  (
    .i0(\u2_Display/n2897 ),
    .i1(\u2_Display/n2910 [10]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2932 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5595  (
    .i0(\u2_Display/n2898 ),
    .i1(\u2_Display/n2910 [9]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2933 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5596  (
    .i0(\u2_Display/n2899 ),
    .i1(\u2_Display/n2910 [8]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2934 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5597  (
    .i0(\u2_Display/n2900 ),
    .i1(\u2_Display/n2910 [7]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2935 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5598  (
    .i0(\u2_Display/n2901 ),
    .i1(\u2_Display/n2910 [6]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2936 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5599  (
    .i0(\u2_Display/n2902 ),
    .i1(\u2_Display/n2910 [5]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2937 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5600  (
    .i0(\u2_Display/n2903 ),
    .i1(\u2_Display/n2910 [4]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2938 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5601  (
    .i0(\u2_Display/n2904 ),
    .i1(\u2_Display/n2910 [3]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2939 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5602  (
    .i0(\u2_Display/n2905 ),
    .i1(\u2_Display/n2910 [2]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2940 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5603  (
    .i0(\u2_Display/n2906 ),
    .i1(\u2_Display/n2910 [1]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2941 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5604  (
    .i0(\u2_Display/n2907 ),
    .i1(\u2_Display/n2910 [0]),
    .sel(\u2_Display/n2909 ),
    .o(\u2_Display/n2942 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5605  (\u2_Display/n2944 , \u2_Display/n2943 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5638  (
    .i0(\u2_Display/n2911 ),
    .i1(\u2_Display/n2945 [31]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2946 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5639  (
    .i0(\u2_Display/n2912 ),
    .i1(\u2_Display/n2945 [30]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2947 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5640  (
    .i0(\u2_Display/n2913 ),
    .i1(\u2_Display/n2945 [29]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2948 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5641  (
    .i0(\u2_Display/n2914 ),
    .i1(\u2_Display/n2945 [28]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2949 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5642  (
    .i0(\u2_Display/n2915 ),
    .i1(\u2_Display/n2945 [27]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2950 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5643  (
    .i0(\u2_Display/n2916 ),
    .i1(\u2_Display/n2945 [26]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2951 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5644  (
    .i0(\u2_Display/n2917 ),
    .i1(\u2_Display/n2945 [25]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2952 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5645  (
    .i0(\u2_Display/n2918 ),
    .i1(\u2_Display/n2945 [24]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2953 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5646  (
    .i0(\u2_Display/n2919 ),
    .i1(\u2_Display/n2945 [23]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2954 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5647  (
    .i0(\u2_Display/n2920 ),
    .i1(\u2_Display/n2945 [22]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2955 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5648  (
    .i0(\u2_Display/n2921 ),
    .i1(\u2_Display/n2945 [21]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2956 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5649  (
    .i0(\u2_Display/n2922 ),
    .i1(\u2_Display/n2945 [20]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2957 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5650  (
    .i0(\u2_Display/n2923 ),
    .i1(\u2_Display/n2945 [19]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2958 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5651  (
    .i0(\u2_Display/n2924 ),
    .i1(\u2_Display/n2945 [18]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2959 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5652  (
    .i0(\u2_Display/n2925 ),
    .i1(\u2_Display/n2945 [17]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2960 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5653  (
    .i0(\u2_Display/n2926 ),
    .i1(\u2_Display/n2945 [16]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2961 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5654  (
    .i0(\u2_Display/n2927 ),
    .i1(\u2_Display/n2945 [15]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2962 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5655  (
    .i0(\u2_Display/n2928 ),
    .i1(\u2_Display/n2945 [14]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2963 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5656  (
    .i0(\u2_Display/n2929 ),
    .i1(\u2_Display/n2945 [13]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2964 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5657  (
    .i0(\u2_Display/n2930 ),
    .i1(\u2_Display/n2945 [12]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2965 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5658  (
    .i0(\u2_Display/n2931 ),
    .i1(\u2_Display/n2945 [11]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2966 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5659  (
    .i0(\u2_Display/n2932 ),
    .i1(\u2_Display/n2945 [10]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2967 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5660  (
    .i0(\u2_Display/n2933 ),
    .i1(\u2_Display/n2945 [9]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2968 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5661  (
    .i0(\u2_Display/n2934 ),
    .i1(\u2_Display/n2945 [8]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2969 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5662  (
    .i0(\u2_Display/n2935 ),
    .i1(\u2_Display/n2945 [7]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2970 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5663  (
    .i0(\u2_Display/n2936 ),
    .i1(\u2_Display/n2945 [6]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2971 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5664  (
    .i0(\u2_Display/n2937 ),
    .i1(\u2_Display/n2945 [5]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2972 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5665  (
    .i0(\u2_Display/n2938 ),
    .i1(\u2_Display/n2945 [4]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2973 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5666  (
    .i0(\u2_Display/n2939 ),
    .i1(\u2_Display/n2945 [3]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2974 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5667  (
    .i0(\u2_Display/n2940 ),
    .i1(\u2_Display/n2945 [2]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2975 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5668  (
    .i0(\u2_Display/n2941 ),
    .i1(\u2_Display/n2945 [1]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2976 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5669  (
    .i0(\u2_Display/n2942 ),
    .i1(\u2_Display/n2945 [0]),
    .sel(\u2_Display/n2944 ),
    .o(\u2_Display/n2977 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5670  (\u2_Display/n2979 , \u2_Display/n2978 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5703  (
    .i0(\u2_Display/n2946 ),
    .i1(\u2_Display/n2980 [31]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2981 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5704  (
    .i0(\u2_Display/n2947 ),
    .i1(\u2_Display/n2980 [30]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2982 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5705  (
    .i0(\u2_Display/n2948 ),
    .i1(\u2_Display/n2980 [29]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2983 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5706  (
    .i0(\u2_Display/n2949 ),
    .i1(\u2_Display/n2980 [28]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2984 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5707  (
    .i0(\u2_Display/n2950 ),
    .i1(\u2_Display/n2980 [27]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2985 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5708  (
    .i0(\u2_Display/n2951 ),
    .i1(\u2_Display/n2980 [26]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2986 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5709  (
    .i0(\u2_Display/n2952 ),
    .i1(\u2_Display/n2980 [25]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2987 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5710  (
    .i0(\u2_Display/n2953 ),
    .i1(\u2_Display/n2980 [24]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2988 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5711  (
    .i0(\u2_Display/n2954 ),
    .i1(\u2_Display/n2980 [23]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2989 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5712  (
    .i0(\u2_Display/n2955 ),
    .i1(\u2_Display/n2980 [22]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2990 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5713  (
    .i0(\u2_Display/n2956 ),
    .i1(\u2_Display/n2980 [21]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2991 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5714  (
    .i0(\u2_Display/n2957 ),
    .i1(\u2_Display/n2980 [20]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2992 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5715  (
    .i0(\u2_Display/n2958 ),
    .i1(\u2_Display/n2980 [19]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2993 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5716  (
    .i0(\u2_Display/n2959 ),
    .i1(\u2_Display/n2980 [18]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2994 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5717  (
    .i0(\u2_Display/n2960 ),
    .i1(\u2_Display/n2980 [17]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2995 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5718  (
    .i0(\u2_Display/n2961 ),
    .i1(\u2_Display/n2980 [16]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2996 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5719  (
    .i0(\u2_Display/n2962 ),
    .i1(\u2_Display/n2980 [15]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2997 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5720  (
    .i0(\u2_Display/n2963 ),
    .i1(\u2_Display/n2980 [14]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2998 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5721  (
    .i0(\u2_Display/n2964 ),
    .i1(\u2_Display/n2980 [13]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n2999 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5722  (
    .i0(\u2_Display/n2965 ),
    .i1(\u2_Display/n2980 [12]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n3000 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5723  (
    .i0(\u2_Display/n2966 ),
    .i1(\u2_Display/n2980 [11]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n3001 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5724  (
    .i0(\u2_Display/n2967 ),
    .i1(\u2_Display/n2980 [10]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n3002 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5725  (
    .i0(\u2_Display/n2968 ),
    .i1(\u2_Display/n2980 [9]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n3003 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5726  (
    .i0(\u2_Display/n2969 ),
    .i1(\u2_Display/n2980 [8]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n3004 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5727  (
    .i0(\u2_Display/n2970 ),
    .i1(\u2_Display/n2980 [7]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n3005 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5728  (
    .i0(\u2_Display/n2971 ),
    .i1(\u2_Display/n2980 [6]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n3006 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5729  (
    .i0(\u2_Display/n2972 ),
    .i1(\u2_Display/n2980 [5]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n3007 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5730  (
    .i0(\u2_Display/n2973 ),
    .i1(\u2_Display/n2980 [4]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n3008 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5731  (
    .i0(\u2_Display/n2974 ),
    .i1(\u2_Display/n2980 [3]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n3009 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5732  (
    .i0(\u2_Display/n2975 ),
    .i1(\u2_Display/n2980 [2]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n3010 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5733  (
    .i0(\u2_Display/n2976 ),
    .i1(\u2_Display/n2980 [1]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n3011 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5734  (
    .i0(\u2_Display/n2977 ),
    .i1(\u2_Display/n2980 [0]),
    .sel(\u2_Display/n2979 ),
    .o(\u2_Display/n3012 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5735  (\u2_Display/n3014 , \u2_Display/n3013 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5768  (
    .i0(\u2_Display/n2981 ),
    .i1(\u2_Display/n3015 [31]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3016 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5769  (
    .i0(\u2_Display/n2982 ),
    .i1(\u2_Display/n3015 [30]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3017 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5770  (
    .i0(\u2_Display/n2983 ),
    .i1(\u2_Display/n3015 [29]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3018 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5771  (
    .i0(\u2_Display/n2984 ),
    .i1(\u2_Display/n3015 [28]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3019 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5772  (
    .i0(\u2_Display/n2985 ),
    .i1(\u2_Display/n3015 [27]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3020 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5773  (
    .i0(\u2_Display/n2986 ),
    .i1(\u2_Display/n3015 [26]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3021 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5774  (
    .i0(\u2_Display/n2987 ),
    .i1(\u2_Display/n3015 [25]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3022 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5775  (
    .i0(\u2_Display/n2988 ),
    .i1(\u2_Display/n3015 [24]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3023 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5776  (
    .i0(\u2_Display/n2989 ),
    .i1(\u2_Display/n3015 [23]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3024 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5777  (
    .i0(\u2_Display/n2990 ),
    .i1(\u2_Display/n3015 [22]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3025 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5778  (
    .i0(\u2_Display/n2991 ),
    .i1(\u2_Display/n3015 [21]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3026 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5779  (
    .i0(\u2_Display/n2992 ),
    .i1(\u2_Display/n3015 [20]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3027 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5780  (
    .i0(\u2_Display/n2993 ),
    .i1(\u2_Display/n3015 [19]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3028 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5781  (
    .i0(\u2_Display/n2994 ),
    .i1(\u2_Display/n3015 [18]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3029 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5782  (
    .i0(\u2_Display/n2995 ),
    .i1(\u2_Display/n3015 [17]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3030 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5783  (
    .i0(\u2_Display/n2996 ),
    .i1(\u2_Display/n3015 [16]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3031 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5784  (
    .i0(\u2_Display/n2997 ),
    .i1(\u2_Display/n3015 [15]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3032 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5785  (
    .i0(\u2_Display/n2998 ),
    .i1(\u2_Display/n3015 [14]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3033 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5786  (
    .i0(\u2_Display/n2999 ),
    .i1(\u2_Display/n3015 [13]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3034 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5787  (
    .i0(\u2_Display/n3000 ),
    .i1(\u2_Display/n3015 [12]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3035 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5788  (
    .i0(\u2_Display/n3001 ),
    .i1(\u2_Display/n3015 [11]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3036 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5789  (
    .i0(\u2_Display/n3002 ),
    .i1(\u2_Display/n3015 [10]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3037 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5790  (
    .i0(\u2_Display/n3003 ),
    .i1(\u2_Display/n3015 [9]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3038 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5791  (
    .i0(\u2_Display/n3004 ),
    .i1(\u2_Display/n3015 [8]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3039 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5792  (
    .i0(\u2_Display/n3005 ),
    .i1(\u2_Display/n3015 [7]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3040 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5793  (
    .i0(\u2_Display/n3006 ),
    .i1(\u2_Display/n3015 [6]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3041 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5794  (
    .i0(\u2_Display/n3007 ),
    .i1(\u2_Display/n3015 [5]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3042 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5795  (
    .i0(\u2_Display/n3008 ),
    .i1(\u2_Display/n3015 [4]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3043 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5796  (
    .i0(\u2_Display/n3009 ),
    .i1(\u2_Display/n3015 [3]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3044 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5797  (
    .i0(\u2_Display/n3010 ),
    .i1(\u2_Display/n3015 [2]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3045 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5798  (
    .i0(\u2_Display/n3011 ),
    .i1(\u2_Display/n3015 [1]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3046 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5799  (
    .i0(\u2_Display/n3012 ),
    .i1(\u2_Display/n3015 [0]),
    .sel(\u2_Display/n3014 ),
    .o(\u2_Display/n3047 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5800  (\u2_Display/n3049 , \u2_Display/n3048 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5833  (
    .i0(\u2_Display/n3016 ),
    .i1(\u2_Display/n3050 [31]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3051 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5834  (
    .i0(\u2_Display/n3017 ),
    .i1(\u2_Display/n3050 [30]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3052 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5835  (
    .i0(\u2_Display/n3018 ),
    .i1(\u2_Display/n3050 [29]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3053 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5836  (
    .i0(\u2_Display/n3019 ),
    .i1(\u2_Display/n3050 [28]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3054 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5837  (
    .i0(\u2_Display/n3020 ),
    .i1(\u2_Display/n3050 [27]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3055 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5838  (
    .i0(\u2_Display/n3021 ),
    .i1(\u2_Display/n3050 [26]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3056 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5839  (
    .i0(\u2_Display/n3022 ),
    .i1(\u2_Display/n3050 [25]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3057 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5840  (
    .i0(\u2_Display/n3023 ),
    .i1(\u2_Display/n3050 [24]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3058 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5841  (
    .i0(\u2_Display/n3024 ),
    .i1(\u2_Display/n3050 [23]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3059 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5842  (
    .i0(\u2_Display/n3025 ),
    .i1(\u2_Display/n3050 [22]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3060 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5843  (
    .i0(\u2_Display/n3026 ),
    .i1(\u2_Display/n3050 [21]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3061 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5844  (
    .i0(\u2_Display/n3027 ),
    .i1(\u2_Display/n3050 [20]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3062 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5845  (
    .i0(\u2_Display/n3028 ),
    .i1(\u2_Display/n3050 [19]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3063 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5846  (
    .i0(\u2_Display/n3029 ),
    .i1(\u2_Display/n3050 [18]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3064 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5847  (
    .i0(\u2_Display/n3030 ),
    .i1(\u2_Display/n3050 [17]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3065 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5848  (
    .i0(\u2_Display/n3031 ),
    .i1(\u2_Display/n3050 [16]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3066 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5849  (
    .i0(\u2_Display/n3032 ),
    .i1(\u2_Display/n3050 [15]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3067 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5850  (
    .i0(\u2_Display/n3033 ),
    .i1(\u2_Display/n3050 [14]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3068 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5851  (
    .i0(\u2_Display/n3034 ),
    .i1(\u2_Display/n3050 [13]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3069 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5852  (
    .i0(\u2_Display/n3035 ),
    .i1(\u2_Display/n3050 [12]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3070 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5853  (
    .i0(\u2_Display/n3036 ),
    .i1(\u2_Display/n3050 [11]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3071 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5854  (
    .i0(\u2_Display/n3037 ),
    .i1(\u2_Display/n3050 [10]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3072 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5855  (
    .i0(\u2_Display/n3038 ),
    .i1(\u2_Display/n3050 [9]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3073 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5856  (
    .i0(\u2_Display/n3039 ),
    .i1(\u2_Display/n3050 [8]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3074 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5857  (
    .i0(\u2_Display/n3040 ),
    .i1(\u2_Display/n3050 [7]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3075 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5858  (
    .i0(\u2_Display/n3041 ),
    .i1(\u2_Display/n3050 [6]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3076 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5859  (
    .i0(\u2_Display/n3042 ),
    .i1(\u2_Display/n3050 [5]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3077 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5860  (
    .i0(\u2_Display/n3043 ),
    .i1(\u2_Display/n3050 [4]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3078 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5861  (
    .i0(\u2_Display/n3044 ),
    .i1(\u2_Display/n3050 [3]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3079 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5862  (
    .i0(\u2_Display/n3045 ),
    .i1(\u2_Display/n3050 [2]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3080 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5863  (
    .i0(\u2_Display/n3046 ),
    .i1(\u2_Display/n3050 [1]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3081 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5864  (
    .i0(\u2_Display/n3047 ),
    .i1(\u2_Display/n3050 [0]),
    .sel(\u2_Display/n3049 ),
    .o(\u2_Display/n3082 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5865  (\u2_Display/n3084 , \u2_Display/n3083 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5898  (
    .i0(\u2_Display/n3051 ),
    .i1(\u2_Display/n3085 [31]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3086 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5899  (
    .i0(\u2_Display/n3052 ),
    .i1(\u2_Display/n3085 [30]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3087 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5900  (
    .i0(\u2_Display/n3053 ),
    .i1(\u2_Display/n3085 [29]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3088 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5901  (
    .i0(\u2_Display/n3054 ),
    .i1(\u2_Display/n3085 [28]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3089 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5902  (
    .i0(\u2_Display/n3055 ),
    .i1(\u2_Display/n3085 [27]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3090 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5903  (
    .i0(\u2_Display/n3056 ),
    .i1(\u2_Display/n3085 [26]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3091 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5904  (
    .i0(\u2_Display/n3057 ),
    .i1(\u2_Display/n3085 [25]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3092 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5905  (
    .i0(\u2_Display/n3058 ),
    .i1(\u2_Display/n3085 [24]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3093 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5906  (
    .i0(\u2_Display/n3059 ),
    .i1(\u2_Display/n3085 [23]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3094 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5907  (
    .i0(\u2_Display/n3060 ),
    .i1(\u2_Display/n3085 [22]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3095 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5908  (
    .i0(\u2_Display/n3061 ),
    .i1(\u2_Display/n3085 [21]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3096 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5909  (
    .i0(\u2_Display/n3062 ),
    .i1(\u2_Display/n3085 [20]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3097 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5910  (
    .i0(\u2_Display/n3063 ),
    .i1(\u2_Display/n3085 [19]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3098 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5911  (
    .i0(\u2_Display/n3064 ),
    .i1(\u2_Display/n3085 [18]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3099 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5912  (
    .i0(\u2_Display/n3065 ),
    .i1(\u2_Display/n3085 [17]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3100 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5913  (
    .i0(\u2_Display/n3066 ),
    .i1(\u2_Display/n3085 [16]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3101 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5914  (
    .i0(\u2_Display/n3067 ),
    .i1(\u2_Display/n3085 [15]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3102 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5915  (
    .i0(\u2_Display/n3068 ),
    .i1(\u2_Display/n3085 [14]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3103 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5916  (
    .i0(\u2_Display/n3069 ),
    .i1(\u2_Display/n3085 [13]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3104 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5917  (
    .i0(\u2_Display/n3070 ),
    .i1(\u2_Display/n3085 [12]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3105 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5918  (
    .i0(\u2_Display/n3071 ),
    .i1(\u2_Display/n3085 [11]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3106 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5919  (
    .i0(\u2_Display/n3072 ),
    .i1(\u2_Display/n3085 [10]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3107 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5920  (
    .i0(\u2_Display/n3073 ),
    .i1(\u2_Display/n3085 [9]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3108 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5921  (
    .i0(\u2_Display/n3074 ),
    .i1(\u2_Display/n3085 [8]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3109 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5922  (
    .i0(\u2_Display/n3075 ),
    .i1(\u2_Display/n3085 [7]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3110 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5923  (
    .i0(\u2_Display/n3076 ),
    .i1(\u2_Display/n3085 [6]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3111 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5924  (
    .i0(\u2_Display/n3077 ),
    .i1(\u2_Display/n3085 [5]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3112 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5925  (
    .i0(\u2_Display/n3078 ),
    .i1(\u2_Display/n3085 [4]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3113 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5926  (
    .i0(\u2_Display/n3079 ),
    .i1(\u2_Display/n3085 [3]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3114 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5927  (
    .i0(\u2_Display/n3080 ),
    .i1(\u2_Display/n3085 [2]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3115 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5928  (
    .i0(\u2_Display/n3081 ),
    .i1(\u2_Display/n3085 [1]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3116 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5929  (
    .i0(\u2_Display/n3082 ),
    .i1(\u2_Display/n3085 [0]),
    .sel(\u2_Display/n3084 ),
    .o(\u2_Display/n3117 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5930  (\u2_Display/n3119 , \u2_Display/n3118 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5963  (
    .i0(\u2_Display/n3086 ),
    .i1(\u2_Display/n3120 [31]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3121 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5964  (
    .i0(\u2_Display/n3087 ),
    .i1(\u2_Display/n3120 [30]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3122 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5965  (
    .i0(\u2_Display/n3088 ),
    .i1(\u2_Display/n3120 [29]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3123 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5966  (
    .i0(\u2_Display/n3089 ),
    .i1(\u2_Display/n3120 [28]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3124 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5967  (
    .i0(\u2_Display/n3090 ),
    .i1(\u2_Display/n3120 [27]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3125 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5968  (
    .i0(\u2_Display/n3091 ),
    .i1(\u2_Display/n3120 [26]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3126 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5969  (
    .i0(\u2_Display/n3092 ),
    .i1(\u2_Display/n3120 [25]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3127 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5970  (
    .i0(\u2_Display/n3093 ),
    .i1(\u2_Display/n3120 [24]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3128 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5971  (
    .i0(\u2_Display/n3094 ),
    .i1(\u2_Display/n3120 [23]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3129 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5972  (
    .i0(\u2_Display/n3095 ),
    .i1(\u2_Display/n3120 [22]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3130 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5973  (
    .i0(\u2_Display/n3096 ),
    .i1(\u2_Display/n3120 [21]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3131 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5974  (
    .i0(\u2_Display/n3097 ),
    .i1(\u2_Display/n3120 [20]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3132 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5975  (
    .i0(\u2_Display/n3098 ),
    .i1(\u2_Display/n3120 [19]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3133 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5976  (
    .i0(\u2_Display/n3099 ),
    .i1(\u2_Display/n3120 [18]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3134 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5977  (
    .i0(\u2_Display/n3100 ),
    .i1(\u2_Display/n3120 [17]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3135 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5978  (
    .i0(\u2_Display/n3101 ),
    .i1(\u2_Display/n3120 [16]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3136 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5979  (
    .i0(\u2_Display/n3102 ),
    .i1(\u2_Display/n3120 [15]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3137 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5980  (
    .i0(\u2_Display/n3103 ),
    .i1(\u2_Display/n3120 [14]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3138 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5981  (
    .i0(\u2_Display/n3104 ),
    .i1(\u2_Display/n3120 [13]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3139 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5982  (
    .i0(\u2_Display/n3105 ),
    .i1(\u2_Display/n3120 [12]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3140 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5983  (
    .i0(\u2_Display/n3106 ),
    .i1(\u2_Display/n3120 [11]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3141 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5984  (
    .i0(\u2_Display/n3107 ),
    .i1(\u2_Display/n3120 [10]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3142 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5985  (
    .i0(\u2_Display/n3108 ),
    .i1(\u2_Display/n3120 [9]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3143 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5986  (
    .i0(\u2_Display/n3109 ),
    .i1(\u2_Display/n3120 [8]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3144 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5987  (
    .i0(\u2_Display/n3110 ),
    .i1(\u2_Display/n3120 [7]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3145 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5988  (
    .i0(\u2_Display/n3111 ),
    .i1(\u2_Display/n3120 [6]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3146 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5989  (
    .i0(\u2_Display/n3112 ),
    .i1(\u2_Display/n3120 [5]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3147 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5990  (
    .i0(\u2_Display/n3113 ),
    .i1(\u2_Display/n3120 [4]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3148 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5991  (
    .i0(\u2_Display/n3114 ),
    .i1(\u2_Display/n3120 [3]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3149 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5992  (
    .i0(\u2_Display/n3115 ),
    .i1(\u2_Display/n3120 [2]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3150 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5993  (
    .i0(\u2_Display/n3116 ),
    .i1(\u2_Display/n3120 [1]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3151 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u5994  (
    .i0(\u2_Display/n3117 ),
    .i1(\u2_Display/n3120 [0]),
    .sel(\u2_Display/n3119 ),
    .o(\u2_Display/n3152 ));  // source/rtl/Display.v(196)
  not \u2_Display/u5995  (\u2_Display/n3154 , \u2_Display/n3153 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6028  (
    .i0(\u2_Display/n3121 ),
    .i1(\u2_Display/n3155 [31]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3156 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6029  (
    .i0(\u2_Display/n3122 ),
    .i1(\u2_Display/n3155 [30]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3157 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6030  (
    .i0(\u2_Display/n3123 ),
    .i1(\u2_Display/n3155 [29]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3158 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6031  (
    .i0(\u2_Display/n3124 ),
    .i1(\u2_Display/n3155 [28]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3159 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6032  (
    .i0(\u2_Display/n3125 ),
    .i1(\u2_Display/n3155 [27]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3160 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6033  (
    .i0(\u2_Display/n3126 ),
    .i1(\u2_Display/n3155 [26]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3161 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6034  (
    .i0(\u2_Display/n3127 ),
    .i1(\u2_Display/n3155 [25]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3162 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6035  (
    .i0(\u2_Display/n3128 ),
    .i1(\u2_Display/n3155 [24]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3163 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6036  (
    .i0(\u2_Display/n3129 ),
    .i1(\u2_Display/n3155 [23]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3164 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6037  (
    .i0(\u2_Display/n3130 ),
    .i1(\u2_Display/n3155 [22]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3165 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6038  (
    .i0(\u2_Display/n3131 ),
    .i1(\u2_Display/n3155 [21]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3166 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6039  (
    .i0(\u2_Display/n3132 ),
    .i1(\u2_Display/n3155 [20]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3167 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6040  (
    .i0(\u2_Display/n3133 ),
    .i1(\u2_Display/n3155 [19]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3168 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6041  (
    .i0(\u2_Display/n3134 ),
    .i1(\u2_Display/n3155 [18]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3169 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6042  (
    .i0(\u2_Display/n3135 ),
    .i1(\u2_Display/n3155 [17]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3170 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6043  (
    .i0(\u2_Display/n3136 ),
    .i1(\u2_Display/n3155 [16]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3171 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6044  (
    .i0(\u2_Display/n3137 ),
    .i1(\u2_Display/n3155 [15]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3172 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6045  (
    .i0(\u2_Display/n3138 ),
    .i1(\u2_Display/n3155 [14]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3173 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6046  (
    .i0(\u2_Display/n3139 ),
    .i1(\u2_Display/n3155 [13]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3174 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6047  (
    .i0(\u2_Display/n3140 ),
    .i1(\u2_Display/n3155 [12]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3175 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6048  (
    .i0(\u2_Display/n3141 ),
    .i1(\u2_Display/n3155 [11]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3176 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6049  (
    .i0(\u2_Display/n3142 ),
    .i1(\u2_Display/n3155 [10]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3177 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6050  (
    .i0(\u2_Display/n3143 ),
    .i1(\u2_Display/n3155 [9]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3178 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6051  (
    .i0(\u2_Display/n3144 ),
    .i1(\u2_Display/n3155 [8]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3179 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6052  (
    .i0(\u2_Display/n3145 ),
    .i1(\u2_Display/n3155 [7]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3180 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6053  (
    .i0(\u2_Display/n3146 ),
    .i1(\u2_Display/n3155 [6]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3181 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6054  (
    .i0(\u2_Display/n3147 ),
    .i1(\u2_Display/n3155 [5]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3182 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6055  (
    .i0(\u2_Display/n3148 ),
    .i1(\u2_Display/n3155 [4]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3183 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6056  (
    .i0(\u2_Display/n3149 ),
    .i1(\u2_Display/n3155 [3]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3184 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6057  (
    .i0(\u2_Display/n3150 ),
    .i1(\u2_Display/n3155 [2]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3185 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6058  (
    .i0(\u2_Display/n3151 ),
    .i1(\u2_Display/n3155 [1]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3186 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6059  (
    .i0(\u2_Display/n3152 ),
    .i1(\u2_Display/n3155 [0]),
    .sel(\u2_Display/n3154 ),
    .o(\u2_Display/n3187 ));  // source/rtl/Display.v(196)
  not \u2_Display/u6060  (\u2_Display/n3189 , \u2_Display/n3188 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6093  (
    .i0(\u2_Display/n3156 ),
    .i1(\u2_Display/n3190 [31]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3191 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6094  (
    .i0(\u2_Display/n3157 ),
    .i1(\u2_Display/n3190 [30]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3192 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6095  (
    .i0(\u2_Display/n3158 ),
    .i1(\u2_Display/n3190 [29]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3193 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6096  (
    .i0(\u2_Display/n3159 ),
    .i1(\u2_Display/n3190 [28]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3194 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6097  (
    .i0(\u2_Display/n3160 ),
    .i1(\u2_Display/n3190 [27]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3195 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6098  (
    .i0(\u2_Display/n3161 ),
    .i1(\u2_Display/n3190 [26]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3196 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6099  (
    .i0(\u2_Display/n3162 ),
    .i1(\u2_Display/n3190 [25]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3197 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6100  (
    .i0(\u2_Display/n3163 ),
    .i1(\u2_Display/n3190 [24]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3198 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6101  (
    .i0(\u2_Display/n3164 ),
    .i1(\u2_Display/n3190 [23]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3199 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6102  (
    .i0(\u2_Display/n3165 ),
    .i1(\u2_Display/n3190 [22]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3200 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6103  (
    .i0(\u2_Display/n3166 ),
    .i1(\u2_Display/n3190 [21]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3201 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6104  (
    .i0(\u2_Display/n3167 ),
    .i1(\u2_Display/n3190 [20]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3202 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6105  (
    .i0(\u2_Display/n3168 ),
    .i1(\u2_Display/n3190 [19]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3203 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6106  (
    .i0(\u2_Display/n3169 ),
    .i1(\u2_Display/n3190 [18]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3204 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6107  (
    .i0(\u2_Display/n3170 ),
    .i1(\u2_Display/n3190 [17]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3205 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6108  (
    .i0(\u2_Display/n3171 ),
    .i1(\u2_Display/n3190 [16]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3206 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6109  (
    .i0(\u2_Display/n3172 ),
    .i1(\u2_Display/n3190 [15]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3207 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6110  (
    .i0(\u2_Display/n3173 ),
    .i1(\u2_Display/n3190 [14]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3208 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6111  (
    .i0(\u2_Display/n3174 ),
    .i1(\u2_Display/n3190 [13]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3209 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6112  (
    .i0(\u2_Display/n3175 ),
    .i1(\u2_Display/n3190 [12]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3210 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6113  (
    .i0(\u2_Display/n3176 ),
    .i1(\u2_Display/n3190 [11]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3211 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6114  (
    .i0(\u2_Display/n3177 ),
    .i1(\u2_Display/n3190 [10]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3212 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6115  (
    .i0(\u2_Display/n3178 ),
    .i1(\u2_Display/n3190 [9]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3213 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6116  (
    .i0(\u2_Display/n3179 ),
    .i1(\u2_Display/n3190 [8]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3214 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6117  (
    .i0(\u2_Display/n3180 ),
    .i1(\u2_Display/n3190 [7]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3215 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6118  (
    .i0(\u2_Display/n3181 ),
    .i1(\u2_Display/n3190 [6]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3216 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6119  (
    .i0(\u2_Display/n3182 ),
    .i1(\u2_Display/n3190 [5]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3217 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6120  (
    .i0(\u2_Display/n3183 ),
    .i1(\u2_Display/n3190 [4]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3218 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6121  (
    .i0(\u2_Display/n3184 ),
    .i1(\u2_Display/n3190 [3]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3219 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6122  (
    .i0(\u2_Display/n3185 ),
    .i1(\u2_Display/n3190 [2]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3220 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6123  (
    .i0(\u2_Display/n3186 ),
    .i1(\u2_Display/n3190 [1]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3221 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6124  (
    .i0(\u2_Display/n3187 ),
    .i1(\u2_Display/n3190 [0]),
    .sel(\u2_Display/n3189 ),
    .o(\u2_Display/n3222 ));  // source/rtl/Display.v(196)
  not \u2_Display/u6125  (\u2_Display/n3224 , \u2_Display/n3223 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6158  (
    .i0(\u2_Display/n3191 ),
    .i1(\u2_Display/n3225 [31]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3226 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6159  (
    .i0(\u2_Display/n3192 ),
    .i1(\u2_Display/n3225 [30]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3227 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6160  (
    .i0(\u2_Display/n3193 ),
    .i1(\u2_Display/n3225 [29]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3228 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6161  (
    .i0(\u2_Display/n3194 ),
    .i1(\u2_Display/n3225 [28]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3229 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6162  (
    .i0(\u2_Display/n3195 ),
    .i1(\u2_Display/n3225 [27]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3230 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6163  (
    .i0(\u2_Display/n3196 ),
    .i1(\u2_Display/n3225 [26]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3231 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6164  (
    .i0(\u2_Display/n3197 ),
    .i1(\u2_Display/n3225 [25]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3232 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6165  (
    .i0(\u2_Display/n3198 ),
    .i1(\u2_Display/n3225 [24]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3233 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6166  (
    .i0(\u2_Display/n3199 ),
    .i1(\u2_Display/n3225 [23]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3234 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6167  (
    .i0(\u2_Display/n3200 ),
    .i1(\u2_Display/n3225 [22]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3235 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6168  (
    .i0(\u2_Display/n3201 ),
    .i1(\u2_Display/n3225 [21]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3236 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6169  (
    .i0(\u2_Display/n3202 ),
    .i1(\u2_Display/n3225 [20]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3237 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6170  (
    .i0(\u2_Display/n3203 ),
    .i1(\u2_Display/n3225 [19]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3238 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6171  (
    .i0(\u2_Display/n3204 ),
    .i1(\u2_Display/n3225 [18]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3239 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6172  (
    .i0(\u2_Display/n3205 ),
    .i1(\u2_Display/n3225 [17]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3240 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6173  (
    .i0(\u2_Display/n3206 ),
    .i1(\u2_Display/n3225 [16]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3241 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6174  (
    .i0(\u2_Display/n3207 ),
    .i1(\u2_Display/n3225 [15]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3242 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6175  (
    .i0(\u2_Display/n3208 ),
    .i1(\u2_Display/n3225 [14]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3243 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6176  (
    .i0(\u2_Display/n3209 ),
    .i1(\u2_Display/n3225 [13]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3244 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6177  (
    .i0(\u2_Display/n3210 ),
    .i1(\u2_Display/n3225 [12]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3245 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6178  (
    .i0(\u2_Display/n3211 ),
    .i1(\u2_Display/n3225 [11]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3246 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6179  (
    .i0(\u2_Display/n3212 ),
    .i1(\u2_Display/n3225 [10]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3247 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6180  (
    .i0(\u2_Display/n3213 ),
    .i1(\u2_Display/n3225 [9]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3248 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6181  (
    .i0(\u2_Display/n3214 ),
    .i1(\u2_Display/n3225 [8]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3249 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6182  (
    .i0(\u2_Display/n3215 ),
    .i1(\u2_Display/n3225 [7]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3250 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6183  (
    .i0(\u2_Display/n3216 ),
    .i1(\u2_Display/n3225 [6]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3251 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6184  (
    .i0(\u2_Display/n3217 ),
    .i1(\u2_Display/n3225 [5]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3252 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6185  (
    .i0(\u2_Display/n3218 ),
    .i1(\u2_Display/n3225 [4]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3253 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6186  (
    .i0(\u2_Display/n3219 ),
    .i1(\u2_Display/n3225 [3]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3254 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6187  (
    .i0(\u2_Display/n3220 ),
    .i1(\u2_Display/n3225 [2]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3255 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6188  (
    .i0(\u2_Display/n3221 ),
    .i1(\u2_Display/n3225 [1]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3256 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6189  (
    .i0(\u2_Display/n3222 ),
    .i1(\u2_Display/n3225 [0]),
    .sel(\u2_Display/n3224 ),
    .o(\u2_Display/n3257 ));  // source/rtl/Display.v(196)
  not \u2_Display/u6190  (\u2_Display/n3259 , \u2_Display/n3258 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6223  (
    .i0(\u2_Display/n3226 ),
    .i1(\u2_Display/n3260 [31]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3261 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6224  (
    .i0(\u2_Display/n3227 ),
    .i1(\u2_Display/n3260 [30]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3262 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6225  (
    .i0(\u2_Display/n3228 ),
    .i1(\u2_Display/n3260 [29]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3263 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6226  (
    .i0(\u2_Display/n3229 ),
    .i1(\u2_Display/n3260 [28]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3264 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6227  (
    .i0(\u2_Display/n3230 ),
    .i1(\u2_Display/n3260 [27]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3265 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6228  (
    .i0(\u2_Display/n3231 ),
    .i1(\u2_Display/n3260 [26]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3266 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6229  (
    .i0(\u2_Display/n3232 ),
    .i1(\u2_Display/n3260 [25]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3267 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6230  (
    .i0(\u2_Display/n3233 ),
    .i1(\u2_Display/n3260 [24]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3268 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6231  (
    .i0(\u2_Display/n3234 ),
    .i1(\u2_Display/n3260 [23]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3269 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6232  (
    .i0(\u2_Display/n3235 ),
    .i1(\u2_Display/n3260 [22]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3270 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6233  (
    .i0(\u2_Display/n3236 ),
    .i1(\u2_Display/n3260 [21]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3271 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6234  (
    .i0(\u2_Display/n3237 ),
    .i1(\u2_Display/n3260 [20]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3272 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6235  (
    .i0(\u2_Display/n3238 ),
    .i1(\u2_Display/n3260 [19]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3273 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6236  (
    .i0(\u2_Display/n3239 ),
    .i1(\u2_Display/n3260 [18]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3274 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6237  (
    .i0(\u2_Display/n3240 ),
    .i1(\u2_Display/n3260 [17]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3275 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6238  (
    .i0(\u2_Display/n3241 ),
    .i1(\u2_Display/n3260 [16]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3276 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6239  (
    .i0(\u2_Display/n3242 ),
    .i1(\u2_Display/n3260 [15]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3277 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6240  (
    .i0(\u2_Display/n3243 ),
    .i1(\u2_Display/n3260 [14]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3278 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6241  (
    .i0(\u2_Display/n3244 ),
    .i1(\u2_Display/n3260 [13]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3279 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6242  (
    .i0(\u2_Display/n3245 ),
    .i1(\u2_Display/n3260 [12]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3280 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6243  (
    .i0(\u2_Display/n3246 ),
    .i1(\u2_Display/n3260 [11]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3281 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6244  (
    .i0(\u2_Display/n3247 ),
    .i1(\u2_Display/n3260 [10]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3282 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6245  (
    .i0(\u2_Display/n3248 ),
    .i1(\u2_Display/n3260 [9]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3283 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6246  (
    .i0(\u2_Display/n3249 ),
    .i1(\u2_Display/n3260 [8]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3284 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6247  (
    .i0(\u2_Display/n3250 ),
    .i1(\u2_Display/n3260 [7]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3285 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6248  (
    .i0(\u2_Display/n3251 ),
    .i1(\u2_Display/n3260 [6]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3286 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6249  (
    .i0(\u2_Display/n3252 ),
    .i1(\u2_Display/n3260 [5]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3287 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6250  (
    .i0(\u2_Display/n3253 ),
    .i1(\u2_Display/n3260 [4]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3288 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6251  (
    .i0(\u2_Display/n3254 ),
    .i1(\u2_Display/n3260 [3]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3289 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6252  (
    .i0(\u2_Display/n3255 ),
    .i1(\u2_Display/n3260 [2]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3290 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6253  (
    .i0(\u2_Display/n3256 ),
    .i1(\u2_Display/n3260 [1]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3291 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6254  (
    .i0(\u2_Display/n3257 ),
    .i1(\u2_Display/n3260 [0]),
    .sel(\u2_Display/n3259 ),
    .o(\u2_Display/n3292 ));  // source/rtl/Display.v(196)
  not \u2_Display/u6255  (\u2_Display/n3294 , \u2_Display/n3293 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6288  (
    .i0(\u2_Display/n3261 ),
    .i1(\u2_Display/n3295 [31]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3296 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6289  (
    .i0(\u2_Display/n3262 ),
    .i1(\u2_Display/n3295 [30]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3297 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6290  (
    .i0(\u2_Display/n3263 ),
    .i1(\u2_Display/n3295 [29]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3298 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6291  (
    .i0(\u2_Display/n3264 ),
    .i1(\u2_Display/n3295 [28]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3299 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6292  (
    .i0(\u2_Display/n3265 ),
    .i1(\u2_Display/n3295 [27]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3300 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6293  (
    .i0(\u2_Display/n3266 ),
    .i1(\u2_Display/n3295 [26]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3301 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6294  (
    .i0(\u2_Display/n3267 ),
    .i1(\u2_Display/n3295 [25]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3302 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6295  (
    .i0(\u2_Display/n3268 ),
    .i1(\u2_Display/n3295 [24]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3303 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6296  (
    .i0(\u2_Display/n3269 ),
    .i1(\u2_Display/n3295 [23]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3304 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6297  (
    .i0(\u2_Display/n3270 ),
    .i1(\u2_Display/n3295 [22]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3305 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6298  (
    .i0(\u2_Display/n3271 ),
    .i1(\u2_Display/n3295 [21]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3306 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6299  (
    .i0(\u2_Display/n3272 ),
    .i1(\u2_Display/n3295 [20]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3307 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6300  (
    .i0(\u2_Display/n3273 ),
    .i1(\u2_Display/n3295 [19]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3308 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6301  (
    .i0(\u2_Display/n3274 ),
    .i1(\u2_Display/n3295 [18]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3309 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6302  (
    .i0(\u2_Display/n3275 ),
    .i1(\u2_Display/n3295 [17]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3310 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6303  (
    .i0(\u2_Display/n3276 ),
    .i1(\u2_Display/n3295 [16]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3311 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6304  (
    .i0(\u2_Display/n3277 ),
    .i1(\u2_Display/n3295 [15]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3312 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6305  (
    .i0(\u2_Display/n3278 ),
    .i1(\u2_Display/n3295 [14]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3313 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6306  (
    .i0(\u2_Display/n3279 ),
    .i1(\u2_Display/n3295 [13]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3314 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6307  (
    .i0(\u2_Display/n3280 ),
    .i1(\u2_Display/n3295 [12]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3315 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6308  (
    .i0(\u2_Display/n3281 ),
    .i1(\u2_Display/n3295 [11]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3316 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6309  (
    .i0(\u2_Display/n3282 ),
    .i1(\u2_Display/n3295 [10]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3317 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6310  (
    .i0(\u2_Display/n3283 ),
    .i1(\u2_Display/n3295 [9]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3318 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6311  (
    .i0(\u2_Display/n3284 ),
    .i1(\u2_Display/n3295 [8]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3319 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6312  (
    .i0(\u2_Display/n3285 ),
    .i1(\u2_Display/n3295 [7]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3320 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6313  (
    .i0(\u2_Display/n3286 ),
    .i1(\u2_Display/n3295 [6]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3321 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6314  (
    .i0(\u2_Display/n3287 ),
    .i1(\u2_Display/n3295 [5]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3322 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6315  (
    .i0(\u2_Display/n3288 ),
    .i1(\u2_Display/n3295 [4]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3323 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6316  (
    .i0(\u2_Display/n3289 ),
    .i1(\u2_Display/n3295 [3]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3324 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6317  (
    .i0(\u2_Display/n3290 ),
    .i1(\u2_Display/n3295 [2]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3325 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6318  (
    .i0(\u2_Display/n3291 ),
    .i1(\u2_Display/n3295 [1]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3326 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6319  (
    .i0(\u2_Display/n3292 ),
    .i1(\u2_Display/n3295 [0]),
    .sel(\u2_Display/n3294 ),
    .o(\u2_Display/n3327 ));  // source/rtl/Display.v(196)
  not \u2_Display/u6320  (\u2_Display/n3329 , \u2_Display/n3328 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6353  (
    .i0(\u2_Display/n3296 ),
    .i1(\u2_Display/n3330 [31]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3331 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6354  (
    .i0(\u2_Display/n3297 ),
    .i1(\u2_Display/n3330 [30]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3332 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6355  (
    .i0(\u2_Display/n3298 ),
    .i1(\u2_Display/n3330 [29]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3333 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6356  (
    .i0(\u2_Display/n3299 ),
    .i1(\u2_Display/n3330 [28]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3334 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6357  (
    .i0(\u2_Display/n3300 ),
    .i1(\u2_Display/n3330 [27]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3335 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6358  (
    .i0(\u2_Display/n3301 ),
    .i1(\u2_Display/n3330 [26]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3336 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6359  (
    .i0(\u2_Display/n3302 ),
    .i1(\u2_Display/n3330 [25]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3337 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6360  (
    .i0(\u2_Display/n3303 ),
    .i1(\u2_Display/n3330 [24]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3338 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6361  (
    .i0(\u2_Display/n3304 ),
    .i1(\u2_Display/n3330 [23]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3339 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6362  (
    .i0(\u2_Display/n3305 ),
    .i1(\u2_Display/n3330 [22]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3340 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6363  (
    .i0(\u2_Display/n3306 ),
    .i1(\u2_Display/n3330 [21]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3341 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6364  (
    .i0(\u2_Display/n3307 ),
    .i1(\u2_Display/n3330 [20]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3342 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6365  (
    .i0(\u2_Display/n3308 ),
    .i1(\u2_Display/n3330 [19]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3343 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6366  (
    .i0(\u2_Display/n3309 ),
    .i1(\u2_Display/n3330 [18]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3344 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6367  (
    .i0(\u2_Display/n3310 ),
    .i1(\u2_Display/n3330 [17]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3345 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6368  (
    .i0(\u2_Display/n3311 ),
    .i1(\u2_Display/n3330 [16]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3346 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6369  (
    .i0(\u2_Display/n3312 ),
    .i1(\u2_Display/n3330 [15]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3347 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6370  (
    .i0(\u2_Display/n3313 ),
    .i1(\u2_Display/n3330 [14]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3348 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6371  (
    .i0(\u2_Display/n3314 ),
    .i1(\u2_Display/n3330 [13]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3349 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6372  (
    .i0(\u2_Display/n3315 ),
    .i1(\u2_Display/n3330 [12]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3350 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6373  (
    .i0(\u2_Display/n3316 ),
    .i1(\u2_Display/n3330 [11]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3351 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6374  (
    .i0(\u2_Display/n3317 ),
    .i1(\u2_Display/n3330 [10]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3352 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6375  (
    .i0(\u2_Display/n3318 ),
    .i1(\u2_Display/n3330 [9]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3353 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6376  (
    .i0(\u2_Display/n3319 ),
    .i1(\u2_Display/n3330 [8]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3354 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6377  (
    .i0(\u2_Display/n3320 ),
    .i1(\u2_Display/n3330 [7]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3355 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6378  (
    .i0(\u2_Display/n3321 ),
    .i1(\u2_Display/n3330 [6]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3356 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6379  (
    .i0(\u2_Display/n3322 ),
    .i1(\u2_Display/n3330 [5]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3357 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6380  (
    .i0(\u2_Display/n3323 ),
    .i1(\u2_Display/n3330 [4]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3358 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6381  (
    .i0(\u2_Display/n3324 ),
    .i1(\u2_Display/n3330 [3]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3359 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6382  (
    .i0(\u2_Display/n3325 ),
    .i1(\u2_Display/n3330 [2]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3360 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6383  (
    .i0(\u2_Display/n3326 ),
    .i1(\u2_Display/n3330 [1]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3361 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6384  (
    .i0(\u2_Display/n3327 ),
    .i1(\u2_Display/n3330 [0]),
    .sel(\u2_Display/n3329 ),
    .o(\u2_Display/n3362 ));  // source/rtl/Display.v(196)
  not \u2_Display/u6385  (\u2_Display/n3364 , \u2_Display/n3363 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6418  (
    .i0(\u2_Display/n3331 ),
    .i1(\u2_Display/n3365 [31]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3366 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6419  (
    .i0(\u2_Display/n3332 ),
    .i1(\u2_Display/n3365 [30]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3367 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6420  (
    .i0(\u2_Display/n3333 ),
    .i1(\u2_Display/n3365 [29]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3368 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6421  (
    .i0(\u2_Display/n3334 ),
    .i1(\u2_Display/n3365 [28]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3369 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6422  (
    .i0(\u2_Display/n3335 ),
    .i1(\u2_Display/n3365 [27]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3370 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6423  (
    .i0(\u2_Display/n3336 ),
    .i1(\u2_Display/n3365 [26]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3371 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6424  (
    .i0(\u2_Display/n3337 ),
    .i1(\u2_Display/n3365 [25]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3372 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6425  (
    .i0(\u2_Display/n3338 ),
    .i1(\u2_Display/n3365 [24]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3373 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6426  (
    .i0(\u2_Display/n3339 ),
    .i1(\u2_Display/n3365 [23]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3374 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6427  (
    .i0(\u2_Display/n3340 ),
    .i1(\u2_Display/n3365 [22]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3375 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6428  (
    .i0(\u2_Display/n3341 ),
    .i1(\u2_Display/n3365 [21]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3376 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6429  (
    .i0(\u2_Display/n3342 ),
    .i1(\u2_Display/n3365 [20]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3377 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6430  (
    .i0(\u2_Display/n3343 ),
    .i1(\u2_Display/n3365 [19]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3378 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6431  (
    .i0(\u2_Display/n3344 ),
    .i1(\u2_Display/n3365 [18]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3379 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6432  (
    .i0(\u2_Display/n3345 ),
    .i1(\u2_Display/n3365 [17]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3380 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6433  (
    .i0(\u2_Display/n3346 ),
    .i1(\u2_Display/n3365 [16]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3381 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6434  (
    .i0(\u2_Display/n3347 ),
    .i1(\u2_Display/n3365 [15]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3382 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6435  (
    .i0(\u2_Display/n3348 ),
    .i1(\u2_Display/n3365 [14]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3383 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6436  (
    .i0(\u2_Display/n3349 ),
    .i1(\u2_Display/n3365 [13]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3384 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6437  (
    .i0(\u2_Display/n3350 ),
    .i1(\u2_Display/n3365 [12]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3385 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6438  (
    .i0(\u2_Display/n3351 ),
    .i1(\u2_Display/n3365 [11]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3386 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6439  (
    .i0(\u2_Display/n3352 ),
    .i1(\u2_Display/n3365 [10]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3387 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6440  (
    .i0(\u2_Display/n3353 ),
    .i1(\u2_Display/n3365 [9]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3388 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6441  (
    .i0(\u2_Display/n3354 ),
    .i1(\u2_Display/n3365 [8]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3389 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6442  (
    .i0(\u2_Display/n3355 ),
    .i1(\u2_Display/n3365 [7]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3390 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6443  (
    .i0(\u2_Display/n3356 ),
    .i1(\u2_Display/n3365 [6]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3391 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6444  (
    .i0(\u2_Display/n3357 ),
    .i1(\u2_Display/n3365 [5]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3392 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6445  (
    .i0(\u2_Display/n3358 ),
    .i1(\u2_Display/n3365 [4]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3393 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6446  (
    .i0(\u2_Display/n3359 ),
    .i1(\u2_Display/n3365 [3]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3394 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6447  (
    .i0(\u2_Display/n3360 ),
    .i1(\u2_Display/n3365 [2]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3395 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6448  (
    .i0(\u2_Display/n3361 ),
    .i1(\u2_Display/n3365 [1]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3396 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6449  (
    .i0(\u2_Display/n3362 ),
    .i1(\u2_Display/n3365 [0]),
    .sel(\u2_Display/n3364 ),
    .o(\u2_Display/n3397 ));  // source/rtl/Display.v(196)
  not \u2_Display/u6450  (\u2_Display/n3399 , \u2_Display/n3398 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6483  (
    .i0(\u2_Display/n3366 ),
    .i1(\u2_Display/n3400 [31]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3401 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6484  (
    .i0(\u2_Display/n3367 ),
    .i1(\u2_Display/n3400 [30]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3402 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6485  (
    .i0(\u2_Display/n3368 ),
    .i1(\u2_Display/n3400 [29]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3403 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6486  (
    .i0(\u2_Display/n3369 ),
    .i1(\u2_Display/n3400 [28]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3404 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6487  (
    .i0(\u2_Display/n3370 ),
    .i1(\u2_Display/n3400 [27]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3405 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6488  (
    .i0(\u2_Display/n3371 ),
    .i1(\u2_Display/n3400 [26]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3406 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6489  (
    .i0(\u2_Display/n3372 ),
    .i1(\u2_Display/n3400 [25]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3407 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6490  (
    .i0(\u2_Display/n3373 ),
    .i1(\u2_Display/n3400 [24]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3408 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6491  (
    .i0(\u2_Display/n3374 ),
    .i1(\u2_Display/n3400 [23]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3409 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6492  (
    .i0(\u2_Display/n3375 ),
    .i1(\u2_Display/n3400 [22]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3410 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6493  (
    .i0(\u2_Display/n3376 ),
    .i1(\u2_Display/n3400 [21]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3411 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6494  (
    .i0(\u2_Display/n3377 ),
    .i1(\u2_Display/n3400 [20]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3412 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6495  (
    .i0(\u2_Display/n3378 ),
    .i1(\u2_Display/n3400 [19]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3413 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6496  (
    .i0(\u2_Display/n3379 ),
    .i1(\u2_Display/n3400 [18]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3414 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6497  (
    .i0(\u2_Display/n3380 ),
    .i1(\u2_Display/n3400 [17]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3415 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6498  (
    .i0(\u2_Display/n3381 ),
    .i1(\u2_Display/n3400 [16]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3416 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6499  (
    .i0(\u2_Display/n3382 ),
    .i1(\u2_Display/n3400 [15]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3417 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6500  (
    .i0(\u2_Display/n3383 ),
    .i1(\u2_Display/n3400 [14]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3418 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6501  (
    .i0(\u2_Display/n3384 ),
    .i1(\u2_Display/n3400 [13]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3419 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6502  (
    .i0(\u2_Display/n3385 ),
    .i1(\u2_Display/n3400 [12]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3420 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6503  (
    .i0(\u2_Display/n3386 ),
    .i1(\u2_Display/n3400 [11]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3421 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6504  (
    .i0(\u2_Display/n3387 ),
    .i1(\u2_Display/n3400 [10]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3422 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6505  (
    .i0(\u2_Display/n3388 ),
    .i1(\u2_Display/n3400 [9]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3423 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6506  (
    .i0(\u2_Display/n3389 ),
    .i1(\u2_Display/n3400 [8]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3424 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6507  (
    .i0(\u2_Display/n3390 ),
    .i1(\u2_Display/n3400 [7]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3425 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6508  (
    .i0(\u2_Display/n3391 ),
    .i1(\u2_Display/n3400 [6]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3426 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6509  (
    .i0(\u2_Display/n3392 ),
    .i1(\u2_Display/n3400 [5]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3427 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6510  (
    .i0(\u2_Display/n3393 ),
    .i1(\u2_Display/n3400 [4]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3428 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6511  (
    .i0(\u2_Display/n3394 ),
    .i1(\u2_Display/n3400 [3]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3429 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6512  (
    .i0(\u2_Display/n3395 ),
    .i1(\u2_Display/n3400 [2]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3430 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6513  (
    .i0(\u2_Display/n3396 ),
    .i1(\u2_Display/n3400 [1]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3431 ));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6514  (
    .i0(\u2_Display/n3397 ),
    .i1(\u2_Display/n3400 [0]),
    .sel(\u2_Display/n3399 ),
    .o(\u2_Display/n3432 ));  // source/rtl/Display.v(196)
  not \u2_Display/u6515  (\u2_Display/n3434 , \u2_Display/n3433 );  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6548  (
    .i0(\u2_Display/n3423 ),
    .i1(\u2_Display/n3435 [9]),
    .sel(\u2_Display/n3434 ),
    .o(\u2_Display/n134 [9]));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6549  (
    .i0(\u2_Display/n3424 ),
    .i1(\u2_Display/n3435 [8]),
    .sel(\u2_Display/n3434 ),
    .o(\u2_Display/n134 [8]));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6550  (
    .i0(\u2_Display/n3425 ),
    .i1(\u2_Display/n3435 [7]),
    .sel(\u2_Display/n3434 ),
    .o(\u2_Display/n134 [7]));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6551  (
    .i0(\u2_Display/n3426 ),
    .i1(\u2_Display/n3435 [6]),
    .sel(\u2_Display/n3434 ),
    .o(\u2_Display/n134 [6]));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6552  (
    .i0(\u2_Display/n3427 ),
    .i1(\u2_Display/n3435 [5]),
    .sel(\u2_Display/n3434 ),
    .o(\u2_Display/n134 [5]));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6553  (
    .i0(\u2_Display/n3428 ),
    .i1(\u2_Display/n3435 [4]),
    .sel(\u2_Display/n3434 ),
    .o(\u2_Display/n134 [4]));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6554  (
    .i0(\u2_Display/n3429 ),
    .i1(\u2_Display/n3435 [3]),
    .sel(\u2_Display/n3434 ),
    .o(\u2_Display/n134 [3]));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6555  (
    .i0(\u2_Display/n3430 ),
    .i1(\u2_Display/n3435 [2]),
    .sel(\u2_Display/n3434 ),
    .o(\u2_Display/n134 [2]));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6556  (
    .i0(\u2_Display/n3431 ),
    .i1(\u2_Display/n3435 [1]),
    .sel(\u2_Display/n3434 ),
    .o(\u2_Display/n134 [1]));  // source/rtl/Display.v(196)
  AL_MUX \u2_Display/u6557  (
    .i0(\u2_Display/n3432 ),
    .i1(\u2_Display/n3435 [0]),
    .sel(\u2_Display/n3434 ),
    .o(\u2_Display/n134 [0]));  // source/rtl/Display.v(196)
  not \u2_Display/u7264  (\u2_Display/n3787 , \u2_Display/n3786 );  // source/rtl/Display.v(195)
  not \u2_Display/u727  (\u2_Display/n418 , \u2_Display/n417 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7297  (
    .i0(\u2_Display/counta [31]),
    .i1(\u2_Display/n3788 [31]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3789 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7298  (
    .i0(\u2_Display/counta [30]),
    .i1(\u2_Display/n3788 [30]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3790 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7299  (
    .i0(\u2_Display/counta [29]),
    .i1(\u2_Display/n3788 [29]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3791 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7300  (
    .i0(\u2_Display/counta [28]),
    .i1(\u2_Display/n3788 [28]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3792 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7301  (
    .i0(\u2_Display/counta [27]),
    .i1(\u2_Display/n3788 [27]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3793 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7302  (
    .i0(\u2_Display/counta [26]),
    .i1(\u2_Display/n3788 [26]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3794 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7303  (
    .i0(\u2_Display/counta [25]),
    .i1(\u2_Display/n3788 [25]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3795 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7304  (
    .i0(\u2_Display/counta [24]),
    .i1(\u2_Display/n3788 [24]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3796 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7305  (
    .i0(\u2_Display/counta [23]),
    .i1(\u2_Display/n3788 [23]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3797 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7306  (
    .i0(\u2_Display/counta [22]),
    .i1(\u2_Display/n3788 [22]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3798 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7307  (
    .i0(\u2_Display/counta [21]),
    .i1(\u2_Display/n3788 [21]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3799 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7308  (
    .i0(\u2_Display/counta [20]),
    .i1(\u2_Display/n3788 [20]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3800 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7309  (
    .i0(\u2_Display/counta [19]),
    .i1(\u2_Display/n3788 [19]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3801 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7310  (
    .i0(\u2_Display/counta [18]),
    .i1(\u2_Display/n3788 [18]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3802 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7311  (
    .i0(\u2_Display/counta [17]),
    .i1(\u2_Display/n3788 [17]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3803 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7312  (
    .i0(\u2_Display/counta [16]),
    .i1(\u2_Display/n3788 [16]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3804 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7313  (
    .i0(\u2_Display/counta [15]),
    .i1(\u2_Display/n3788 [15]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3805 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7314  (
    .i0(\u2_Display/counta [14]),
    .i1(\u2_Display/n3788 [14]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3806 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7315  (
    .i0(\u2_Display/counta [13]),
    .i1(\u2_Display/n3788 [13]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3807 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7316  (
    .i0(\u2_Display/counta [12]),
    .i1(\u2_Display/n3788 [12]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3808 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7317  (
    .i0(\u2_Display/counta [11]),
    .i1(\u2_Display/n3788 [11]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3809 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7318  (
    .i0(\u2_Display/counta [10]),
    .i1(\u2_Display/n3788 [10]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3810 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7319  (
    .i0(\u2_Display/counta [9]),
    .i1(\u2_Display/n3788 [9]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3811 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7320  (
    .i0(\u2_Display/counta [8]),
    .i1(\u2_Display/n3788 [8]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3812 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7321  (
    .i0(\u2_Display/counta [7]),
    .i1(\u2_Display/n3788 [7]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3813 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7322  (
    .i0(\u2_Display/counta [6]),
    .i1(\u2_Display/n3788 [6]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3814 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7323  (
    .i0(\u2_Display/counta [5]),
    .i1(\u2_Display/n3788 [5]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3815 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7324  (
    .i0(\u2_Display/counta [4]),
    .i1(\u2_Display/n3788 [4]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3816 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7325  (
    .i0(\u2_Display/counta [3]),
    .i1(\u2_Display/n3788 [3]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3817 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7326  (
    .i0(\u2_Display/counta [2]),
    .i1(\u2_Display/n3788 [2]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3818 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7327  (
    .i0(\u2_Display/counta [1]),
    .i1(\u2_Display/n3788 [1]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3819 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7328  (
    .i0(\u2_Display/counta [0]),
    .i1(\u2_Display/n3788 [0]),
    .sel(\u2_Display/n3787 ),
    .o(\u2_Display/n3820 ));  // source/rtl/Display.v(195)
  not \u2_Display/u7329  (\u2_Display/n3822 , \u2_Display/n3821 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7362  (
    .i0(\u2_Display/n3789 ),
    .i1(\u2_Display/n3823 [31]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3824 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7363  (
    .i0(\u2_Display/n3790 ),
    .i1(\u2_Display/n3823 [30]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3825 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7364  (
    .i0(\u2_Display/n3791 ),
    .i1(\u2_Display/n3823 [29]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3826 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7365  (
    .i0(\u2_Display/n3792 ),
    .i1(\u2_Display/n3823 [28]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3827 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7366  (
    .i0(\u2_Display/n3793 ),
    .i1(\u2_Display/n3823 [27]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3828 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7367  (
    .i0(\u2_Display/n3794 ),
    .i1(\u2_Display/n3823 [26]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3829 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7368  (
    .i0(\u2_Display/n3795 ),
    .i1(\u2_Display/n3823 [25]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3830 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7369  (
    .i0(\u2_Display/n3796 ),
    .i1(\u2_Display/n3823 [24]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3831 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7370  (
    .i0(\u2_Display/n3797 ),
    .i1(\u2_Display/n3823 [23]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3832 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7371  (
    .i0(\u2_Display/n3798 ),
    .i1(\u2_Display/n3823 [22]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3833 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7372  (
    .i0(\u2_Display/n3799 ),
    .i1(\u2_Display/n3823 [21]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3834 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7373  (
    .i0(\u2_Display/n3800 ),
    .i1(\u2_Display/n3823 [20]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3835 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7374  (
    .i0(\u2_Display/n3801 ),
    .i1(\u2_Display/n3823 [19]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3836 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7375  (
    .i0(\u2_Display/n3802 ),
    .i1(\u2_Display/n3823 [18]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3837 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7376  (
    .i0(\u2_Display/n3803 ),
    .i1(\u2_Display/n3823 [17]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3838 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7377  (
    .i0(\u2_Display/n3804 ),
    .i1(\u2_Display/n3823 [16]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3839 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7378  (
    .i0(\u2_Display/n3805 ),
    .i1(\u2_Display/n3823 [15]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3840 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7379  (
    .i0(\u2_Display/n3806 ),
    .i1(\u2_Display/n3823 [14]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3841 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7380  (
    .i0(\u2_Display/n3807 ),
    .i1(\u2_Display/n3823 [13]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3842 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7381  (
    .i0(\u2_Display/n3808 ),
    .i1(\u2_Display/n3823 [12]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3843 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7382  (
    .i0(\u2_Display/n3809 ),
    .i1(\u2_Display/n3823 [11]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3844 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7383  (
    .i0(\u2_Display/n3810 ),
    .i1(\u2_Display/n3823 [10]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3845 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7384  (
    .i0(\u2_Display/n3811 ),
    .i1(\u2_Display/n3823 [9]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3846 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7385  (
    .i0(\u2_Display/n3812 ),
    .i1(\u2_Display/n3823 [8]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3847 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7386  (
    .i0(\u2_Display/n3813 ),
    .i1(\u2_Display/n3823 [7]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3848 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7387  (
    .i0(\u2_Display/n3814 ),
    .i1(\u2_Display/n3823 [6]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3849 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7388  (
    .i0(\u2_Display/n3815 ),
    .i1(\u2_Display/n3823 [5]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3850 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7389  (
    .i0(\u2_Display/n3816 ),
    .i1(\u2_Display/n3823 [4]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3851 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7390  (
    .i0(\u2_Display/n3817 ),
    .i1(\u2_Display/n3823 [3]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3852 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7391  (
    .i0(\u2_Display/n3818 ),
    .i1(\u2_Display/n3823 [2]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3853 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7392  (
    .i0(\u2_Display/n3819 ),
    .i1(\u2_Display/n3823 [1]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3854 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7393  (
    .i0(\u2_Display/n3820 ),
    .i1(\u2_Display/n3823 [0]),
    .sel(\u2_Display/n3822 ),
    .o(\u2_Display/n3855 ));  // source/rtl/Display.v(195)
  not \u2_Display/u7394  (\u2_Display/n3857 , \u2_Display/n3856 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7427  (
    .i0(\u2_Display/n3824 ),
    .i1(\u2_Display/n3858 [31]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3859 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7428  (
    .i0(\u2_Display/n3825 ),
    .i1(\u2_Display/n3858 [30]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3860 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7429  (
    .i0(\u2_Display/n3826 ),
    .i1(\u2_Display/n3858 [29]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3861 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7430  (
    .i0(\u2_Display/n3827 ),
    .i1(\u2_Display/n3858 [28]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3862 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7431  (
    .i0(\u2_Display/n3828 ),
    .i1(\u2_Display/n3858 [27]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3863 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7432  (
    .i0(\u2_Display/n3829 ),
    .i1(\u2_Display/n3858 [26]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3864 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7433  (
    .i0(\u2_Display/n3830 ),
    .i1(\u2_Display/n3858 [25]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3865 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7434  (
    .i0(\u2_Display/n3831 ),
    .i1(\u2_Display/n3858 [24]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3866 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7435  (
    .i0(\u2_Display/n3832 ),
    .i1(\u2_Display/n3858 [23]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3867 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7436  (
    .i0(\u2_Display/n3833 ),
    .i1(\u2_Display/n3858 [22]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3868 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7437  (
    .i0(\u2_Display/n3834 ),
    .i1(\u2_Display/n3858 [21]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3869 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7438  (
    .i0(\u2_Display/n3835 ),
    .i1(\u2_Display/n3858 [20]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3870 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7439  (
    .i0(\u2_Display/n3836 ),
    .i1(\u2_Display/n3858 [19]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3871 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7440  (
    .i0(\u2_Display/n3837 ),
    .i1(\u2_Display/n3858 [18]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3872 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7441  (
    .i0(\u2_Display/n3838 ),
    .i1(\u2_Display/n3858 [17]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3873 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7442  (
    .i0(\u2_Display/n3839 ),
    .i1(\u2_Display/n3858 [16]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3874 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7443  (
    .i0(\u2_Display/n3840 ),
    .i1(\u2_Display/n3858 [15]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3875 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7444  (
    .i0(\u2_Display/n3841 ),
    .i1(\u2_Display/n3858 [14]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3876 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7445  (
    .i0(\u2_Display/n3842 ),
    .i1(\u2_Display/n3858 [13]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3877 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7446  (
    .i0(\u2_Display/n3843 ),
    .i1(\u2_Display/n3858 [12]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3878 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7447  (
    .i0(\u2_Display/n3844 ),
    .i1(\u2_Display/n3858 [11]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3879 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7448  (
    .i0(\u2_Display/n3845 ),
    .i1(\u2_Display/n3858 [10]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3880 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7449  (
    .i0(\u2_Display/n3846 ),
    .i1(\u2_Display/n3858 [9]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3881 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7450  (
    .i0(\u2_Display/n3847 ),
    .i1(\u2_Display/n3858 [8]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3882 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7451  (
    .i0(\u2_Display/n3848 ),
    .i1(\u2_Display/n3858 [7]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3883 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7452  (
    .i0(\u2_Display/n3849 ),
    .i1(\u2_Display/n3858 [6]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3884 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7453  (
    .i0(\u2_Display/n3850 ),
    .i1(\u2_Display/n3858 [5]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3885 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7454  (
    .i0(\u2_Display/n3851 ),
    .i1(\u2_Display/n3858 [4]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3886 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7455  (
    .i0(\u2_Display/n3852 ),
    .i1(\u2_Display/n3858 [3]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3887 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7456  (
    .i0(\u2_Display/n3853 ),
    .i1(\u2_Display/n3858 [2]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3888 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7457  (
    .i0(\u2_Display/n3854 ),
    .i1(\u2_Display/n3858 [1]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3889 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7458  (
    .i0(\u2_Display/n3855 ),
    .i1(\u2_Display/n3858 [0]),
    .sel(\u2_Display/n3857 ),
    .o(\u2_Display/n3890 ));  // source/rtl/Display.v(195)
  not \u2_Display/u7459  (\u2_Display/n3892 , \u2_Display/n3891 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7492  (
    .i0(\u2_Display/n3859 ),
    .i1(\u2_Display/n3893 [31]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3894 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7493  (
    .i0(\u2_Display/n3860 ),
    .i1(\u2_Display/n3893 [30]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3895 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7494  (
    .i0(\u2_Display/n3861 ),
    .i1(\u2_Display/n3893 [29]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3896 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7495  (
    .i0(\u2_Display/n3862 ),
    .i1(\u2_Display/n3893 [28]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3897 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7496  (
    .i0(\u2_Display/n3863 ),
    .i1(\u2_Display/n3893 [27]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3898 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7497  (
    .i0(\u2_Display/n3864 ),
    .i1(\u2_Display/n3893 [26]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3899 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7498  (
    .i0(\u2_Display/n3865 ),
    .i1(\u2_Display/n3893 [25]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3900 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7499  (
    .i0(\u2_Display/n3866 ),
    .i1(\u2_Display/n3893 [24]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3901 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7500  (
    .i0(\u2_Display/n3867 ),
    .i1(\u2_Display/n3893 [23]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3902 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7501  (
    .i0(\u2_Display/n3868 ),
    .i1(\u2_Display/n3893 [22]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3903 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7502  (
    .i0(\u2_Display/n3869 ),
    .i1(\u2_Display/n3893 [21]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3904 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7503  (
    .i0(\u2_Display/n3870 ),
    .i1(\u2_Display/n3893 [20]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3905 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7504  (
    .i0(\u2_Display/n3871 ),
    .i1(\u2_Display/n3893 [19]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3906 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7505  (
    .i0(\u2_Display/n3872 ),
    .i1(\u2_Display/n3893 [18]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3907 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7506  (
    .i0(\u2_Display/n3873 ),
    .i1(\u2_Display/n3893 [17]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3908 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7507  (
    .i0(\u2_Display/n3874 ),
    .i1(\u2_Display/n3893 [16]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3909 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7508  (
    .i0(\u2_Display/n3875 ),
    .i1(\u2_Display/n3893 [15]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3910 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7509  (
    .i0(\u2_Display/n3876 ),
    .i1(\u2_Display/n3893 [14]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3911 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7510  (
    .i0(\u2_Display/n3877 ),
    .i1(\u2_Display/n3893 [13]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3912 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7511  (
    .i0(\u2_Display/n3878 ),
    .i1(\u2_Display/n3893 [12]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3913 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7512  (
    .i0(\u2_Display/n3879 ),
    .i1(\u2_Display/n3893 [11]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3914 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7513  (
    .i0(\u2_Display/n3880 ),
    .i1(\u2_Display/n3893 [10]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3915 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7514  (
    .i0(\u2_Display/n3881 ),
    .i1(\u2_Display/n3893 [9]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3916 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7515  (
    .i0(\u2_Display/n3882 ),
    .i1(\u2_Display/n3893 [8]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3917 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7516  (
    .i0(\u2_Display/n3883 ),
    .i1(\u2_Display/n3893 [7]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3918 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7517  (
    .i0(\u2_Display/n3884 ),
    .i1(\u2_Display/n3893 [6]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3919 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7518  (
    .i0(\u2_Display/n3885 ),
    .i1(\u2_Display/n3893 [5]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3920 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7519  (
    .i0(\u2_Display/n3886 ),
    .i1(\u2_Display/n3893 [4]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3921 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7520  (
    .i0(\u2_Display/n3887 ),
    .i1(\u2_Display/n3893 [3]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3922 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7521  (
    .i0(\u2_Display/n3888 ),
    .i1(\u2_Display/n3893 [2]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3923 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7522  (
    .i0(\u2_Display/n3889 ),
    .i1(\u2_Display/n3893 [1]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3924 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7523  (
    .i0(\u2_Display/n3890 ),
    .i1(\u2_Display/n3893 [0]),
    .sel(\u2_Display/n3892 ),
    .o(\u2_Display/n3925 ));  // source/rtl/Display.v(195)
  not \u2_Display/u7524  (\u2_Display/n3927 , \u2_Display/n3926 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7557  (
    .i0(\u2_Display/n3894 ),
    .i1(\u2_Display/n3928 [31]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3929 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7558  (
    .i0(\u2_Display/n3895 ),
    .i1(\u2_Display/n3928 [30]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3930 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7559  (
    .i0(\u2_Display/n3896 ),
    .i1(\u2_Display/n3928 [29]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3931 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7560  (
    .i0(\u2_Display/n3897 ),
    .i1(\u2_Display/n3928 [28]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3932 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7561  (
    .i0(\u2_Display/n3898 ),
    .i1(\u2_Display/n3928 [27]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3933 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7562  (
    .i0(\u2_Display/n3899 ),
    .i1(\u2_Display/n3928 [26]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3934 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7563  (
    .i0(\u2_Display/n3900 ),
    .i1(\u2_Display/n3928 [25]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3935 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7564  (
    .i0(\u2_Display/n3901 ),
    .i1(\u2_Display/n3928 [24]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3936 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7565  (
    .i0(\u2_Display/n3902 ),
    .i1(\u2_Display/n3928 [23]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3937 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7566  (
    .i0(\u2_Display/n3903 ),
    .i1(\u2_Display/n3928 [22]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3938 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7567  (
    .i0(\u2_Display/n3904 ),
    .i1(\u2_Display/n3928 [21]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3939 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7568  (
    .i0(\u2_Display/n3905 ),
    .i1(\u2_Display/n3928 [20]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3940 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7569  (
    .i0(\u2_Display/n3906 ),
    .i1(\u2_Display/n3928 [19]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3941 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7570  (
    .i0(\u2_Display/n3907 ),
    .i1(\u2_Display/n3928 [18]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3942 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7571  (
    .i0(\u2_Display/n3908 ),
    .i1(\u2_Display/n3928 [17]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3943 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7572  (
    .i0(\u2_Display/n3909 ),
    .i1(\u2_Display/n3928 [16]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3944 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7573  (
    .i0(\u2_Display/n3910 ),
    .i1(\u2_Display/n3928 [15]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3945 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7574  (
    .i0(\u2_Display/n3911 ),
    .i1(\u2_Display/n3928 [14]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3946 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7575  (
    .i0(\u2_Display/n3912 ),
    .i1(\u2_Display/n3928 [13]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3947 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7576  (
    .i0(\u2_Display/n3913 ),
    .i1(\u2_Display/n3928 [12]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3948 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7577  (
    .i0(\u2_Display/n3914 ),
    .i1(\u2_Display/n3928 [11]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3949 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7578  (
    .i0(\u2_Display/n3915 ),
    .i1(\u2_Display/n3928 [10]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3950 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7579  (
    .i0(\u2_Display/n3916 ),
    .i1(\u2_Display/n3928 [9]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3951 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7580  (
    .i0(\u2_Display/n3917 ),
    .i1(\u2_Display/n3928 [8]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3952 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7581  (
    .i0(\u2_Display/n3918 ),
    .i1(\u2_Display/n3928 [7]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3953 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7582  (
    .i0(\u2_Display/n3919 ),
    .i1(\u2_Display/n3928 [6]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3954 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7583  (
    .i0(\u2_Display/n3920 ),
    .i1(\u2_Display/n3928 [5]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3955 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7584  (
    .i0(\u2_Display/n3921 ),
    .i1(\u2_Display/n3928 [4]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3956 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7585  (
    .i0(\u2_Display/n3922 ),
    .i1(\u2_Display/n3928 [3]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3957 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7586  (
    .i0(\u2_Display/n3923 ),
    .i1(\u2_Display/n3928 [2]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3958 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7587  (
    .i0(\u2_Display/n3924 ),
    .i1(\u2_Display/n3928 [1]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3959 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7588  (
    .i0(\u2_Display/n3925 ),
    .i1(\u2_Display/n3928 [0]),
    .sel(\u2_Display/n3927 ),
    .o(\u2_Display/n3960 ));  // source/rtl/Display.v(195)
  not \u2_Display/u7589  (\u2_Display/n3962 , \u2_Display/n3961 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u760  (
    .i0(\u2_Display/counta [31]),
    .i1(\u2_Display/n419 [31]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n420 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u761  (
    .i0(\u2_Display/counta [30]),
    .i1(\u2_Display/n419 [30]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n421 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u762  (
    .i0(\u2_Display/counta [29]),
    .i1(\u2_Display/n419 [29]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n422 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7622  (
    .i0(\u2_Display/n3929 ),
    .i1(\u2_Display/n3963 [31]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3964 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7623  (
    .i0(\u2_Display/n3930 ),
    .i1(\u2_Display/n3963 [30]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3965 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7624  (
    .i0(\u2_Display/n3931 ),
    .i1(\u2_Display/n3963 [29]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3966 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7625  (
    .i0(\u2_Display/n3932 ),
    .i1(\u2_Display/n3963 [28]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3967 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7626  (
    .i0(\u2_Display/n3933 ),
    .i1(\u2_Display/n3963 [27]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3968 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7627  (
    .i0(\u2_Display/n3934 ),
    .i1(\u2_Display/n3963 [26]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3969 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7628  (
    .i0(\u2_Display/n3935 ),
    .i1(\u2_Display/n3963 [25]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3970 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7629  (
    .i0(\u2_Display/n3936 ),
    .i1(\u2_Display/n3963 [24]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3971 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u763  (
    .i0(\u2_Display/counta [28]),
    .i1(\u2_Display/n419 [28]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n423 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7630  (
    .i0(\u2_Display/n3937 ),
    .i1(\u2_Display/n3963 [23]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3972 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7631  (
    .i0(\u2_Display/n3938 ),
    .i1(\u2_Display/n3963 [22]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3973 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7632  (
    .i0(\u2_Display/n3939 ),
    .i1(\u2_Display/n3963 [21]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3974 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7633  (
    .i0(\u2_Display/n3940 ),
    .i1(\u2_Display/n3963 [20]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3975 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7634  (
    .i0(\u2_Display/n3941 ),
    .i1(\u2_Display/n3963 [19]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3976 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7635  (
    .i0(\u2_Display/n3942 ),
    .i1(\u2_Display/n3963 [18]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3977 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7636  (
    .i0(\u2_Display/n3943 ),
    .i1(\u2_Display/n3963 [17]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3978 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7637  (
    .i0(\u2_Display/n3944 ),
    .i1(\u2_Display/n3963 [16]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3979 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7638  (
    .i0(\u2_Display/n3945 ),
    .i1(\u2_Display/n3963 [15]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3980 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7639  (
    .i0(\u2_Display/n3946 ),
    .i1(\u2_Display/n3963 [14]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3981 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u764  (
    .i0(\u2_Display/counta [27]),
    .i1(\u2_Display/n419 [27]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n424 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7640  (
    .i0(\u2_Display/n3947 ),
    .i1(\u2_Display/n3963 [13]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3982 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7641  (
    .i0(\u2_Display/n3948 ),
    .i1(\u2_Display/n3963 [12]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3983 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7642  (
    .i0(\u2_Display/n3949 ),
    .i1(\u2_Display/n3963 [11]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3984 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7643  (
    .i0(\u2_Display/n3950 ),
    .i1(\u2_Display/n3963 [10]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3985 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7644  (
    .i0(\u2_Display/n3951 ),
    .i1(\u2_Display/n3963 [9]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3986 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7645  (
    .i0(\u2_Display/n3952 ),
    .i1(\u2_Display/n3963 [8]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3987 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7646  (
    .i0(\u2_Display/n3953 ),
    .i1(\u2_Display/n3963 [7]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3988 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7647  (
    .i0(\u2_Display/n3954 ),
    .i1(\u2_Display/n3963 [6]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3989 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7648  (
    .i0(\u2_Display/n3955 ),
    .i1(\u2_Display/n3963 [5]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3990 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7649  (
    .i0(\u2_Display/n3956 ),
    .i1(\u2_Display/n3963 [4]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3991 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u765  (
    .i0(\u2_Display/counta [26]),
    .i1(\u2_Display/n419 [26]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n425 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7650  (
    .i0(\u2_Display/n3957 ),
    .i1(\u2_Display/n3963 [3]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3992 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7651  (
    .i0(\u2_Display/n3958 ),
    .i1(\u2_Display/n3963 [2]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3993 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7652  (
    .i0(\u2_Display/n3959 ),
    .i1(\u2_Display/n3963 [1]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3994 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7653  (
    .i0(\u2_Display/n3960 ),
    .i1(\u2_Display/n3963 [0]),
    .sel(\u2_Display/n3962 ),
    .o(\u2_Display/n3995 ));  // source/rtl/Display.v(195)
  not \u2_Display/u7654  (\u2_Display/n3997 , \u2_Display/n3996 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u766  (
    .i0(\u2_Display/counta [25]),
    .i1(\u2_Display/n419 [25]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n426 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u767  (
    .i0(\u2_Display/counta [24]),
    .i1(\u2_Display/n419 [24]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n427 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u768  (
    .i0(\u2_Display/counta [23]),
    .i1(\u2_Display/n419 [23]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n428 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7687  (
    .i0(\u2_Display/n3964 ),
    .i1(\u2_Display/n3998 [31]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n3999 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7688  (
    .i0(\u2_Display/n3965 ),
    .i1(\u2_Display/n3998 [30]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4000 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7689  (
    .i0(\u2_Display/n3966 ),
    .i1(\u2_Display/n3998 [29]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4001 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u769  (
    .i0(\u2_Display/counta [22]),
    .i1(\u2_Display/n419 [22]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n429 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7690  (
    .i0(\u2_Display/n3967 ),
    .i1(\u2_Display/n3998 [28]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4002 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7691  (
    .i0(\u2_Display/n3968 ),
    .i1(\u2_Display/n3998 [27]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4003 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7692  (
    .i0(\u2_Display/n3969 ),
    .i1(\u2_Display/n3998 [26]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4004 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7693  (
    .i0(\u2_Display/n3970 ),
    .i1(\u2_Display/n3998 [25]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4005 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7694  (
    .i0(\u2_Display/n3971 ),
    .i1(\u2_Display/n3998 [24]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4006 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7695  (
    .i0(\u2_Display/n3972 ),
    .i1(\u2_Display/n3998 [23]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4007 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7696  (
    .i0(\u2_Display/n3973 ),
    .i1(\u2_Display/n3998 [22]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4008 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7697  (
    .i0(\u2_Display/n3974 ),
    .i1(\u2_Display/n3998 [21]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4009 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7698  (
    .i0(\u2_Display/n3975 ),
    .i1(\u2_Display/n3998 [20]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4010 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7699  (
    .i0(\u2_Display/n3976 ),
    .i1(\u2_Display/n3998 [19]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4011 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u770  (
    .i0(\u2_Display/counta [21]),
    .i1(\u2_Display/n419 [21]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n430 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7700  (
    .i0(\u2_Display/n3977 ),
    .i1(\u2_Display/n3998 [18]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4012 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7701  (
    .i0(\u2_Display/n3978 ),
    .i1(\u2_Display/n3998 [17]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4013 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7702  (
    .i0(\u2_Display/n3979 ),
    .i1(\u2_Display/n3998 [16]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4014 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7703  (
    .i0(\u2_Display/n3980 ),
    .i1(\u2_Display/n3998 [15]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4015 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7704  (
    .i0(\u2_Display/n3981 ),
    .i1(\u2_Display/n3998 [14]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4016 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7705  (
    .i0(\u2_Display/n3982 ),
    .i1(\u2_Display/n3998 [13]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4017 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7706  (
    .i0(\u2_Display/n3983 ),
    .i1(\u2_Display/n3998 [12]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4018 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7707  (
    .i0(\u2_Display/n3984 ),
    .i1(\u2_Display/n3998 [11]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4019 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7708  (
    .i0(\u2_Display/n3985 ),
    .i1(\u2_Display/n3998 [10]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4020 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7709  (
    .i0(\u2_Display/n3986 ),
    .i1(\u2_Display/n3998 [9]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4021 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u771  (
    .i0(\u2_Display/counta [20]),
    .i1(\u2_Display/n419 [20]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n431 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7710  (
    .i0(\u2_Display/n3987 ),
    .i1(\u2_Display/n3998 [8]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4022 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7711  (
    .i0(\u2_Display/n3988 ),
    .i1(\u2_Display/n3998 [7]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4023 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7712  (
    .i0(\u2_Display/n3989 ),
    .i1(\u2_Display/n3998 [6]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4024 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7713  (
    .i0(\u2_Display/n3990 ),
    .i1(\u2_Display/n3998 [5]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4025 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7714  (
    .i0(\u2_Display/n3991 ),
    .i1(\u2_Display/n3998 [4]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4026 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7715  (
    .i0(\u2_Display/n3992 ),
    .i1(\u2_Display/n3998 [3]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4027 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7716  (
    .i0(\u2_Display/n3993 ),
    .i1(\u2_Display/n3998 [2]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4028 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7717  (
    .i0(\u2_Display/n3994 ),
    .i1(\u2_Display/n3998 [1]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4029 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7718  (
    .i0(\u2_Display/n3995 ),
    .i1(\u2_Display/n3998 [0]),
    .sel(\u2_Display/n3997 ),
    .o(\u2_Display/n4030 ));  // source/rtl/Display.v(195)
  not \u2_Display/u7719  (\u2_Display/n4032 , \u2_Display/n4031 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u772  (
    .i0(\u2_Display/counta [19]),
    .i1(\u2_Display/n419 [19]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n432 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u773  (
    .i0(\u2_Display/counta [18]),
    .i1(\u2_Display/n419 [18]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n433 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u774  (
    .i0(\u2_Display/counta [17]),
    .i1(\u2_Display/n419 [17]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n434 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u775  (
    .i0(\u2_Display/counta [16]),
    .i1(\u2_Display/n419 [16]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n435 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7752  (
    .i0(\u2_Display/n3999 ),
    .i1(\u2_Display/n4033 [31]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4034 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7753  (
    .i0(\u2_Display/n4000 ),
    .i1(\u2_Display/n4033 [30]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4035 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7754  (
    .i0(\u2_Display/n4001 ),
    .i1(\u2_Display/n4033 [29]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4036 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7755  (
    .i0(\u2_Display/n4002 ),
    .i1(\u2_Display/n4033 [28]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4037 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7756  (
    .i0(\u2_Display/n4003 ),
    .i1(\u2_Display/n4033 [27]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4038 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7757  (
    .i0(\u2_Display/n4004 ),
    .i1(\u2_Display/n4033 [26]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4039 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7758  (
    .i0(\u2_Display/n4005 ),
    .i1(\u2_Display/n4033 [25]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4040 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7759  (
    .i0(\u2_Display/n4006 ),
    .i1(\u2_Display/n4033 [24]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4041 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u776  (
    .i0(\u2_Display/counta [15]),
    .i1(\u2_Display/n419 [15]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n436 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7760  (
    .i0(\u2_Display/n4007 ),
    .i1(\u2_Display/n4033 [23]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4042 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7761  (
    .i0(\u2_Display/n4008 ),
    .i1(\u2_Display/n4033 [22]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4043 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7762  (
    .i0(\u2_Display/n4009 ),
    .i1(\u2_Display/n4033 [21]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4044 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7763  (
    .i0(\u2_Display/n4010 ),
    .i1(\u2_Display/n4033 [20]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4045 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7764  (
    .i0(\u2_Display/n4011 ),
    .i1(\u2_Display/n4033 [19]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4046 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7765  (
    .i0(\u2_Display/n4012 ),
    .i1(\u2_Display/n4033 [18]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4047 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7766  (
    .i0(\u2_Display/n4013 ),
    .i1(\u2_Display/n4033 [17]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4048 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7767  (
    .i0(\u2_Display/n4014 ),
    .i1(\u2_Display/n4033 [16]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4049 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7768  (
    .i0(\u2_Display/n4015 ),
    .i1(\u2_Display/n4033 [15]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4050 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7769  (
    .i0(\u2_Display/n4016 ),
    .i1(\u2_Display/n4033 [14]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4051 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u777  (
    .i0(\u2_Display/counta [14]),
    .i1(\u2_Display/n419 [14]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n437 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7770  (
    .i0(\u2_Display/n4017 ),
    .i1(\u2_Display/n4033 [13]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4052 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7771  (
    .i0(\u2_Display/n4018 ),
    .i1(\u2_Display/n4033 [12]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4053 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7772  (
    .i0(\u2_Display/n4019 ),
    .i1(\u2_Display/n4033 [11]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4054 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7773  (
    .i0(\u2_Display/n4020 ),
    .i1(\u2_Display/n4033 [10]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4055 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7774  (
    .i0(\u2_Display/n4021 ),
    .i1(\u2_Display/n4033 [9]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4056 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7775  (
    .i0(\u2_Display/n4022 ),
    .i1(\u2_Display/n4033 [8]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4057 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7776  (
    .i0(\u2_Display/n4023 ),
    .i1(\u2_Display/n4033 [7]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4058 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7777  (
    .i0(\u2_Display/n4024 ),
    .i1(\u2_Display/n4033 [6]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4059 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7778  (
    .i0(\u2_Display/n4025 ),
    .i1(\u2_Display/n4033 [5]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4060 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7779  (
    .i0(\u2_Display/n4026 ),
    .i1(\u2_Display/n4033 [4]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4061 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u778  (
    .i0(\u2_Display/counta [13]),
    .i1(\u2_Display/n419 [13]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n438 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7780  (
    .i0(\u2_Display/n4027 ),
    .i1(\u2_Display/n4033 [3]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4062 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7781  (
    .i0(\u2_Display/n4028 ),
    .i1(\u2_Display/n4033 [2]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4063 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7782  (
    .i0(\u2_Display/n4029 ),
    .i1(\u2_Display/n4033 [1]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4064 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7783  (
    .i0(\u2_Display/n4030 ),
    .i1(\u2_Display/n4033 [0]),
    .sel(\u2_Display/n4032 ),
    .o(\u2_Display/n4065 ));  // source/rtl/Display.v(195)
  not \u2_Display/u7784  (\u2_Display/n4067 , \u2_Display/n4066 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u779  (
    .i0(\u2_Display/counta [12]),
    .i1(\u2_Display/n419 [12]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n439 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u780  (
    .i0(\u2_Display/counta [11]),
    .i1(\u2_Display/n419 [11]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n440 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u781  (
    .i0(\u2_Display/counta [10]),
    .i1(\u2_Display/n419 [10]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n441 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7817  (
    .i0(\u2_Display/n4034 ),
    .i1(\u2_Display/n4068 [31]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4069 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7818  (
    .i0(\u2_Display/n4035 ),
    .i1(\u2_Display/n4068 [30]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4070 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7819  (
    .i0(\u2_Display/n4036 ),
    .i1(\u2_Display/n4068 [29]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4071 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u782  (
    .i0(\u2_Display/counta [9]),
    .i1(\u2_Display/n419 [9]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n442 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7820  (
    .i0(\u2_Display/n4037 ),
    .i1(\u2_Display/n4068 [28]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4072 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7821  (
    .i0(\u2_Display/n4038 ),
    .i1(\u2_Display/n4068 [27]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4073 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7822  (
    .i0(\u2_Display/n4039 ),
    .i1(\u2_Display/n4068 [26]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4074 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7823  (
    .i0(\u2_Display/n4040 ),
    .i1(\u2_Display/n4068 [25]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4075 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7824  (
    .i0(\u2_Display/n4041 ),
    .i1(\u2_Display/n4068 [24]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4076 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7825  (
    .i0(\u2_Display/n4042 ),
    .i1(\u2_Display/n4068 [23]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4077 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7826  (
    .i0(\u2_Display/n4043 ),
    .i1(\u2_Display/n4068 [22]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4078 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7827  (
    .i0(\u2_Display/n4044 ),
    .i1(\u2_Display/n4068 [21]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4079 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7828  (
    .i0(\u2_Display/n4045 ),
    .i1(\u2_Display/n4068 [20]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4080 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7829  (
    .i0(\u2_Display/n4046 ),
    .i1(\u2_Display/n4068 [19]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4081 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u783  (
    .i0(\u2_Display/counta [8]),
    .i1(\u2_Display/n419 [8]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n443 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7830  (
    .i0(\u2_Display/n4047 ),
    .i1(\u2_Display/n4068 [18]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4082 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7831  (
    .i0(\u2_Display/n4048 ),
    .i1(\u2_Display/n4068 [17]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4083 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7832  (
    .i0(\u2_Display/n4049 ),
    .i1(\u2_Display/n4068 [16]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4084 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7833  (
    .i0(\u2_Display/n4050 ),
    .i1(\u2_Display/n4068 [15]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4085 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7834  (
    .i0(\u2_Display/n4051 ),
    .i1(\u2_Display/n4068 [14]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4086 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7835  (
    .i0(\u2_Display/n4052 ),
    .i1(\u2_Display/n4068 [13]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4087 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7836  (
    .i0(\u2_Display/n4053 ),
    .i1(\u2_Display/n4068 [12]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4088 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7837  (
    .i0(\u2_Display/n4054 ),
    .i1(\u2_Display/n4068 [11]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4089 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7838  (
    .i0(\u2_Display/n4055 ),
    .i1(\u2_Display/n4068 [10]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4090 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7839  (
    .i0(\u2_Display/n4056 ),
    .i1(\u2_Display/n4068 [9]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4091 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u784  (
    .i0(\u2_Display/counta [7]),
    .i1(\u2_Display/n419 [7]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n444 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7840  (
    .i0(\u2_Display/n4057 ),
    .i1(\u2_Display/n4068 [8]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4092 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7841  (
    .i0(\u2_Display/n4058 ),
    .i1(\u2_Display/n4068 [7]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4093 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7842  (
    .i0(\u2_Display/n4059 ),
    .i1(\u2_Display/n4068 [6]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4094 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7843  (
    .i0(\u2_Display/n4060 ),
    .i1(\u2_Display/n4068 [5]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4095 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7844  (
    .i0(\u2_Display/n4061 ),
    .i1(\u2_Display/n4068 [4]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4096 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7845  (
    .i0(\u2_Display/n4062 ),
    .i1(\u2_Display/n4068 [3]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4097 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7846  (
    .i0(\u2_Display/n4063 ),
    .i1(\u2_Display/n4068 [2]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4098 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7847  (
    .i0(\u2_Display/n4064 ),
    .i1(\u2_Display/n4068 [1]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4099 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7848  (
    .i0(\u2_Display/n4065 ),
    .i1(\u2_Display/n4068 [0]),
    .sel(\u2_Display/n4067 ),
    .o(\u2_Display/n4100 ));  // source/rtl/Display.v(195)
  not \u2_Display/u7849  (\u2_Display/n4102 , \u2_Display/n4101 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u785  (
    .i0(\u2_Display/counta [6]),
    .i1(\u2_Display/n419 [6]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n445 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u786  (
    .i0(\u2_Display/counta [5]),
    .i1(\u2_Display/n419 [5]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n446 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u787  (
    .i0(\u2_Display/counta [4]),
    .i1(\u2_Display/n419 [4]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n447 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u788  (
    .i0(\u2_Display/counta [3]),
    .i1(\u2_Display/n419 [3]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n448 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7882  (
    .i0(\u2_Display/n4069 ),
    .i1(\u2_Display/n4103 [31]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4104 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7883  (
    .i0(\u2_Display/n4070 ),
    .i1(\u2_Display/n4103 [30]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4105 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7884  (
    .i0(\u2_Display/n4071 ),
    .i1(\u2_Display/n4103 [29]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4106 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7885  (
    .i0(\u2_Display/n4072 ),
    .i1(\u2_Display/n4103 [28]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4107 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7886  (
    .i0(\u2_Display/n4073 ),
    .i1(\u2_Display/n4103 [27]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4108 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7887  (
    .i0(\u2_Display/n4074 ),
    .i1(\u2_Display/n4103 [26]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4109 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7888  (
    .i0(\u2_Display/n4075 ),
    .i1(\u2_Display/n4103 [25]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4110 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7889  (
    .i0(\u2_Display/n4076 ),
    .i1(\u2_Display/n4103 [24]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4111 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u789  (
    .i0(\u2_Display/counta [2]),
    .i1(\u2_Display/n419 [2]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n449 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7890  (
    .i0(\u2_Display/n4077 ),
    .i1(\u2_Display/n4103 [23]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4112 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7891  (
    .i0(\u2_Display/n4078 ),
    .i1(\u2_Display/n4103 [22]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4113 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7892  (
    .i0(\u2_Display/n4079 ),
    .i1(\u2_Display/n4103 [21]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4114 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7893  (
    .i0(\u2_Display/n4080 ),
    .i1(\u2_Display/n4103 [20]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4115 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7894  (
    .i0(\u2_Display/n4081 ),
    .i1(\u2_Display/n4103 [19]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4116 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7895  (
    .i0(\u2_Display/n4082 ),
    .i1(\u2_Display/n4103 [18]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4117 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7896  (
    .i0(\u2_Display/n4083 ),
    .i1(\u2_Display/n4103 [17]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4118 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7897  (
    .i0(\u2_Display/n4084 ),
    .i1(\u2_Display/n4103 [16]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4119 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7898  (
    .i0(\u2_Display/n4085 ),
    .i1(\u2_Display/n4103 [15]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4120 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7899  (
    .i0(\u2_Display/n4086 ),
    .i1(\u2_Display/n4103 [14]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4121 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u790  (
    .i0(\u2_Display/counta [1]),
    .i1(\u2_Display/n419 [1]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n450 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7900  (
    .i0(\u2_Display/n4087 ),
    .i1(\u2_Display/n4103 [13]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4122 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7901  (
    .i0(\u2_Display/n4088 ),
    .i1(\u2_Display/n4103 [12]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4123 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7902  (
    .i0(\u2_Display/n4089 ),
    .i1(\u2_Display/n4103 [11]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4124 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7903  (
    .i0(\u2_Display/n4090 ),
    .i1(\u2_Display/n4103 [10]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4125 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7904  (
    .i0(\u2_Display/n4091 ),
    .i1(\u2_Display/n4103 [9]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4126 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7905  (
    .i0(\u2_Display/n4092 ),
    .i1(\u2_Display/n4103 [8]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4127 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7906  (
    .i0(\u2_Display/n4093 ),
    .i1(\u2_Display/n4103 [7]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4128 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7907  (
    .i0(\u2_Display/n4094 ),
    .i1(\u2_Display/n4103 [6]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4129 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7908  (
    .i0(\u2_Display/n4095 ),
    .i1(\u2_Display/n4103 [5]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4130 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7909  (
    .i0(\u2_Display/n4096 ),
    .i1(\u2_Display/n4103 [4]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4131 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u791  (
    .i0(\u2_Display/counta [0]),
    .i1(\u2_Display/n419 [0]),
    .sel(\u2_Display/n418 ),
    .o(\u2_Display/n451 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7910  (
    .i0(\u2_Display/n4097 ),
    .i1(\u2_Display/n4103 [3]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4132 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7911  (
    .i0(\u2_Display/n4098 ),
    .i1(\u2_Display/n4103 [2]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4133 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7912  (
    .i0(\u2_Display/n4099 ),
    .i1(\u2_Display/n4103 [1]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4134 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7913  (
    .i0(\u2_Display/n4100 ),
    .i1(\u2_Display/n4103 [0]),
    .sel(\u2_Display/n4102 ),
    .o(\u2_Display/n4135 ));  // source/rtl/Display.v(195)
  not \u2_Display/u7914  (\u2_Display/n4137 , \u2_Display/n4136 );  // source/rtl/Display.v(195)
  not \u2_Display/u792  (\u2_Display/n453 , \u2_Display/n452 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u7947  (
    .i0(\u2_Display/n4104 ),
    .i1(\u2_Display/n4138 [31]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4139 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7948  (
    .i0(\u2_Display/n4105 ),
    .i1(\u2_Display/n4138 [30]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4140 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7949  (
    .i0(\u2_Display/n4106 ),
    .i1(\u2_Display/n4138 [29]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4141 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7950  (
    .i0(\u2_Display/n4107 ),
    .i1(\u2_Display/n4138 [28]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4142 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7951  (
    .i0(\u2_Display/n4108 ),
    .i1(\u2_Display/n4138 [27]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4143 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7952  (
    .i0(\u2_Display/n4109 ),
    .i1(\u2_Display/n4138 [26]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4144 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7953  (
    .i0(\u2_Display/n4110 ),
    .i1(\u2_Display/n4138 [25]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4145 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7954  (
    .i0(\u2_Display/n4111 ),
    .i1(\u2_Display/n4138 [24]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4146 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7955  (
    .i0(\u2_Display/n4112 ),
    .i1(\u2_Display/n4138 [23]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4147 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7956  (
    .i0(\u2_Display/n4113 ),
    .i1(\u2_Display/n4138 [22]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4148 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7957  (
    .i0(\u2_Display/n4114 ),
    .i1(\u2_Display/n4138 [21]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4149 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7958  (
    .i0(\u2_Display/n4115 ),
    .i1(\u2_Display/n4138 [20]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4150 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7959  (
    .i0(\u2_Display/n4116 ),
    .i1(\u2_Display/n4138 [19]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4151 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7960  (
    .i0(\u2_Display/n4117 ),
    .i1(\u2_Display/n4138 [18]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4152 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7961  (
    .i0(\u2_Display/n4118 ),
    .i1(\u2_Display/n4138 [17]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4153 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7962  (
    .i0(\u2_Display/n4119 ),
    .i1(\u2_Display/n4138 [16]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4154 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7963  (
    .i0(\u2_Display/n4120 ),
    .i1(\u2_Display/n4138 [15]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4155 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7964  (
    .i0(\u2_Display/n4121 ),
    .i1(\u2_Display/n4138 [14]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4156 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7965  (
    .i0(\u2_Display/n4122 ),
    .i1(\u2_Display/n4138 [13]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4157 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7966  (
    .i0(\u2_Display/n4123 ),
    .i1(\u2_Display/n4138 [12]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4158 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7967  (
    .i0(\u2_Display/n4124 ),
    .i1(\u2_Display/n4138 [11]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4159 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7968  (
    .i0(\u2_Display/n4125 ),
    .i1(\u2_Display/n4138 [10]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4160 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7969  (
    .i0(\u2_Display/n4126 ),
    .i1(\u2_Display/n4138 [9]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4161 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7970  (
    .i0(\u2_Display/n4127 ),
    .i1(\u2_Display/n4138 [8]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4162 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7971  (
    .i0(\u2_Display/n4128 ),
    .i1(\u2_Display/n4138 [7]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4163 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7972  (
    .i0(\u2_Display/n4129 ),
    .i1(\u2_Display/n4138 [6]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4164 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7973  (
    .i0(\u2_Display/n4130 ),
    .i1(\u2_Display/n4138 [5]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4165 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7974  (
    .i0(\u2_Display/n4131 ),
    .i1(\u2_Display/n4138 [4]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4166 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7975  (
    .i0(\u2_Display/n4132 ),
    .i1(\u2_Display/n4138 [3]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4167 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7976  (
    .i0(\u2_Display/n4133 ),
    .i1(\u2_Display/n4138 [2]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4168 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7977  (
    .i0(\u2_Display/n4134 ),
    .i1(\u2_Display/n4138 [1]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4169 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u7978  (
    .i0(\u2_Display/n4135 ),
    .i1(\u2_Display/n4138 [0]),
    .sel(\u2_Display/n4137 ),
    .o(\u2_Display/n4170 ));  // source/rtl/Display.v(195)
  not \u2_Display/u7979  (\u2_Display/n4172 , \u2_Display/n4171 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8012  (
    .i0(\u2_Display/n4139 ),
    .i1(\u2_Display/n4173 [31]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4174 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8013  (
    .i0(\u2_Display/n4140 ),
    .i1(\u2_Display/n4173 [30]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4175 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8014  (
    .i0(\u2_Display/n4141 ),
    .i1(\u2_Display/n4173 [29]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4176 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8015  (
    .i0(\u2_Display/n4142 ),
    .i1(\u2_Display/n4173 [28]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4177 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8016  (
    .i0(\u2_Display/n4143 ),
    .i1(\u2_Display/n4173 [27]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4178 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8017  (
    .i0(\u2_Display/n4144 ),
    .i1(\u2_Display/n4173 [26]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4179 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8018  (
    .i0(\u2_Display/n4145 ),
    .i1(\u2_Display/n4173 [25]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4180 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8019  (
    .i0(\u2_Display/n4146 ),
    .i1(\u2_Display/n4173 [24]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4181 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8020  (
    .i0(\u2_Display/n4147 ),
    .i1(\u2_Display/n4173 [23]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4182 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8021  (
    .i0(\u2_Display/n4148 ),
    .i1(\u2_Display/n4173 [22]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4183 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8022  (
    .i0(\u2_Display/n4149 ),
    .i1(\u2_Display/n4173 [21]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4184 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8023  (
    .i0(\u2_Display/n4150 ),
    .i1(\u2_Display/n4173 [20]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4185 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8024  (
    .i0(\u2_Display/n4151 ),
    .i1(\u2_Display/n4173 [19]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4186 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8025  (
    .i0(\u2_Display/n4152 ),
    .i1(\u2_Display/n4173 [18]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4187 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8026  (
    .i0(\u2_Display/n4153 ),
    .i1(\u2_Display/n4173 [17]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4188 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8027  (
    .i0(\u2_Display/n4154 ),
    .i1(\u2_Display/n4173 [16]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4189 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8028  (
    .i0(\u2_Display/n4155 ),
    .i1(\u2_Display/n4173 [15]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4190 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8029  (
    .i0(\u2_Display/n4156 ),
    .i1(\u2_Display/n4173 [14]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4191 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8030  (
    .i0(\u2_Display/n4157 ),
    .i1(\u2_Display/n4173 [13]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4192 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8031  (
    .i0(\u2_Display/n4158 ),
    .i1(\u2_Display/n4173 [12]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4193 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8032  (
    .i0(\u2_Display/n4159 ),
    .i1(\u2_Display/n4173 [11]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4194 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8033  (
    .i0(\u2_Display/n4160 ),
    .i1(\u2_Display/n4173 [10]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4195 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8034  (
    .i0(\u2_Display/n4161 ),
    .i1(\u2_Display/n4173 [9]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4196 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8035  (
    .i0(\u2_Display/n4162 ),
    .i1(\u2_Display/n4173 [8]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4197 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8036  (
    .i0(\u2_Display/n4163 ),
    .i1(\u2_Display/n4173 [7]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4198 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8037  (
    .i0(\u2_Display/n4164 ),
    .i1(\u2_Display/n4173 [6]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4199 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8038  (
    .i0(\u2_Display/n4165 ),
    .i1(\u2_Display/n4173 [5]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4200 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8039  (
    .i0(\u2_Display/n4166 ),
    .i1(\u2_Display/n4173 [4]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4201 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8040  (
    .i0(\u2_Display/n4167 ),
    .i1(\u2_Display/n4173 [3]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4202 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8041  (
    .i0(\u2_Display/n4168 ),
    .i1(\u2_Display/n4173 [2]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4203 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8042  (
    .i0(\u2_Display/n4169 ),
    .i1(\u2_Display/n4173 [1]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4204 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8043  (
    .i0(\u2_Display/n4170 ),
    .i1(\u2_Display/n4173 [0]),
    .sel(\u2_Display/n4172 ),
    .o(\u2_Display/n4205 ));  // source/rtl/Display.v(195)
  not \u2_Display/u8044  (\u2_Display/n4207 , \u2_Display/n4206 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8077  (
    .i0(\u2_Display/n4174 ),
    .i1(\u2_Display/n4208 [31]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4209 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8078  (
    .i0(\u2_Display/n4175 ),
    .i1(\u2_Display/n4208 [30]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4210 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8079  (
    .i0(\u2_Display/n4176 ),
    .i1(\u2_Display/n4208 [29]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4211 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8080  (
    .i0(\u2_Display/n4177 ),
    .i1(\u2_Display/n4208 [28]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4212 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8081  (
    .i0(\u2_Display/n4178 ),
    .i1(\u2_Display/n4208 [27]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4213 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8082  (
    .i0(\u2_Display/n4179 ),
    .i1(\u2_Display/n4208 [26]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4214 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8083  (
    .i0(\u2_Display/n4180 ),
    .i1(\u2_Display/n4208 [25]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4215 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8084  (
    .i0(\u2_Display/n4181 ),
    .i1(\u2_Display/n4208 [24]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4216 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8085  (
    .i0(\u2_Display/n4182 ),
    .i1(\u2_Display/n4208 [23]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4217 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8086  (
    .i0(\u2_Display/n4183 ),
    .i1(\u2_Display/n4208 [22]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4218 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8087  (
    .i0(\u2_Display/n4184 ),
    .i1(\u2_Display/n4208 [21]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4219 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8088  (
    .i0(\u2_Display/n4185 ),
    .i1(\u2_Display/n4208 [20]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4220 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8089  (
    .i0(\u2_Display/n4186 ),
    .i1(\u2_Display/n4208 [19]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4221 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8090  (
    .i0(\u2_Display/n4187 ),
    .i1(\u2_Display/n4208 [18]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4222 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8091  (
    .i0(\u2_Display/n4188 ),
    .i1(\u2_Display/n4208 [17]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4223 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8092  (
    .i0(\u2_Display/n4189 ),
    .i1(\u2_Display/n4208 [16]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4224 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8093  (
    .i0(\u2_Display/n4190 ),
    .i1(\u2_Display/n4208 [15]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4225 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8094  (
    .i0(\u2_Display/n4191 ),
    .i1(\u2_Display/n4208 [14]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4226 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8095  (
    .i0(\u2_Display/n4192 ),
    .i1(\u2_Display/n4208 [13]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4227 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8096  (
    .i0(\u2_Display/n4193 ),
    .i1(\u2_Display/n4208 [12]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4228 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8097  (
    .i0(\u2_Display/n4194 ),
    .i1(\u2_Display/n4208 [11]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4229 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8098  (
    .i0(\u2_Display/n4195 ),
    .i1(\u2_Display/n4208 [10]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4230 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8099  (
    .i0(\u2_Display/n4196 ),
    .i1(\u2_Display/n4208 [9]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4231 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8100  (
    .i0(\u2_Display/n4197 ),
    .i1(\u2_Display/n4208 [8]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4232 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8101  (
    .i0(\u2_Display/n4198 ),
    .i1(\u2_Display/n4208 [7]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4233 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8102  (
    .i0(\u2_Display/n4199 ),
    .i1(\u2_Display/n4208 [6]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4234 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8103  (
    .i0(\u2_Display/n4200 ),
    .i1(\u2_Display/n4208 [5]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4235 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8104  (
    .i0(\u2_Display/n4201 ),
    .i1(\u2_Display/n4208 [4]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4236 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8105  (
    .i0(\u2_Display/n4202 ),
    .i1(\u2_Display/n4208 [3]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4237 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8106  (
    .i0(\u2_Display/n4203 ),
    .i1(\u2_Display/n4208 [2]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4238 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8107  (
    .i0(\u2_Display/n4204 ),
    .i1(\u2_Display/n4208 [1]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4239 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8108  (
    .i0(\u2_Display/n4205 ),
    .i1(\u2_Display/n4208 [0]),
    .sel(\u2_Display/n4207 ),
    .o(\u2_Display/n4240 ));  // source/rtl/Display.v(195)
  not \u2_Display/u8109  (\u2_Display/n4242 , \u2_Display/n4241 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8142  (
    .i0(\u2_Display/n4209 ),
    .i1(\u2_Display/n4243 [31]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4244 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8143  (
    .i0(\u2_Display/n4210 ),
    .i1(\u2_Display/n4243 [30]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4245 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8144  (
    .i0(\u2_Display/n4211 ),
    .i1(\u2_Display/n4243 [29]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4246 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8145  (
    .i0(\u2_Display/n4212 ),
    .i1(\u2_Display/n4243 [28]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4247 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8146  (
    .i0(\u2_Display/n4213 ),
    .i1(\u2_Display/n4243 [27]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4248 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8147  (
    .i0(\u2_Display/n4214 ),
    .i1(\u2_Display/n4243 [26]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4249 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8148  (
    .i0(\u2_Display/n4215 ),
    .i1(\u2_Display/n4243 [25]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4250 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8149  (
    .i0(\u2_Display/n4216 ),
    .i1(\u2_Display/n4243 [24]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4251 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8150  (
    .i0(\u2_Display/n4217 ),
    .i1(\u2_Display/n4243 [23]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4252 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8151  (
    .i0(\u2_Display/n4218 ),
    .i1(\u2_Display/n4243 [22]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4253 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8152  (
    .i0(\u2_Display/n4219 ),
    .i1(\u2_Display/n4243 [21]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4254 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8153  (
    .i0(\u2_Display/n4220 ),
    .i1(\u2_Display/n4243 [20]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4255 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8154  (
    .i0(\u2_Display/n4221 ),
    .i1(\u2_Display/n4243 [19]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4256 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8155  (
    .i0(\u2_Display/n4222 ),
    .i1(\u2_Display/n4243 [18]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4257 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8156  (
    .i0(\u2_Display/n4223 ),
    .i1(\u2_Display/n4243 [17]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4258 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8157  (
    .i0(\u2_Display/n4224 ),
    .i1(\u2_Display/n4243 [16]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4259 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8158  (
    .i0(\u2_Display/n4225 ),
    .i1(\u2_Display/n4243 [15]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4260 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8159  (
    .i0(\u2_Display/n4226 ),
    .i1(\u2_Display/n4243 [14]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4261 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8160  (
    .i0(\u2_Display/n4227 ),
    .i1(\u2_Display/n4243 [13]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4262 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8161  (
    .i0(\u2_Display/n4228 ),
    .i1(\u2_Display/n4243 [12]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4263 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8162  (
    .i0(\u2_Display/n4229 ),
    .i1(\u2_Display/n4243 [11]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4264 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8163  (
    .i0(\u2_Display/n4230 ),
    .i1(\u2_Display/n4243 [10]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4265 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8164  (
    .i0(\u2_Display/n4231 ),
    .i1(\u2_Display/n4243 [9]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4266 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8165  (
    .i0(\u2_Display/n4232 ),
    .i1(\u2_Display/n4243 [8]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4267 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8166  (
    .i0(\u2_Display/n4233 ),
    .i1(\u2_Display/n4243 [7]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4268 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8167  (
    .i0(\u2_Display/n4234 ),
    .i1(\u2_Display/n4243 [6]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4269 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8168  (
    .i0(\u2_Display/n4235 ),
    .i1(\u2_Display/n4243 [5]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4270 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8169  (
    .i0(\u2_Display/n4236 ),
    .i1(\u2_Display/n4243 [4]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4271 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8170  (
    .i0(\u2_Display/n4237 ),
    .i1(\u2_Display/n4243 [3]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4272 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8171  (
    .i0(\u2_Display/n4238 ),
    .i1(\u2_Display/n4243 [2]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4273 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8172  (
    .i0(\u2_Display/n4239 ),
    .i1(\u2_Display/n4243 [1]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4274 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8173  (
    .i0(\u2_Display/n4240 ),
    .i1(\u2_Display/n4243 [0]),
    .sel(\u2_Display/n4242 ),
    .o(\u2_Display/n4275 ));  // source/rtl/Display.v(195)
  not \u2_Display/u8174  (\u2_Display/n4277 , \u2_Display/n4276 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8207  (
    .i0(\u2_Display/n4244 ),
    .i1(\u2_Display/n4278 [31]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4279 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8208  (
    .i0(\u2_Display/n4245 ),
    .i1(\u2_Display/n4278 [30]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4280 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8209  (
    .i0(\u2_Display/n4246 ),
    .i1(\u2_Display/n4278 [29]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4281 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8210  (
    .i0(\u2_Display/n4247 ),
    .i1(\u2_Display/n4278 [28]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4282 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8211  (
    .i0(\u2_Display/n4248 ),
    .i1(\u2_Display/n4278 [27]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4283 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8212  (
    .i0(\u2_Display/n4249 ),
    .i1(\u2_Display/n4278 [26]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4284 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8213  (
    .i0(\u2_Display/n4250 ),
    .i1(\u2_Display/n4278 [25]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4285 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8214  (
    .i0(\u2_Display/n4251 ),
    .i1(\u2_Display/n4278 [24]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4286 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8215  (
    .i0(\u2_Display/n4252 ),
    .i1(\u2_Display/n4278 [23]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4287 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8216  (
    .i0(\u2_Display/n4253 ),
    .i1(\u2_Display/n4278 [22]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4288 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8217  (
    .i0(\u2_Display/n4254 ),
    .i1(\u2_Display/n4278 [21]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4289 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8218  (
    .i0(\u2_Display/n4255 ),
    .i1(\u2_Display/n4278 [20]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4290 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8219  (
    .i0(\u2_Display/n4256 ),
    .i1(\u2_Display/n4278 [19]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4291 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8220  (
    .i0(\u2_Display/n4257 ),
    .i1(\u2_Display/n4278 [18]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4292 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8221  (
    .i0(\u2_Display/n4258 ),
    .i1(\u2_Display/n4278 [17]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4293 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8222  (
    .i0(\u2_Display/n4259 ),
    .i1(\u2_Display/n4278 [16]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4294 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8223  (
    .i0(\u2_Display/n4260 ),
    .i1(\u2_Display/n4278 [15]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4295 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8224  (
    .i0(\u2_Display/n4261 ),
    .i1(\u2_Display/n4278 [14]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4296 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8225  (
    .i0(\u2_Display/n4262 ),
    .i1(\u2_Display/n4278 [13]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4297 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8226  (
    .i0(\u2_Display/n4263 ),
    .i1(\u2_Display/n4278 [12]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4298 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8227  (
    .i0(\u2_Display/n4264 ),
    .i1(\u2_Display/n4278 [11]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4299 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8228  (
    .i0(\u2_Display/n4265 ),
    .i1(\u2_Display/n4278 [10]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4300 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8229  (
    .i0(\u2_Display/n4266 ),
    .i1(\u2_Display/n4278 [9]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4301 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8230  (
    .i0(\u2_Display/n4267 ),
    .i1(\u2_Display/n4278 [8]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4302 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8231  (
    .i0(\u2_Display/n4268 ),
    .i1(\u2_Display/n4278 [7]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4303 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8232  (
    .i0(\u2_Display/n4269 ),
    .i1(\u2_Display/n4278 [6]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4304 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8233  (
    .i0(\u2_Display/n4270 ),
    .i1(\u2_Display/n4278 [5]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4305 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8234  (
    .i0(\u2_Display/n4271 ),
    .i1(\u2_Display/n4278 [4]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4306 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8235  (
    .i0(\u2_Display/n4272 ),
    .i1(\u2_Display/n4278 [3]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4307 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8236  (
    .i0(\u2_Display/n4273 ),
    .i1(\u2_Display/n4278 [2]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4308 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8237  (
    .i0(\u2_Display/n4274 ),
    .i1(\u2_Display/n4278 [1]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4309 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8238  (
    .i0(\u2_Display/n4275 ),
    .i1(\u2_Display/n4278 [0]),
    .sel(\u2_Display/n4277 ),
    .o(\u2_Display/n4310 ));  // source/rtl/Display.v(195)
  not \u2_Display/u8239  (\u2_Display/n4312 , \u2_Display/n4311 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u825  (
    .i0(\u2_Display/n420 ),
    .i1(\u2_Display/n454 [31]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n455 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u826  (
    .i0(\u2_Display/n421 ),
    .i1(\u2_Display/n454 [30]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n456 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u827  (
    .i0(\u2_Display/n422 ),
    .i1(\u2_Display/n454 [29]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n457 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8272  (
    .i0(\u2_Display/n4279 ),
    .i1(\u2_Display/n4313 [31]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4314 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8273  (
    .i0(\u2_Display/n4280 ),
    .i1(\u2_Display/n4313 [30]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4315 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8274  (
    .i0(\u2_Display/n4281 ),
    .i1(\u2_Display/n4313 [29]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4316 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8275  (
    .i0(\u2_Display/n4282 ),
    .i1(\u2_Display/n4313 [28]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4317 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8276  (
    .i0(\u2_Display/n4283 ),
    .i1(\u2_Display/n4313 [27]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4318 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8277  (
    .i0(\u2_Display/n4284 ),
    .i1(\u2_Display/n4313 [26]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4319 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8278  (
    .i0(\u2_Display/n4285 ),
    .i1(\u2_Display/n4313 [25]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4320 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8279  (
    .i0(\u2_Display/n4286 ),
    .i1(\u2_Display/n4313 [24]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4321 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u828  (
    .i0(\u2_Display/n423 ),
    .i1(\u2_Display/n454 [28]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n458 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8280  (
    .i0(\u2_Display/n4287 ),
    .i1(\u2_Display/n4313 [23]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4322 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8281  (
    .i0(\u2_Display/n4288 ),
    .i1(\u2_Display/n4313 [22]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4323 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8282  (
    .i0(\u2_Display/n4289 ),
    .i1(\u2_Display/n4313 [21]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4324 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8283  (
    .i0(\u2_Display/n4290 ),
    .i1(\u2_Display/n4313 [20]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4325 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8284  (
    .i0(\u2_Display/n4291 ),
    .i1(\u2_Display/n4313 [19]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4326 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8285  (
    .i0(\u2_Display/n4292 ),
    .i1(\u2_Display/n4313 [18]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4327 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8286  (
    .i0(\u2_Display/n4293 ),
    .i1(\u2_Display/n4313 [17]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4328 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8287  (
    .i0(\u2_Display/n4294 ),
    .i1(\u2_Display/n4313 [16]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4329 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8288  (
    .i0(\u2_Display/n4295 ),
    .i1(\u2_Display/n4313 [15]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4330 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8289  (
    .i0(\u2_Display/n4296 ),
    .i1(\u2_Display/n4313 [14]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4331 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u829  (
    .i0(\u2_Display/n424 ),
    .i1(\u2_Display/n454 [27]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n459 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8290  (
    .i0(\u2_Display/n4297 ),
    .i1(\u2_Display/n4313 [13]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4332 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8291  (
    .i0(\u2_Display/n4298 ),
    .i1(\u2_Display/n4313 [12]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4333 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8292  (
    .i0(\u2_Display/n4299 ),
    .i1(\u2_Display/n4313 [11]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4334 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8293  (
    .i0(\u2_Display/n4300 ),
    .i1(\u2_Display/n4313 [10]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4335 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8294  (
    .i0(\u2_Display/n4301 ),
    .i1(\u2_Display/n4313 [9]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4336 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8295  (
    .i0(\u2_Display/n4302 ),
    .i1(\u2_Display/n4313 [8]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4337 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8296  (
    .i0(\u2_Display/n4303 ),
    .i1(\u2_Display/n4313 [7]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4338 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8297  (
    .i0(\u2_Display/n4304 ),
    .i1(\u2_Display/n4313 [6]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4339 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8298  (
    .i0(\u2_Display/n4305 ),
    .i1(\u2_Display/n4313 [5]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4340 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8299  (
    .i0(\u2_Display/n4306 ),
    .i1(\u2_Display/n4313 [4]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4341 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u830  (
    .i0(\u2_Display/n425 ),
    .i1(\u2_Display/n454 [26]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n460 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8300  (
    .i0(\u2_Display/n4307 ),
    .i1(\u2_Display/n4313 [3]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4342 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8301  (
    .i0(\u2_Display/n4308 ),
    .i1(\u2_Display/n4313 [2]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4343 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8302  (
    .i0(\u2_Display/n4309 ),
    .i1(\u2_Display/n4313 [1]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4344 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8303  (
    .i0(\u2_Display/n4310 ),
    .i1(\u2_Display/n4313 [0]),
    .sel(\u2_Display/n4312 ),
    .o(\u2_Display/n4345 ));  // source/rtl/Display.v(195)
  not \u2_Display/u8304  (\u2_Display/n4347 , \u2_Display/n4346 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u831  (
    .i0(\u2_Display/n426 ),
    .i1(\u2_Display/n454 [25]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n461 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u832  (
    .i0(\u2_Display/n427 ),
    .i1(\u2_Display/n454 [24]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n462 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u833  (
    .i0(\u2_Display/n428 ),
    .i1(\u2_Display/n454 [23]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n463 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8337  (
    .i0(\u2_Display/n4314 ),
    .i1(\u2_Display/n4348 [31]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4349 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8338  (
    .i0(\u2_Display/n4315 ),
    .i1(\u2_Display/n4348 [30]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4350 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8339  (
    .i0(\u2_Display/n4316 ),
    .i1(\u2_Display/n4348 [29]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4351 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u834  (
    .i0(\u2_Display/n429 ),
    .i1(\u2_Display/n454 [22]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n464 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8340  (
    .i0(\u2_Display/n4317 ),
    .i1(\u2_Display/n4348 [28]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4352 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8341  (
    .i0(\u2_Display/n4318 ),
    .i1(\u2_Display/n4348 [27]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4353 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8342  (
    .i0(\u2_Display/n4319 ),
    .i1(\u2_Display/n4348 [26]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4354 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8343  (
    .i0(\u2_Display/n4320 ),
    .i1(\u2_Display/n4348 [25]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4355 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8344  (
    .i0(\u2_Display/n4321 ),
    .i1(\u2_Display/n4348 [24]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4356 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8345  (
    .i0(\u2_Display/n4322 ),
    .i1(\u2_Display/n4348 [23]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4357 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8346  (
    .i0(\u2_Display/n4323 ),
    .i1(\u2_Display/n4348 [22]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4358 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8347  (
    .i0(\u2_Display/n4324 ),
    .i1(\u2_Display/n4348 [21]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4359 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8348  (
    .i0(\u2_Display/n4325 ),
    .i1(\u2_Display/n4348 [20]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4360 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8349  (
    .i0(\u2_Display/n4326 ),
    .i1(\u2_Display/n4348 [19]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4361 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u835  (
    .i0(\u2_Display/n430 ),
    .i1(\u2_Display/n454 [21]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n465 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8350  (
    .i0(\u2_Display/n4327 ),
    .i1(\u2_Display/n4348 [18]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4362 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8351  (
    .i0(\u2_Display/n4328 ),
    .i1(\u2_Display/n4348 [17]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4363 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8352  (
    .i0(\u2_Display/n4329 ),
    .i1(\u2_Display/n4348 [16]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4364 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8353  (
    .i0(\u2_Display/n4330 ),
    .i1(\u2_Display/n4348 [15]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4365 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8354  (
    .i0(\u2_Display/n4331 ),
    .i1(\u2_Display/n4348 [14]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4366 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8355  (
    .i0(\u2_Display/n4332 ),
    .i1(\u2_Display/n4348 [13]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4367 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8356  (
    .i0(\u2_Display/n4333 ),
    .i1(\u2_Display/n4348 [12]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4368 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8357  (
    .i0(\u2_Display/n4334 ),
    .i1(\u2_Display/n4348 [11]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4369 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8358  (
    .i0(\u2_Display/n4335 ),
    .i1(\u2_Display/n4348 [10]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4370 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8359  (
    .i0(\u2_Display/n4336 ),
    .i1(\u2_Display/n4348 [9]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4371 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u836  (
    .i0(\u2_Display/n431 ),
    .i1(\u2_Display/n454 [20]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n466 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8360  (
    .i0(\u2_Display/n4337 ),
    .i1(\u2_Display/n4348 [8]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4372 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8361  (
    .i0(\u2_Display/n4338 ),
    .i1(\u2_Display/n4348 [7]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4373 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8362  (
    .i0(\u2_Display/n4339 ),
    .i1(\u2_Display/n4348 [6]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4374 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8363  (
    .i0(\u2_Display/n4340 ),
    .i1(\u2_Display/n4348 [5]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4375 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8364  (
    .i0(\u2_Display/n4341 ),
    .i1(\u2_Display/n4348 [4]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4376 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8365  (
    .i0(\u2_Display/n4342 ),
    .i1(\u2_Display/n4348 [3]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4377 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8366  (
    .i0(\u2_Display/n4343 ),
    .i1(\u2_Display/n4348 [2]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4378 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8367  (
    .i0(\u2_Display/n4344 ),
    .i1(\u2_Display/n4348 [1]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4379 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8368  (
    .i0(\u2_Display/n4345 ),
    .i1(\u2_Display/n4348 [0]),
    .sel(\u2_Display/n4347 ),
    .o(\u2_Display/n4380 ));  // source/rtl/Display.v(195)
  not \u2_Display/u8369  (\u2_Display/n4382 , \u2_Display/n4381 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u837  (
    .i0(\u2_Display/n432 ),
    .i1(\u2_Display/n454 [19]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n467 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u838  (
    .i0(\u2_Display/n433 ),
    .i1(\u2_Display/n454 [18]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n468 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u839  (
    .i0(\u2_Display/n434 ),
    .i1(\u2_Display/n454 [17]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n469 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u840  (
    .i0(\u2_Display/n435 ),
    .i1(\u2_Display/n454 [16]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n470 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8402  (
    .i0(\u2_Display/n4349 ),
    .i1(\u2_Display/n4383 [31]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4384 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8403  (
    .i0(\u2_Display/n4350 ),
    .i1(\u2_Display/n4383 [30]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4385 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8404  (
    .i0(\u2_Display/n4351 ),
    .i1(\u2_Display/n4383 [29]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4386 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8405  (
    .i0(\u2_Display/n4352 ),
    .i1(\u2_Display/n4383 [28]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4387 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8406  (
    .i0(\u2_Display/n4353 ),
    .i1(\u2_Display/n4383 [27]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4388 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8407  (
    .i0(\u2_Display/n4354 ),
    .i1(\u2_Display/n4383 [26]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4389 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8408  (
    .i0(\u2_Display/n4355 ),
    .i1(\u2_Display/n4383 [25]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4390 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8409  (
    .i0(\u2_Display/n4356 ),
    .i1(\u2_Display/n4383 [24]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4391 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u841  (
    .i0(\u2_Display/n436 ),
    .i1(\u2_Display/n454 [15]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n471 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8410  (
    .i0(\u2_Display/n4357 ),
    .i1(\u2_Display/n4383 [23]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4392 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8411  (
    .i0(\u2_Display/n4358 ),
    .i1(\u2_Display/n4383 [22]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4393 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8412  (
    .i0(\u2_Display/n4359 ),
    .i1(\u2_Display/n4383 [21]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4394 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8413  (
    .i0(\u2_Display/n4360 ),
    .i1(\u2_Display/n4383 [20]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4395 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8414  (
    .i0(\u2_Display/n4361 ),
    .i1(\u2_Display/n4383 [19]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4396 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8415  (
    .i0(\u2_Display/n4362 ),
    .i1(\u2_Display/n4383 [18]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4397 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8416  (
    .i0(\u2_Display/n4363 ),
    .i1(\u2_Display/n4383 [17]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4398 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8417  (
    .i0(\u2_Display/n4364 ),
    .i1(\u2_Display/n4383 [16]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4399 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8418  (
    .i0(\u2_Display/n4365 ),
    .i1(\u2_Display/n4383 [15]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4400 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8419  (
    .i0(\u2_Display/n4366 ),
    .i1(\u2_Display/n4383 [14]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4401 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u842  (
    .i0(\u2_Display/n437 ),
    .i1(\u2_Display/n454 [14]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n472 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8420  (
    .i0(\u2_Display/n4367 ),
    .i1(\u2_Display/n4383 [13]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4402 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8421  (
    .i0(\u2_Display/n4368 ),
    .i1(\u2_Display/n4383 [12]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4403 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8422  (
    .i0(\u2_Display/n4369 ),
    .i1(\u2_Display/n4383 [11]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4404 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8423  (
    .i0(\u2_Display/n4370 ),
    .i1(\u2_Display/n4383 [10]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4405 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8424  (
    .i0(\u2_Display/n4371 ),
    .i1(\u2_Display/n4383 [9]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4406 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8425  (
    .i0(\u2_Display/n4372 ),
    .i1(\u2_Display/n4383 [8]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4407 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8426  (
    .i0(\u2_Display/n4373 ),
    .i1(\u2_Display/n4383 [7]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4408 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8427  (
    .i0(\u2_Display/n4374 ),
    .i1(\u2_Display/n4383 [6]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4409 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8428  (
    .i0(\u2_Display/n4375 ),
    .i1(\u2_Display/n4383 [5]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4410 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8429  (
    .i0(\u2_Display/n4376 ),
    .i1(\u2_Display/n4383 [4]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4411 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u843  (
    .i0(\u2_Display/n438 ),
    .i1(\u2_Display/n454 [13]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n473 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8430  (
    .i0(\u2_Display/n4377 ),
    .i1(\u2_Display/n4383 [3]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4412 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8431  (
    .i0(\u2_Display/n4378 ),
    .i1(\u2_Display/n4383 [2]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4413 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8432  (
    .i0(\u2_Display/n4379 ),
    .i1(\u2_Display/n4383 [1]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4414 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8433  (
    .i0(\u2_Display/n4380 ),
    .i1(\u2_Display/n4383 [0]),
    .sel(\u2_Display/n4382 ),
    .o(\u2_Display/n4415 ));  // source/rtl/Display.v(195)
  not \u2_Display/u8434  (\u2_Display/n4417 , \u2_Display/n4416 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u844  (
    .i0(\u2_Display/n439 ),
    .i1(\u2_Display/n454 [12]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n474 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u845  (
    .i0(\u2_Display/n440 ),
    .i1(\u2_Display/n454 [11]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n475 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u846  (
    .i0(\u2_Display/n441 ),
    .i1(\u2_Display/n454 [10]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n476 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8467  (
    .i0(\u2_Display/n4384 ),
    .i1(\u2_Display/n4418 [31]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4419 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8468  (
    .i0(\u2_Display/n4385 ),
    .i1(\u2_Display/n4418 [30]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4420 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8469  (
    .i0(\u2_Display/n4386 ),
    .i1(\u2_Display/n4418 [29]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4421 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u847  (
    .i0(\u2_Display/n442 ),
    .i1(\u2_Display/n454 [9]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n477 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8470  (
    .i0(\u2_Display/n4387 ),
    .i1(\u2_Display/n4418 [28]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4422 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8471  (
    .i0(\u2_Display/n4388 ),
    .i1(\u2_Display/n4418 [27]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4423 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8472  (
    .i0(\u2_Display/n4389 ),
    .i1(\u2_Display/n4418 [26]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4424 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8473  (
    .i0(\u2_Display/n4390 ),
    .i1(\u2_Display/n4418 [25]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4425 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8474  (
    .i0(\u2_Display/n4391 ),
    .i1(\u2_Display/n4418 [24]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4426 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8475  (
    .i0(\u2_Display/n4392 ),
    .i1(\u2_Display/n4418 [23]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4427 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8476  (
    .i0(\u2_Display/n4393 ),
    .i1(\u2_Display/n4418 [22]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4428 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8477  (
    .i0(\u2_Display/n4394 ),
    .i1(\u2_Display/n4418 [21]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4429 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8478  (
    .i0(\u2_Display/n4395 ),
    .i1(\u2_Display/n4418 [20]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4430 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8479  (
    .i0(\u2_Display/n4396 ),
    .i1(\u2_Display/n4418 [19]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4431 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u848  (
    .i0(\u2_Display/n443 ),
    .i1(\u2_Display/n454 [8]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n478 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8480  (
    .i0(\u2_Display/n4397 ),
    .i1(\u2_Display/n4418 [18]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4432 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8481  (
    .i0(\u2_Display/n4398 ),
    .i1(\u2_Display/n4418 [17]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4433 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8482  (
    .i0(\u2_Display/n4399 ),
    .i1(\u2_Display/n4418 [16]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4434 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8483  (
    .i0(\u2_Display/n4400 ),
    .i1(\u2_Display/n4418 [15]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4435 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8484  (
    .i0(\u2_Display/n4401 ),
    .i1(\u2_Display/n4418 [14]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4436 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8485  (
    .i0(\u2_Display/n4402 ),
    .i1(\u2_Display/n4418 [13]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4437 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8486  (
    .i0(\u2_Display/n4403 ),
    .i1(\u2_Display/n4418 [12]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4438 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8487  (
    .i0(\u2_Display/n4404 ),
    .i1(\u2_Display/n4418 [11]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4439 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8488  (
    .i0(\u2_Display/n4405 ),
    .i1(\u2_Display/n4418 [10]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4440 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8489  (
    .i0(\u2_Display/n4406 ),
    .i1(\u2_Display/n4418 [9]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4441 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u849  (
    .i0(\u2_Display/n444 ),
    .i1(\u2_Display/n454 [7]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n479 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8490  (
    .i0(\u2_Display/n4407 ),
    .i1(\u2_Display/n4418 [8]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4442 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8491  (
    .i0(\u2_Display/n4408 ),
    .i1(\u2_Display/n4418 [7]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4443 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8492  (
    .i0(\u2_Display/n4409 ),
    .i1(\u2_Display/n4418 [6]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4444 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8493  (
    .i0(\u2_Display/n4410 ),
    .i1(\u2_Display/n4418 [5]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4445 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8494  (
    .i0(\u2_Display/n4411 ),
    .i1(\u2_Display/n4418 [4]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4446 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8495  (
    .i0(\u2_Display/n4412 ),
    .i1(\u2_Display/n4418 [3]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4447 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8496  (
    .i0(\u2_Display/n4413 ),
    .i1(\u2_Display/n4418 [2]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4448 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8497  (
    .i0(\u2_Display/n4414 ),
    .i1(\u2_Display/n4418 [1]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4449 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8498  (
    .i0(\u2_Display/n4415 ),
    .i1(\u2_Display/n4418 [0]),
    .sel(\u2_Display/n4417 ),
    .o(\u2_Display/n4450 ));  // source/rtl/Display.v(195)
  not \u2_Display/u8499  (\u2_Display/n4452 , \u2_Display/n4451 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u850  (
    .i0(\u2_Display/n445 ),
    .i1(\u2_Display/n454 [6]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n480 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u851  (
    .i0(\u2_Display/n446 ),
    .i1(\u2_Display/n454 [5]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n481 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u852  (
    .i0(\u2_Display/n447 ),
    .i1(\u2_Display/n454 [4]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n482 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u853  (
    .i0(\u2_Display/n448 ),
    .i1(\u2_Display/n454 [3]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n483 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8532  (
    .i0(\u2_Display/n4419 ),
    .i1(\u2_Display/n4453 [31]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4454 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8533  (
    .i0(\u2_Display/n4420 ),
    .i1(\u2_Display/n4453 [30]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4455 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8534  (
    .i0(\u2_Display/n4421 ),
    .i1(\u2_Display/n4453 [29]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4456 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8535  (
    .i0(\u2_Display/n4422 ),
    .i1(\u2_Display/n4453 [28]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4457 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8536  (
    .i0(\u2_Display/n4423 ),
    .i1(\u2_Display/n4453 [27]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4458 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8537  (
    .i0(\u2_Display/n4424 ),
    .i1(\u2_Display/n4453 [26]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4459 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8538  (
    .i0(\u2_Display/n4425 ),
    .i1(\u2_Display/n4453 [25]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4460 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8539  (
    .i0(\u2_Display/n4426 ),
    .i1(\u2_Display/n4453 [24]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4461 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u854  (
    .i0(\u2_Display/n449 ),
    .i1(\u2_Display/n454 [2]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n484 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8540  (
    .i0(\u2_Display/n4427 ),
    .i1(\u2_Display/n4453 [23]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4462 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8541  (
    .i0(\u2_Display/n4428 ),
    .i1(\u2_Display/n4453 [22]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4463 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8542  (
    .i0(\u2_Display/n4429 ),
    .i1(\u2_Display/n4453 [21]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4464 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8543  (
    .i0(\u2_Display/n4430 ),
    .i1(\u2_Display/n4453 [20]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4465 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8544  (
    .i0(\u2_Display/n4431 ),
    .i1(\u2_Display/n4453 [19]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4466 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8545  (
    .i0(\u2_Display/n4432 ),
    .i1(\u2_Display/n4453 [18]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4467 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8546  (
    .i0(\u2_Display/n4433 ),
    .i1(\u2_Display/n4453 [17]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4468 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8547  (
    .i0(\u2_Display/n4434 ),
    .i1(\u2_Display/n4453 [16]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4469 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8548  (
    .i0(\u2_Display/n4435 ),
    .i1(\u2_Display/n4453 [15]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4470 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8549  (
    .i0(\u2_Display/n4436 ),
    .i1(\u2_Display/n4453 [14]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4471 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u855  (
    .i0(\u2_Display/n450 ),
    .i1(\u2_Display/n454 [1]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n485 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8550  (
    .i0(\u2_Display/n4437 ),
    .i1(\u2_Display/n4453 [13]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4472 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8551  (
    .i0(\u2_Display/n4438 ),
    .i1(\u2_Display/n4453 [12]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4473 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8552  (
    .i0(\u2_Display/n4439 ),
    .i1(\u2_Display/n4453 [11]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4474 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8553  (
    .i0(\u2_Display/n4440 ),
    .i1(\u2_Display/n4453 [10]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4475 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8554  (
    .i0(\u2_Display/n4441 ),
    .i1(\u2_Display/n4453 [9]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4476 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8555  (
    .i0(\u2_Display/n4442 ),
    .i1(\u2_Display/n4453 [8]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4477 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8556  (
    .i0(\u2_Display/n4443 ),
    .i1(\u2_Display/n4453 [7]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4478 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8557  (
    .i0(\u2_Display/n4444 ),
    .i1(\u2_Display/n4453 [6]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4479 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8558  (
    .i0(\u2_Display/n4445 ),
    .i1(\u2_Display/n4453 [5]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4480 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8559  (
    .i0(\u2_Display/n4446 ),
    .i1(\u2_Display/n4453 [4]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4481 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u856  (
    .i0(\u2_Display/n451 ),
    .i1(\u2_Display/n454 [0]),
    .sel(\u2_Display/n453 ),
    .o(\u2_Display/n486 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8560  (
    .i0(\u2_Display/n4447 ),
    .i1(\u2_Display/n4453 [3]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4482 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8561  (
    .i0(\u2_Display/n4448 ),
    .i1(\u2_Display/n4453 [2]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4483 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8562  (
    .i0(\u2_Display/n4449 ),
    .i1(\u2_Display/n4453 [1]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4484 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8563  (
    .i0(\u2_Display/n4450 ),
    .i1(\u2_Display/n4453 [0]),
    .sel(\u2_Display/n4452 ),
    .o(\u2_Display/n4485 ));  // source/rtl/Display.v(195)
  not \u2_Display/u8564  (\u2_Display/n4487 , \u2_Display/n4486 );  // source/rtl/Display.v(195)
  not \u2_Display/u857  (\u2_Display/n488 , \u2_Display/n487 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u8597  (
    .i0(\u2_Display/n4454 ),
    .i1(\u2_Display/n4488 [31]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4489 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8598  (
    .i0(\u2_Display/n4455 ),
    .i1(\u2_Display/n4488 [30]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4490 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8599  (
    .i0(\u2_Display/n4456 ),
    .i1(\u2_Display/n4488 [29]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4491 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8600  (
    .i0(\u2_Display/n4457 ),
    .i1(\u2_Display/n4488 [28]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4492 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8601  (
    .i0(\u2_Display/n4458 ),
    .i1(\u2_Display/n4488 [27]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4493 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8602  (
    .i0(\u2_Display/n4459 ),
    .i1(\u2_Display/n4488 [26]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4494 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8603  (
    .i0(\u2_Display/n4460 ),
    .i1(\u2_Display/n4488 [25]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4495 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8604  (
    .i0(\u2_Display/n4461 ),
    .i1(\u2_Display/n4488 [24]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4496 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8605  (
    .i0(\u2_Display/n4462 ),
    .i1(\u2_Display/n4488 [23]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4497 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8606  (
    .i0(\u2_Display/n4463 ),
    .i1(\u2_Display/n4488 [22]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4498 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8607  (
    .i0(\u2_Display/n4464 ),
    .i1(\u2_Display/n4488 [21]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4499 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8608  (
    .i0(\u2_Display/n4465 ),
    .i1(\u2_Display/n4488 [20]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4500 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8609  (
    .i0(\u2_Display/n4466 ),
    .i1(\u2_Display/n4488 [19]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4501 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8610  (
    .i0(\u2_Display/n4467 ),
    .i1(\u2_Display/n4488 [18]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4502 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8611  (
    .i0(\u2_Display/n4468 ),
    .i1(\u2_Display/n4488 [17]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4503 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8612  (
    .i0(\u2_Display/n4469 ),
    .i1(\u2_Display/n4488 [16]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4504 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8613  (
    .i0(\u2_Display/n4470 ),
    .i1(\u2_Display/n4488 [15]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4505 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8614  (
    .i0(\u2_Display/n4471 ),
    .i1(\u2_Display/n4488 [14]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4506 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8615  (
    .i0(\u2_Display/n4472 ),
    .i1(\u2_Display/n4488 [13]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4507 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8616  (
    .i0(\u2_Display/n4473 ),
    .i1(\u2_Display/n4488 [12]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4508 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8617  (
    .i0(\u2_Display/n4474 ),
    .i1(\u2_Display/n4488 [11]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4509 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8618  (
    .i0(\u2_Display/n4475 ),
    .i1(\u2_Display/n4488 [10]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4510 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8619  (
    .i0(\u2_Display/n4476 ),
    .i1(\u2_Display/n4488 [9]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4511 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8620  (
    .i0(\u2_Display/n4477 ),
    .i1(\u2_Display/n4488 [8]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4512 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8621  (
    .i0(\u2_Display/n4478 ),
    .i1(\u2_Display/n4488 [7]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4513 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8622  (
    .i0(\u2_Display/n4479 ),
    .i1(\u2_Display/n4488 [6]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4514 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8623  (
    .i0(\u2_Display/n4480 ),
    .i1(\u2_Display/n4488 [5]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4515 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8624  (
    .i0(\u2_Display/n4481 ),
    .i1(\u2_Display/n4488 [4]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4516 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8625  (
    .i0(\u2_Display/n4482 ),
    .i1(\u2_Display/n4488 [3]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4517 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8626  (
    .i0(\u2_Display/n4483 ),
    .i1(\u2_Display/n4488 [2]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4518 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8627  (
    .i0(\u2_Display/n4484 ),
    .i1(\u2_Display/n4488 [1]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4519 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8628  (
    .i0(\u2_Display/n4485 ),
    .i1(\u2_Display/n4488 [0]),
    .sel(\u2_Display/n4487 ),
    .o(\u2_Display/n4520 ));  // source/rtl/Display.v(195)
  not \u2_Display/u8629  (\u2_Display/n4522 , \u2_Display/n4521 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8662  (
    .i0(\u2_Display/n4489 ),
    .i1(\u2_Display/n4523 [31]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4524 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8663  (
    .i0(\u2_Display/n4490 ),
    .i1(\u2_Display/n4523 [30]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4525 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8664  (
    .i0(\u2_Display/n4491 ),
    .i1(\u2_Display/n4523 [29]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4526 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8665  (
    .i0(\u2_Display/n4492 ),
    .i1(\u2_Display/n4523 [28]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4527 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8666  (
    .i0(\u2_Display/n4493 ),
    .i1(\u2_Display/n4523 [27]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4528 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8667  (
    .i0(\u2_Display/n4494 ),
    .i1(\u2_Display/n4523 [26]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4529 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8668  (
    .i0(\u2_Display/n4495 ),
    .i1(\u2_Display/n4523 [25]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4530 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8669  (
    .i0(\u2_Display/n4496 ),
    .i1(\u2_Display/n4523 [24]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4531 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8670  (
    .i0(\u2_Display/n4497 ),
    .i1(\u2_Display/n4523 [23]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4532 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8671  (
    .i0(\u2_Display/n4498 ),
    .i1(\u2_Display/n4523 [22]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4533 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8672  (
    .i0(\u2_Display/n4499 ),
    .i1(\u2_Display/n4523 [21]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4534 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8673  (
    .i0(\u2_Display/n4500 ),
    .i1(\u2_Display/n4523 [20]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4535 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8674  (
    .i0(\u2_Display/n4501 ),
    .i1(\u2_Display/n4523 [19]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4536 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8675  (
    .i0(\u2_Display/n4502 ),
    .i1(\u2_Display/n4523 [18]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4537 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8676  (
    .i0(\u2_Display/n4503 ),
    .i1(\u2_Display/n4523 [17]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4538 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8677  (
    .i0(\u2_Display/n4504 ),
    .i1(\u2_Display/n4523 [16]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4539 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8678  (
    .i0(\u2_Display/n4505 ),
    .i1(\u2_Display/n4523 [15]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4540 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8679  (
    .i0(\u2_Display/n4506 ),
    .i1(\u2_Display/n4523 [14]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4541 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8680  (
    .i0(\u2_Display/n4507 ),
    .i1(\u2_Display/n4523 [13]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4542 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8681  (
    .i0(\u2_Display/n4508 ),
    .i1(\u2_Display/n4523 [12]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4543 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8682  (
    .i0(\u2_Display/n4509 ),
    .i1(\u2_Display/n4523 [11]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4544 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8683  (
    .i0(\u2_Display/n4510 ),
    .i1(\u2_Display/n4523 [10]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4545 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8684  (
    .i0(\u2_Display/n4511 ),
    .i1(\u2_Display/n4523 [9]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4546 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8685  (
    .i0(\u2_Display/n4512 ),
    .i1(\u2_Display/n4523 [8]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4547 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8686  (
    .i0(\u2_Display/n4513 ),
    .i1(\u2_Display/n4523 [7]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4548 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8687  (
    .i0(\u2_Display/n4514 ),
    .i1(\u2_Display/n4523 [6]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4549 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8688  (
    .i0(\u2_Display/n4515 ),
    .i1(\u2_Display/n4523 [5]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4550 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8689  (
    .i0(\u2_Display/n4516 ),
    .i1(\u2_Display/n4523 [4]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4551 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8690  (
    .i0(\u2_Display/n4517 ),
    .i1(\u2_Display/n4523 [3]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4552 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8691  (
    .i0(\u2_Display/n4518 ),
    .i1(\u2_Display/n4523 [2]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4553 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8692  (
    .i0(\u2_Display/n4519 ),
    .i1(\u2_Display/n4523 [1]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4554 ));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8693  (
    .i0(\u2_Display/n4520 ),
    .i1(\u2_Display/n4523 [0]),
    .sel(\u2_Display/n4522 ),
    .o(\u2_Display/n4555 ));  // source/rtl/Display.v(195)
  not \u2_Display/u8694  (\u2_Display/n4557 , \u2_Display/n4556 );  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8727  (
    .i0(\u2_Display/n4546 ),
    .i1(\u2_Display/n4558 [9]),
    .sel(\u2_Display/n4557 ),
    .o(\u2_Display/n133 [9]));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8728  (
    .i0(\u2_Display/n4547 ),
    .i1(\u2_Display/n4558 [8]),
    .sel(\u2_Display/n4557 ),
    .o(\u2_Display/n133 [8]));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8729  (
    .i0(\u2_Display/n4548 ),
    .i1(\u2_Display/n4558 [7]),
    .sel(\u2_Display/n4557 ),
    .o(\u2_Display/n133 [7]));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8730  (
    .i0(\u2_Display/n4549 ),
    .i1(\u2_Display/n4558 [6]),
    .sel(\u2_Display/n4557 ),
    .o(\u2_Display/n133 [6]));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8731  (
    .i0(\u2_Display/n4550 ),
    .i1(\u2_Display/n4558 [5]),
    .sel(\u2_Display/n4557 ),
    .o(\u2_Display/n133 [5]));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8732  (
    .i0(\u2_Display/n4551 ),
    .i1(\u2_Display/n4558 [4]),
    .sel(\u2_Display/n4557 ),
    .o(\u2_Display/n133 [4]));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8733  (
    .i0(\u2_Display/n4552 ),
    .i1(\u2_Display/n4558 [3]),
    .sel(\u2_Display/n4557 ),
    .o(\u2_Display/n133 [3]));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8734  (
    .i0(\u2_Display/n4553 ),
    .i1(\u2_Display/n4558 [2]),
    .sel(\u2_Display/n4557 ),
    .o(\u2_Display/n133 [2]));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8735  (
    .i0(\u2_Display/n4554 ),
    .i1(\u2_Display/n4558 [1]),
    .sel(\u2_Display/n4557 ),
    .o(\u2_Display/n133 [1]));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u8736  (
    .i0(\u2_Display/n4555 ),
    .i1(\u2_Display/n4558 [0]),
    .sel(\u2_Display/n4557 ),
    .o(\u2_Display/n133 [0]));  // source/rtl/Display.v(195)
  AL_MUX \u2_Display/u890  (
    .i0(\u2_Display/n455 ),
    .i1(\u2_Display/n489 [31]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n490 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u891  (
    .i0(\u2_Display/n456 ),
    .i1(\u2_Display/n489 [30]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n491 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u892  (
    .i0(\u2_Display/n457 ),
    .i1(\u2_Display/n489 [29]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n492 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u893  (
    .i0(\u2_Display/n458 ),
    .i1(\u2_Display/n489 [28]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n493 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u894  (
    .i0(\u2_Display/n459 ),
    .i1(\u2_Display/n489 [27]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n494 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u895  (
    .i0(\u2_Display/n460 ),
    .i1(\u2_Display/n489 [26]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n495 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u896  (
    .i0(\u2_Display/n461 ),
    .i1(\u2_Display/n489 [25]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n496 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u897  (
    .i0(\u2_Display/n462 ),
    .i1(\u2_Display/n489 [24]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n497 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u898  (
    .i0(\u2_Display/n463 ),
    .i1(\u2_Display/n489 [23]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n498 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u899  (
    .i0(\u2_Display/n464 ),
    .i1(\u2_Display/n489 [22]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n499 ));  // source/rtl/Display.v(230)
  and \u2_Display/u9  (\u2_Display/n46 , \u2_Display/n44 , \u2_Display/n45 );  // source/rtl/Display.v(165)
  AL_MUX \u2_Display/u900  (
    .i0(\u2_Display/n465 ),
    .i1(\u2_Display/n489 [21]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n500 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u901  (
    .i0(\u2_Display/n466 ),
    .i1(\u2_Display/n489 [20]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n501 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u902  (
    .i0(\u2_Display/n467 ),
    .i1(\u2_Display/n489 [19]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n502 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u903  (
    .i0(\u2_Display/n468 ),
    .i1(\u2_Display/n489 [18]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n503 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u904  (
    .i0(\u2_Display/n469 ),
    .i1(\u2_Display/n489 [17]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n504 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u905  (
    .i0(\u2_Display/n470 ),
    .i1(\u2_Display/n489 [16]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n505 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u906  (
    .i0(\u2_Display/n471 ),
    .i1(\u2_Display/n489 [15]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n506 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u907  (
    .i0(\u2_Display/n472 ),
    .i1(\u2_Display/n489 [14]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n507 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u908  (
    .i0(\u2_Display/n473 ),
    .i1(\u2_Display/n489 [13]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n508 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u909  (
    .i0(\u2_Display/n474 ),
    .i1(\u2_Display/n489 [12]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n509 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u910  (
    .i0(\u2_Display/n475 ),
    .i1(\u2_Display/n489 [11]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n510 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u911  (
    .i0(\u2_Display/n476 ),
    .i1(\u2_Display/n489 [10]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n511 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u912  (
    .i0(\u2_Display/n477 ),
    .i1(\u2_Display/n489 [9]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n512 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u913  (
    .i0(\u2_Display/n478 ),
    .i1(\u2_Display/n489 [8]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n513 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u914  (
    .i0(\u2_Display/n479 ),
    .i1(\u2_Display/n489 [7]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n514 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u915  (
    .i0(\u2_Display/n480 ),
    .i1(\u2_Display/n489 [6]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n515 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u916  (
    .i0(\u2_Display/n481 ),
    .i1(\u2_Display/n489 [5]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n516 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u917  (
    .i0(\u2_Display/n482 ),
    .i1(\u2_Display/n489 [4]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n517 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u918  (
    .i0(\u2_Display/n483 ),
    .i1(\u2_Display/n489 [3]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n518 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u919  (
    .i0(\u2_Display/n484 ),
    .i1(\u2_Display/n489 [2]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n519 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u920  (
    .i0(\u2_Display/n485 ),
    .i1(\u2_Display/n489 [1]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n520 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u921  (
    .i0(\u2_Display/n486 ),
    .i1(\u2_Display/n489 [0]),
    .sel(\u2_Display/n488 ),
    .o(\u2_Display/n521 ));  // source/rtl/Display.v(230)
  not \u2_Display/u922  (\u2_Display/n523 , \u2_Display/n522 );  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u955  (
    .i0(\u2_Display/n490 ),
    .i1(\u2_Display/n524 [31]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n525 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u956  (
    .i0(\u2_Display/n491 ),
    .i1(\u2_Display/n524 [30]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n526 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u957  (
    .i0(\u2_Display/n492 ),
    .i1(\u2_Display/n524 [29]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n527 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u958  (
    .i0(\u2_Display/n493 ),
    .i1(\u2_Display/n524 [28]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n528 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u959  (
    .i0(\u2_Display/n494 ),
    .i1(\u2_Display/n524 [27]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n529 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u960  (
    .i0(\u2_Display/n495 ),
    .i1(\u2_Display/n524 [26]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n530 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u961  (
    .i0(\u2_Display/n496 ),
    .i1(\u2_Display/n524 [25]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n531 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u962  (
    .i0(\u2_Display/n497 ),
    .i1(\u2_Display/n524 [24]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n532 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u963  (
    .i0(\u2_Display/n498 ),
    .i1(\u2_Display/n524 [23]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n533 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u964  (
    .i0(\u2_Display/n499 ),
    .i1(\u2_Display/n524 [22]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n534 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u965  (
    .i0(\u2_Display/n500 ),
    .i1(\u2_Display/n524 [21]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n535 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u966  (
    .i0(\u2_Display/n501 ),
    .i1(\u2_Display/n524 [20]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n536 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u967  (
    .i0(\u2_Display/n502 ),
    .i1(\u2_Display/n524 [19]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n537 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u968  (
    .i0(\u2_Display/n503 ),
    .i1(\u2_Display/n524 [18]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n538 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u969  (
    .i0(\u2_Display/n504 ),
    .i1(\u2_Display/n524 [17]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n539 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u970  (
    .i0(\u2_Display/n505 ),
    .i1(\u2_Display/n524 [16]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n540 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u971  (
    .i0(\u2_Display/n506 ),
    .i1(\u2_Display/n524 [15]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n541 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u972  (
    .i0(\u2_Display/n507 ),
    .i1(\u2_Display/n524 [14]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n542 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u973  (
    .i0(\u2_Display/n508 ),
    .i1(\u2_Display/n524 [13]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n543 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u974  (
    .i0(\u2_Display/n509 ),
    .i1(\u2_Display/n524 [12]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n544 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u975  (
    .i0(\u2_Display/n510 ),
    .i1(\u2_Display/n524 [11]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n545 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u976  (
    .i0(\u2_Display/n511 ),
    .i1(\u2_Display/n524 [10]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n546 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u977  (
    .i0(\u2_Display/n512 ),
    .i1(\u2_Display/n524 [9]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n547 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u978  (
    .i0(\u2_Display/n513 ),
    .i1(\u2_Display/n524 [8]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n548 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u979  (
    .i0(\u2_Display/n514 ),
    .i1(\u2_Display/n524 [7]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n549 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u980  (
    .i0(\u2_Display/n515 ),
    .i1(\u2_Display/n524 [6]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n550 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u981  (
    .i0(\u2_Display/n516 ),
    .i1(\u2_Display/n524 [5]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n551 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u982  (
    .i0(\u2_Display/n517 ),
    .i1(\u2_Display/n524 [4]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n552 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u983  (
    .i0(\u2_Display/n518 ),
    .i1(\u2_Display/n524 [3]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n553 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u984  (
    .i0(\u2_Display/n519 ),
    .i1(\u2_Display/n524 [2]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n554 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u985  (
    .i0(\u2_Display/n520 ),
    .i1(\u2_Display/n524 [1]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n555 ));  // source/rtl/Display.v(230)
  AL_MUX \u2_Display/u986  (
    .i0(\u2_Display/n521 ),
    .i1(\u2_Display/n524 [0]),
    .sel(\u2_Display/n523 ),
    .o(\u2_Display/n556 ));  // source/rtl/Display.v(230)
  not \u2_Display/u987  (\u2_Display/n558 , \u2_Display/n557 );  // source/rtl/Display.v(230)

endmodule 

module add_pu12_pu12_o12
  (
  i0,
  i1,
  o
  );

  input [11:0] i0;
  input [11:0] i1;
  output [11:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module eq_w12
  (
  i0,
  i1,
  o
  );

  input [11:0] i0;
  input [11:0] i1;
  output o;

  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[6]_i1[6_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[10]_i1[10]_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[7]_i1[7]_o_o ;
  wire \or_xor_i0[9]_i1[9]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, \or_or_or_xor_i0[0]_i_o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[6]_i1[6_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[3]_i1[3]_o_o );
  or \or_or_xor_i0[6]_i1[6  (\or_or_xor_i0[6]_i1[6_o , \or_xor_i0[6]_i1[6]_o_o , \or_xor_i0[9]_i1[9]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[10]_i1[10]  (\or_xor_i0[10]_i1[10]_o , \xor_i0[10]_i1[10]_o , \xor_i0[11]_i1[11]_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \or_xor_i0[4]_i1[4]_o_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \or_xor_i0[7]_i1[7]_o_o );
  or \or_xor_i0[7]_i1[7]_o  (\or_xor_i0[7]_i1[7]_o_o , \xor_i0[7]_i1[7]_o , \xor_i0[8]_i1[8]_o );
  or \or_xor_i0[9]_i1[9]_o  (\or_xor_i0[9]_i1[9]_o_o , \xor_i0[9]_i1[9]_o , \or_xor_i0[10]_i1[10]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module lt_u12_u12
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [11:0] i0;
  input [11:0] i1;
  output o;

  wire [11:0] diff;
  wire diff_6_11;
  wire less_6_11;
  wire \less_6_11_inst/diff_0 ;
  wire \less_6_11_inst/diff_1 ;
  wire \less_6_11_inst/diff_2 ;
  wire \less_6_11_inst/diff_3 ;
  wire \less_6_11_inst/diff_4 ;
  wire \less_6_11_inst/diff_5 ;
  wire \less_6_11_inst/o_0 ;
  wire \less_6_11_inst/o_1 ;
  wire \less_6_11_inst/o_2 ;
  wire \less_6_11_inst/o_3 ;
  wire \less_6_11_inst/o_4 ;
  wire o_0;
  wire o_1;
  wire o_2;
  wire o_3;
  wire o_4;
  wire o_5;

  or any_diff_6_11 (diff_6_11, diff[6], diff[7], diff[8], diff[9], diff[10], diff[11]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);
  AL_MUX \less_6_11_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[6]),
    .sel(\less_6_11_inst/diff_0 ),
    .o(\less_6_11_inst/o_0 ));
  AL_MUX \less_6_11_inst/mux_1  (
    .i0(\less_6_11_inst/o_0 ),
    .i1(i1[7]),
    .sel(\less_6_11_inst/diff_1 ),
    .o(\less_6_11_inst/o_1 ));
  AL_MUX \less_6_11_inst/mux_2  (
    .i0(\less_6_11_inst/o_1 ),
    .i1(i1[8]),
    .sel(\less_6_11_inst/diff_2 ),
    .o(\less_6_11_inst/o_2 ));
  AL_MUX \less_6_11_inst/mux_3  (
    .i0(\less_6_11_inst/o_2 ),
    .i1(i1[9]),
    .sel(\less_6_11_inst/diff_3 ),
    .o(\less_6_11_inst/o_3 ));
  AL_MUX \less_6_11_inst/mux_4  (
    .i0(\less_6_11_inst/o_3 ),
    .i1(i1[10]),
    .sel(\less_6_11_inst/diff_4 ),
    .o(\less_6_11_inst/o_4 ));
  AL_MUX \less_6_11_inst/mux_5  (
    .i0(\less_6_11_inst/o_4 ),
    .i1(i1[11]),
    .sel(\less_6_11_inst/diff_5 ),
    .o(less_6_11));
  xor \less_6_11_inst/xor_0  (\less_6_11_inst/diff_0 , i0[6], i1[6]);
  xor \less_6_11_inst/xor_1  (\less_6_11_inst/diff_1 , i0[7], i1[7]);
  xor \less_6_11_inst/xor_2  (\less_6_11_inst/diff_2 , i0[8], i1[8]);
  xor \less_6_11_inst/xor_3  (\less_6_11_inst/diff_3 , i0[9], i1[9]);
  xor \less_6_11_inst/xor_4  (\less_6_11_inst/diff_4 , i0[10], i1[10]);
  xor \less_6_11_inst/xor_5  (\less_6_11_inst/diff_5 , i0[11], i1[11]);
  AL_MUX mux_0 (
    .i0(ci),
    .i1(i1[0]),
    .sel(diff[0]),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(i1[1]),
    .sel(diff[1]),
    .o(o_1));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(i1[2]),
    .sel(diff[2]),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(i1[3]),
    .sel(diff[3]),
    .o(o_3));
  AL_MUX mux_4 (
    .i0(o_3),
    .i1(i1[4]),
    .sel(diff[4]),
    .o(o_4));
  AL_MUX mux_5 (
    .i0(o_4),
    .i1(i1[5]),
    .sel(diff[5]),
    .o(o_5));
  AL_MUX mux_6 (
    .i0(o_5),
    .i1(less_6_11),
    .sel(diff_6_11),
    .o(o));

endmodule 

module binary_mux_s1_w1
  (
  i0,
  i1,
  sel,
  o
  );

  input i0;
  input i1;
  input sel;
  output o;


  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel),
    .o(o));

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module add_pu12_mu12_o12
  (
  i0,
  i1,
  o
  );

  input [11:0] i0;
  input [11:0] i1;
  output [11:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_nb0;
  wire net_nb1;
  wire net_nb10;
  wire net_nb11;
  wire net_nb2;
  wire net_nb3;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_nb9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_nb10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_nb11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_nb9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b10 (net_nb10, net_b10);
  not inv_b11 (net_nb11, net_b11);
  not inv_b2 (net_nb2, net_b2);
  not inv_b3 (net_nb3, net_b3);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);
  not inv_b9 (net_nb9, net_b9);

endmodule 

module add_pu31_pu31_o31
  (
  i0,
  i1,
  o
  );

  input [30:0] i0;
  input [30:0] i1;
  output [30:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module add_pu32_pu32_o32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output [31:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_b31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module add_pu32_pu32_pu1_o32
  (
  i0,
  i1,
  i2,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  input i2;
  output [31:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cin;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign net_cin = i2;
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(net_cin),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_b31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module add_pu10_pu10_pu1_o10
  (
  i0,
  i1,
  i2,
  o
  );

  input [9:0] i0;
  input [9:0] i1;
  input i2;
  output [9:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cin;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign net_cin = i2;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(net_cin),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module add_pu11_pu11_pu1_o11
  (
  i0,
  i1,
  i2,
  o
  );

  input [10:0] i0;
  input [10:0] i1;
  input i2;
  output [10:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cin;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign net_cin = i2;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(net_cin),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module add_pu3_pu3_o4
  (
  i0,
  i1,
  o
  );

  input [2:0] i0;
  input [2:0] i1;
  output [3:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;

  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[3] = net_cout2;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));

endmodule 

module add_pu4_pu4_o5
  (
  i0,
  i1,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  output [4:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;

  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[4] = net_cout3;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));

endmodule 

module add_pu1_pu1_o2
  (
  i0,
  i1,
  o
  );

  input i0;
  input i1;
  output [1:0] o;

  wire net_a0;
  wire net_cin;
  wire net_cout0;
  wire net_sum0;

  assign net_a0 = i0;
  assign net_cin = i1;
  assign o[1] = net_cout0;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(1'b0),
    .c(net_cin),
    .cout(net_cout0),
    .sum(net_sum0));

endmodule 

module add_pu2_pu2_o3
  (
  i0,
  i1,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  output [2:0] o;

  wire net_a0;
  wire net_a1;
  wire net_b0;
  wire net_b1;
  wire net_cout0;
  wire net_cout1;
  wire net_sum0;
  wire net_sum1;

  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[2] = net_cout1;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));

endmodule 

module eq_w31
  (
  i0,
  i1,
  o
  );

  input [30:0] i0;
  input [30:0] i1;
  output o;

  wire \or_or_or_or_xor_i0[0_o ;
  wire \or_or_or_or_xor_i0[1_o ;
  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_or_xor_i0[15]__o ;
  wire \or_or_or_xor_i0[23]__o ;
  wire \or_or_or_xor_i0[7]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[11]_i1[_o ;
  wire \or_or_xor_i0[15]_i1[_o ;
  wire \or_or_xor_i0[19]_i1[_o ;
  wire \or_or_xor_i0[23]_i1[_o ;
  wire \or_or_xor_i0[27]_i1[_o ;
  wire \or_or_xor_i0[3]_i1[3_o ;
  wire \or_or_xor_i0[7]_i1[7_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[11]_i1[11]_o ;
  wire \or_xor_i0[13]_i1[13]_o ;
  wire \or_xor_i0[15]_i1[15]_o ;
  wire \or_xor_i0[17]_i1[17]_o ;
  wire \or_xor_i0[19]_i1[19]_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \or_xor_i0[21]_i1[21]_o ;
  wire \or_xor_i0[23]_i1[23]_o ;
  wire \or_xor_i0[25]_i1[25]_o ;
  wire \or_xor_i0[27]_i1[27]_o ;
  wire \or_xor_i0[29]_i1[29]_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[5]_i1[5]_o_o ;
  wire \or_xor_i0[7]_i1[7]_o_o ;
  wire \or_xor_i0[9]_i1[9]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[12]_i1[12]_o ;
  wire \xor_i0[13]_i1[13]_o ;
  wire \xor_i0[14]_i1[14]_o ;
  wire \xor_i0[15]_i1[15]_o ;
  wire \xor_i0[16]_i1[16]_o ;
  wire \xor_i0[17]_i1[17]_o ;
  wire \xor_i0[18]_i1[18]_o ;
  wire \xor_i0[19]_i1[19]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[20]_i1[20]_o ;
  wire \xor_i0[21]_i1[21]_o ;
  wire \xor_i0[22]_i1[22]_o ;
  wire \xor_i0[23]_i1[23]_o ;
  wire \xor_i0[24]_i1[24]_o ;
  wire \xor_i0[25]_i1[25]_o ;
  wire \xor_i0[26]_i1[26]_o ;
  wire \xor_i0[27]_i1[27]_o ;
  wire \xor_i0[28]_i1[28]_o ;
  wire \xor_i0[29]_i1[29]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[30]_i1[30]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, \or_or_or_or_xor_i0[0_o );
  or \or_or_or_or_xor_i0[0  (\or_or_or_or_xor_i0[0_o , \or_or_or_xor_i0[0]_i_o , \or_or_or_or_xor_i0[1_o );
  or \or_or_or_or_xor_i0[1  (\or_or_or_or_xor_i0[1_o , \or_or_or_xor_i0[15]__o , \or_or_or_xor_i0[23]__o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_or_xor_i0[7]_i_o );
  or \or_or_or_xor_i0[15]_  (\or_or_or_xor_i0[15]__o , \or_or_xor_i0[15]_i1[_o , \or_or_xor_i0[19]_i1[_o );
  or \or_or_or_xor_i0[23]_  (\or_or_or_xor_i0[23]__o , \or_or_xor_i0[23]_i1[_o , \or_or_xor_i0[27]_i1[_o );
  or \or_or_or_xor_i0[7]_i  (\or_or_or_xor_i0[7]_i_o , \or_or_xor_i0[7]_i1[7_o , \or_or_xor_i0[11]_i1[_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_or_xor_i0[3]_i1[3_o );
  or \or_or_xor_i0[11]_i1[  (\or_or_xor_i0[11]_i1[_o , \or_xor_i0[11]_i1[11]_o , \or_xor_i0[13]_i1[13]_o );
  or \or_or_xor_i0[15]_i1[  (\or_or_xor_i0[15]_i1[_o , \or_xor_i0[15]_i1[15]_o , \or_xor_i0[17]_i1[17]_o );
  or \or_or_xor_i0[19]_i1[  (\or_or_xor_i0[19]_i1[_o , \or_xor_i0[19]_i1[19]_o , \or_xor_i0[21]_i1[21]_o );
  or \or_or_xor_i0[23]_i1[  (\or_or_xor_i0[23]_i1[_o , \or_xor_i0[23]_i1[23]_o , \or_xor_i0[25]_i1[25]_o );
  or \or_or_xor_i0[27]_i1[  (\or_or_xor_i0[27]_i1[_o , \or_xor_i0[27]_i1[27]_o , \or_xor_i0[29]_i1[29]_o );
  or \or_or_xor_i0[3]_i1[3  (\or_or_xor_i0[3]_i1[3_o , \or_xor_i0[3]_i1[3]_o_o , \or_xor_i0[5]_i1[5]_o_o );
  or \or_or_xor_i0[7]_i1[7  (\or_or_xor_i0[7]_i1[7_o , \or_xor_i0[7]_i1[7]_o_o , \or_xor_i0[9]_i1[9]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[11]_i1[11]  (\or_xor_i0[11]_i1[11]_o , \xor_i0[11]_i1[11]_o , \xor_i0[12]_i1[12]_o );
  or \or_xor_i0[13]_i1[13]  (\or_xor_i0[13]_i1[13]_o , \xor_i0[13]_i1[13]_o , \xor_i0[14]_i1[14]_o );
  or \or_xor_i0[15]_i1[15]  (\or_xor_i0[15]_i1[15]_o , \xor_i0[15]_i1[15]_o , \xor_i0[16]_i1[16]_o );
  or \or_xor_i0[17]_i1[17]  (\or_xor_i0[17]_i1[17]_o , \xor_i0[17]_i1[17]_o , \xor_i0[18]_i1[18]_o );
  or \or_xor_i0[19]_i1[19]  (\or_xor_i0[19]_i1[19]_o , \xor_i0[19]_i1[19]_o , \xor_i0[20]_i1[20]_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  or \or_xor_i0[21]_i1[21]  (\or_xor_i0[21]_i1[21]_o , \xor_i0[21]_i1[21]_o , \xor_i0[22]_i1[22]_o );
  or \or_xor_i0[23]_i1[23]  (\or_xor_i0[23]_i1[23]_o , \xor_i0[23]_i1[23]_o , \xor_i0[24]_i1[24]_o );
  or \or_xor_i0[25]_i1[25]  (\or_xor_i0[25]_i1[25]_o , \xor_i0[25]_i1[25]_o , \xor_i0[26]_i1[26]_o );
  or \or_xor_i0[27]_i1[27]  (\or_xor_i0[27]_i1[27]_o , \xor_i0[27]_i1[27]_o , \xor_i0[28]_i1[28]_o );
  or \or_xor_i0[29]_i1[29]  (\or_xor_i0[29]_i1[29]_o , \xor_i0[29]_i1[29]_o , \xor_i0[30]_i1[30]_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \xor_i0[4]_i1[4]_o );
  or \or_xor_i0[5]_i1[5]_o  (\or_xor_i0[5]_i1[5]_o_o , \xor_i0[5]_i1[5]_o , \xor_i0[6]_i1[6]_o );
  or \or_xor_i0[7]_i1[7]_o  (\or_xor_i0[7]_i1[7]_o_o , \xor_i0[7]_i1[7]_o , \xor_i0[8]_i1[8]_o );
  or \or_xor_i0[9]_i1[9]_o  (\or_xor_i0[9]_i1[9]_o_o , \xor_i0[9]_i1[9]_o , \xor_i0[10]_i1[10]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (\xor_i0[12]_i1[12]_o , i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (\xor_i0[13]_i1[13]_o , i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (\xor_i0[14]_i1[14]_o , i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (\xor_i0[15]_i1[15]_o , i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (\xor_i0[16]_i1[16]_o , i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (\xor_i0[17]_i1[17]_o , i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (\xor_i0[18]_i1[18]_o , i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (\xor_i0[19]_i1[19]_o , i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[20]_i1[20]  (\xor_i0[20]_i1[20]_o , i0[20], i1[20]);
  xor \xor_i0[21]_i1[21]  (\xor_i0[21]_i1[21]_o , i0[21], i1[21]);
  xor \xor_i0[22]_i1[22]  (\xor_i0[22]_i1[22]_o , i0[22], i1[22]);
  xor \xor_i0[23]_i1[23]  (\xor_i0[23]_i1[23]_o , i0[23], i1[23]);
  xor \xor_i0[24]_i1[24]  (\xor_i0[24]_i1[24]_o , i0[24], i1[24]);
  xor \xor_i0[25]_i1[25]  (\xor_i0[25]_i1[25]_o , i0[25], i1[25]);
  xor \xor_i0[26]_i1[26]  (\xor_i0[26]_i1[26]_o , i0[26], i1[26]);
  xor \xor_i0[27]_i1[27]  (\xor_i0[27]_i1[27]_o , i0[27], i1[27]);
  xor \xor_i0[28]_i1[28]  (\xor_i0[28]_i1[28]_o , i0[28], i1[28]);
  xor \xor_i0[29]_i1[29]  (\xor_i0[29]_i1[29]_o , i0[29], i1[29]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[30]_i1[30]  (\xor_i0[30]_i1[30]_o , i0[30], i1[30]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module lt_u32_u32
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [31:0] i0;
  input [31:0] i1;
  output o;

  wire [31:0] diff;
  wire diff_12_18;
  wire diff_19_26;
  wire diff_27_31;
  wire diff_6_11;
  wire less_12_18;
  wire \less_12_18_inst/diff_0 ;
  wire \less_12_18_inst/diff_1 ;
  wire \less_12_18_inst/diff_2 ;
  wire \less_12_18_inst/diff_3 ;
  wire \less_12_18_inst/diff_4 ;
  wire \less_12_18_inst/diff_5 ;
  wire \less_12_18_inst/diff_6 ;
  wire \less_12_18_inst/o_0 ;
  wire \less_12_18_inst/o_1 ;
  wire \less_12_18_inst/o_2 ;
  wire \less_12_18_inst/o_3 ;
  wire \less_12_18_inst/o_4 ;
  wire \less_12_18_inst/o_5 ;
  wire less_19_26;
  wire \less_19_26_inst/diff_0 ;
  wire \less_19_26_inst/diff_1 ;
  wire \less_19_26_inst/diff_2 ;
  wire \less_19_26_inst/diff_3 ;
  wire \less_19_26_inst/diff_4 ;
  wire \less_19_26_inst/diff_5 ;
  wire \less_19_26_inst/diff_6 ;
  wire \less_19_26_inst/diff_7 ;
  wire \less_19_26_inst/o_0 ;
  wire \less_19_26_inst/o_1 ;
  wire \less_19_26_inst/o_2 ;
  wire \less_19_26_inst/o_3 ;
  wire \less_19_26_inst/o_4 ;
  wire \less_19_26_inst/o_5 ;
  wire \less_19_26_inst/o_6 ;
  wire less_27_31;
  wire \less_27_31_inst/diff_0 ;
  wire \less_27_31_inst/diff_1 ;
  wire \less_27_31_inst/diff_2 ;
  wire \less_27_31_inst/diff_3 ;
  wire \less_27_31_inst/diff_4 ;
  wire \less_27_31_inst/o_0 ;
  wire \less_27_31_inst/o_1 ;
  wire \less_27_31_inst/o_2 ;
  wire \less_27_31_inst/o_3 ;
  wire less_6_11;
  wire \less_6_11_inst/diff_0 ;
  wire \less_6_11_inst/diff_1 ;
  wire \less_6_11_inst/diff_2 ;
  wire \less_6_11_inst/diff_3 ;
  wire \less_6_11_inst/diff_4 ;
  wire \less_6_11_inst/diff_5 ;
  wire \less_6_11_inst/o_0 ;
  wire \less_6_11_inst/o_1 ;
  wire \less_6_11_inst/o_2 ;
  wire \less_6_11_inst/o_3 ;
  wire \less_6_11_inst/o_4 ;
  wire o_0;
  wire o_1;
  wire o_2;
  wire o_3;
  wire o_4;
  wire o_5;
  wire o_6;
  wire o_7;
  wire o_8;

  or any_diff_12_18 (diff_12_18, diff[12], diff[13], diff[14], diff[15], diff[16], diff[17], diff[18]);
  or any_diff_19_26 (diff_19_26, diff[19], diff[20], diff[21], diff[22], diff[23], diff[24], diff[25], diff[26]);
  or any_diff_27_31 (diff_27_31, diff[27], diff[28], diff[29], diff[30], diff[31]);
  or any_diff_6_11 (diff_6_11, diff[6], diff[7], diff[8], diff[9], diff[10], diff[11]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_12 (diff[12], i0[12], i1[12]);
  xor diff_13 (diff[13], i0[13], i1[13]);
  xor diff_14 (diff[14], i0[14], i1[14]);
  xor diff_15 (diff[15], i0[15], i1[15]);
  xor diff_16 (diff[16], i0[16], i1[16]);
  xor diff_17 (diff[17], i0[17], i1[17]);
  xor diff_18 (diff[18], i0[18], i1[18]);
  xor diff_19 (diff[19], i0[19], i1[19]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_20 (diff[20], i0[20], i1[20]);
  xor diff_21 (diff[21], i0[21], i1[21]);
  xor diff_22 (diff[22], i0[22], i1[22]);
  xor diff_23 (diff[23], i0[23], i1[23]);
  xor diff_24 (diff[24], i0[24], i1[24]);
  xor diff_25 (diff[25], i0[25], i1[25]);
  xor diff_26 (diff[26], i0[26], i1[26]);
  xor diff_27 (diff[27], i0[27], i1[27]);
  xor diff_28 (diff[28], i0[28], i1[28]);
  xor diff_29 (diff[29], i0[29], i1[29]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_30 (diff[30], i0[30], i1[30]);
  xor diff_31 (diff[31], i0[31], i1[31]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);
  AL_MUX \less_12_18_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[12]),
    .sel(\less_12_18_inst/diff_0 ),
    .o(\less_12_18_inst/o_0 ));
  AL_MUX \less_12_18_inst/mux_1  (
    .i0(\less_12_18_inst/o_0 ),
    .i1(i1[13]),
    .sel(\less_12_18_inst/diff_1 ),
    .o(\less_12_18_inst/o_1 ));
  AL_MUX \less_12_18_inst/mux_2  (
    .i0(\less_12_18_inst/o_1 ),
    .i1(i1[14]),
    .sel(\less_12_18_inst/diff_2 ),
    .o(\less_12_18_inst/o_2 ));
  AL_MUX \less_12_18_inst/mux_3  (
    .i0(\less_12_18_inst/o_2 ),
    .i1(i1[15]),
    .sel(\less_12_18_inst/diff_3 ),
    .o(\less_12_18_inst/o_3 ));
  AL_MUX \less_12_18_inst/mux_4  (
    .i0(\less_12_18_inst/o_3 ),
    .i1(i1[16]),
    .sel(\less_12_18_inst/diff_4 ),
    .o(\less_12_18_inst/o_4 ));
  AL_MUX \less_12_18_inst/mux_5  (
    .i0(\less_12_18_inst/o_4 ),
    .i1(i1[17]),
    .sel(\less_12_18_inst/diff_5 ),
    .o(\less_12_18_inst/o_5 ));
  AL_MUX \less_12_18_inst/mux_6  (
    .i0(\less_12_18_inst/o_5 ),
    .i1(i1[18]),
    .sel(\less_12_18_inst/diff_6 ),
    .o(less_12_18));
  xor \less_12_18_inst/xor_0  (\less_12_18_inst/diff_0 , i0[12], i1[12]);
  xor \less_12_18_inst/xor_1  (\less_12_18_inst/diff_1 , i0[13], i1[13]);
  xor \less_12_18_inst/xor_2  (\less_12_18_inst/diff_2 , i0[14], i1[14]);
  xor \less_12_18_inst/xor_3  (\less_12_18_inst/diff_3 , i0[15], i1[15]);
  xor \less_12_18_inst/xor_4  (\less_12_18_inst/diff_4 , i0[16], i1[16]);
  xor \less_12_18_inst/xor_5  (\less_12_18_inst/diff_5 , i0[17], i1[17]);
  xor \less_12_18_inst/xor_6  (\less_12_18_inst/diff_6 , i0[18], i1[18]);
  AL_MUX \less_19_26_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[19]),
    .sel(\less_19_26_inst/diff_0 ),
    .o(\less_19_26_inst/o_0 ));
  AL_MUX \less_19_26_inst/mux_1  (
    .i0(\less_19_26_inst/o_0 ),
    .i1(i1[20]),
    .sel(\less_19_26_inst/diff_1 ),
    .o(\less_19_26_inst/o_1 ));
  AL_MUX \less_19_26_inst/mux_2  (
    .i0(\less_19_26_inst/o_1 ),
    .i1(i1[21]),
    .sel(\less_19_26_inst/diff_2 ),
    .o(\less_19_26_inst/o_2 ));
  AL_MUX \less_19_26_inst/mux_3  (
    .i0(\less_19_26_inst/o_2 ),
    .i1(i1[22]),
    .sel(\less_19_26_inst/diff_3 ),
    .o(\less_19_26_inst/o_3 ));
  AL_MUX \less_19_26_inst/mux_4  (
    .i0(\less_19_26_inst/o_3 ),
    .i1(i1[23]),
    .sel(\less_19_26_inst/diff_4 ),
    .o(\less_19_26_inst/o_4 ));
  AL_MUX \less_19_26_inst/mux_5  (
    .i0(\less_19_26_inst/o_4 ),
    .i1(i1[24]),
    .sel(\less_19_26_inst/diff_5 ),
    .o(\less_19_26_inst/o_5 ));
  AL_MUX \less_19_26_inst/mux_6  (
    .i0(\less_19_26_inst/o_5 ),
    .i1(i1[25]),
    .sel(\less_19_26_inst/diff_6 ),
    .o(\less_19_26_inst/o_6 ));
  AL_MUX \less_19_26_inst/mux_7  (
    .i0(\less_19_26_inst/o_6 ),
    .i1(i1[26]),
    .sel(\less_19_26_inst/diff_7 ),
    .o(less_19_26));
  xor \less_19_26_inst/xor_0  (\less_19_26_inst/diff_0 , i0[19], i1[19]);
  xor \less_19_26_inst/xor_1  (\less_19_26_inst/diff_1 , i0[20], i1[20]);
  xor \less_19_26_inst/xor_2  (\less_19_26_inst/diff_2 , i0[21], i1[21]);
  xor \less_19_26_inst/xor_3  (\less_19_26_inst/diff_3 , i0[22], i1[22]);
  xor \less_19_26_inst/xor_4  (\less_19_26_inst/diff_4 , i0[23], i1[23]);
  xor \less_19_26_inst/xor_5  (\less_19_26_inst/diff_5 , i0[24], i1[24]);
  xor \less_19_26_inst/xor_6  (\less_19_26_inst/diff_6 , i0[25], i1[25]);
  xor \less_19_26_inst/xor_7  (\less_19_26_inst/diff_7 , i0[26], i1[26]);
  AL_MUX \less_27_31_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[27]),
    .sel(\less_27_31_inst/diff_0 ),
    .o(\less_27_31_inst/o_0 ));
  AL_MUX \less_27_31_inst/mux_1  (
    .i0(\less_27_31_inst/o_0 ),
    .i1(i1[28]),
    .sel(\less_27_31_inst/diff_1 ),
    .o(\less_27_31_inst/o_1 ));
  AL_MUX \less_27_31_inst/mux_2  (
    .i0(\less_27_31_inst/o_1 ),
    .i1(i1[29]),
    .sel(\less_27_31_inst/diff_2 ),
    .o(\less_27_31_inst/o_2 ));
  AL_MUX \less_27_31_inst/mux_3  (
    .i0(\less_27_31_inst/o_2 ),
    .i1(i1[30]),
    .sel(\less_27_31_inst/diff_3 ),
    .o(\less_27_31_inst/o_3 ));
  AL_MUX \less_27_31_inst/mux_4  (
    .i0(\less_27_31_inst/o_3 ),
    .i1(i1[31]),
    .sel(\less_27_31_inst/diff_4 ),
    .o(less_27_31));
  xor \less_27_31_inst/xor_0  (\less_27_31_inst/diff_0 , i0[27], i1[27]);
  xor \less_27_31_inst/xor_1  (\less_27_31_inst/diff_1 , i0[28], i1[28]);
  xor \less_27_31_inst/xor_2  (\less_27_31_inst/diff_2 , i0[29], i1[29]);
  xor \less_27_31_inst/xor_3  (\less_27_31_inst/diff_3 , i0[30], i1[30]);
  xor \less_27_31_inst/xor_4  (\less_27_31_inst/diff_4 , i0[31], i1[31]);
  AL_MUX \less_6_11_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[6]),
    .sel(\less_6_11_inst/diff_0 ),
    .o(\less_6_11_inst/o_0 ));
  AL_MUX \less_6_11_inst/mux_1  (
    .i0(\less_6_11_inst/o_0 ),
    .i1(i1[7]),
    .sel(\less_6_11_inst/diff_1 ),
    .o(\less_6_11_inst/o_1 ));
  AL_MUX \less_6_11_inst/mux_2  (
    .i0(\less_6_11_inst/o_1 ),
    .i1(i1[8]),
    .sel(\less_6_11_inst/diff_2 ),
    .o(\less_6_11_inst/o_2 ));
  AL_MUX \less_6_11_inst/mux_3  (
    .i0(\less_6_11_inst/o_2 ),
    .i1(i1[9]),
    .sel(\less_6_11_inst/diff_3 ),
    .o(\less_6_11_inst/o_3 ));
  AL_MUX \less_6_11_inst/mux_4  (
    .i0(\less_6_11_inst/o_3 ),
    .i1(i1[10]),
    .sel(\less_6_11_inst/diff_4 ),
    .o(\less_6_11_inst/o_4 ));
  AL_MUX \less_6_11_inst/mux_5  (
    .i0(\less_6_11_inst/o_4 ),
    .i1(i1[11]),
    .sel(\less_6_11_inst/diff_5 ),
    .o(less_6_11));
  xor \less_6_11_inst/xor_0  (\less_6_11_inst/diff_0 , i0[6], i1[6]);
  xor \less_6_11_inst/xor_1  (\less_6_11_inst/diff_1 , i0[7], i1[7]);
  xor \less_6_11_inst/xor_2  (\less_6_11_inst/diff_2 , i0[8], i1[8]);
  xor \less_6_11_inst/xor_3  (\less_6_11_inst/diff_3 , i0[9], i1[9]);
  xor \less_6_11_inst/xor_4  (\less_6_11_inst/diff_4 , i0[10], i1[10]);
  xor \less_6_11_inst/xor_5  (\less_6_11_inst/diff_5 , i0[11], i1[11]);
  AL_MUX mux_0 (
    .i0(ci),
    .i1(i1[0]),
    .sel(diff[0]),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(i1[1]),
    .sel(diff[1]),
    .o(o_1));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(i1[2]),
    .sel(diff[2]),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(i1[3]),
    .sel(diff[3]),
    .o(o_3));
  AL_MUX mux_4 (
    .i0(o_3),
    .i1(i1[4]),
    .sel(diff[4]),
    .o(o_4));
  AL_MUX mux_5 (
    .i0(o_4),
    .i1(i1[5]),
    .sel(diff[5]),
    .o(o_5));
  AL_MUX mux_6 (
    .i0(o_5),
    .i1(less_6_11),
    .sel(diff_6_11),
    .o(o_6));
  AL_MUX mux_7 (
    .i0(o_6),
    .i1(less_12_18),
    .sel(diff_12_18),
    .o(o_7));
  AL_MUX mux_8 (
    .i0(o_7),
    .i1(less_19_26),
    .sel(diff_19_26),
    .o(o_8));
  AL_MUX mux_9 (
    .i0(o_8),
    .i1(less_27_31),
    .sel(diff_27_31),
    .o(o));

endmodule 

module lt_u13_u13
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [12:0] i0;
  input [12:0] i1;
  output o;

  wire [12:0] diff;
  wire diff_6_11;
  wire less_6_11;
  wire \less_6_11_inst/diff_0 ;
  wire \less_6_11_inst/diff_1 ;
  wire \less_6_11_inst/diff_2 ;
  wire \less_6_11_inst/diff_3 ;
  wire \less_6_11_inst/diff_4 ;
  wire \less_6_11_inst/diff_5 ;
  wire \less_6_11_inst/o_0 ;
  wire \less_6_11_inst/o_1 ;
  wire \less_6_11_inst/o_2 ;
  wire \less_6_11_inst/o_3 ;
  wire \less_6_11_inst/o_4 ;
  wire o_0;
  wire o_1;
  wire o_2;
  wire o_3;
  wire o_4;
  wire o_5;
  wire o_6;

  or any_diff_6_11 (diff_6_11, diff[6], diff[7], diff[8], diff[9], diff[10], diff[11]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_12 (diff[12], i0[12], i1[12]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);
  AL_MUX \less_6_11_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[6]),
    .sel(\less_6_11_inst/diff_0 ),
    .o(\less_6_11_inst/o_0 ));
  AL_MUX \less_6_11_inst/mux_1  (
    .i0(\less_6_11_inst/o_0 ),
    .i1(i1[7]),
    .sel(\less_6_11_inst/diff_1 ),
    .o(\less_6_11_inst/o_1 ));
  AL_MUX \less_6_11_inst/mux_2  (
    .i0(\less_6_11_inst/o_1 ),
    .i1(i1[8]),
    .sel(\less_6_11_inst/diff_2 ),
    .o(\less_6_11_inst/o_2 ));
  AL_MUX \less_6_11_inst/mux_3  (
    .i0(\less_6_11_inst/o_2 ),
    .i1(i1[9]),
    .sel(\less_6_11_inst/diff_3 ),
    .o(\less_6_11_inst/o_3 ));
  AL_MUX \less_6_11_inst/mux_4  (
    .i0(\less_6_11_inst/o_3 ),
    .i1(i1[10]),
    .sel(\less_6_11_inst/diff_4 ),
    .o(\less_6_11_inst/o_4 ));
  AL_MUX \less_6_11_inst/mux_5  (
    .i0(\less_6_11_inst/o_4 ),
    .i1(i1[11]),
    .sel(\less_6_11_inst/diff_5 ),
    .o(less_6_11));
  xor \less_6_11_inst/xor_0  (\less_6_11_inst/diff_0 , i0[6], i1[6]);
  xor \less_6_11_inst/xor_1  (\less_6_11_inst/diff_1 , i0[7], i1[7]);
  xor \less_6_11_inst/xor_2  (\less_6_11_inst/diff_2 , i0[8], i1[8]);
  xor \less_6_11_inst/xor_3  (\less_6_11_inst/diff_3 , i0[9], i1[9]);
  xor \less_6_11_inst/xor_4  (\less_6_11_inst/diff_4 , i0[10], i1[10]);
  xor \less_6_11_inst/xor_5  (\less_6_11_inst/diff_5 , i0[11], i1[11]);
  AL_MUX mux_0 (
    .i0(ci),
    .i1(i1[0]),
    .sel(diff[0]),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(i1[1]),
    .sel(diff[1]),
    .o(o_1));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(i1[2]),
    .sel(diff[2]),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(i1[3]),
    .sel(diff[3]),
    .o(o_3));
  AL_MUX mux_4 (
    .i0(o_3),
    .i1(i1[4]),
    .sel(diff[4]),
    .o(o_4));
  AL_MUX mux_5 (
    .i0(o_4),
    .i1(i1[5]),
    .sel(diff[5]),
    .o(o_5));
  AL_MUX mux_6 (
    .i0(o_5),
    .i1(less_6_11),
    .sel(diff_6_11),
    .o(o_6));
  AL_MUX mux_7 (
    .i0(o_6),
    .i1(i1[12]),
    .sel(diff[12]),
    .o(o));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module add_pu11_mu11_o12
  (
  i0,
  i1,
  o
  );

  input [10:0] i0;
  input [10:0] i1;
  output [11:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_nb0;
  wire net_nb1;
  wire net_nb10;
  wire net_nb2;
  wire net_nb3;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_nb9;
  wire net_ncout;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[11] = net_ncout;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_nb10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_nb9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b10 (net_nb10, net_b10);
  not inv_b2 (net_nb2, net_b2);
  not inv_b3 (net_nb3, net_b3);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);
  not inv_b9 (net_nb9, net_b9);
  not inv_cout (net_ncout, net_cout10);

endmodule 

module add_pu10_mu10_o11
  (
  i0,
  i1,
  o
  );

  input [9:0] i0;
  input [9:0] i1;
  output [10:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_nb0;
  wire net_nb1;
  wire net_nb2;
  wire net_nb3;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_nb9;
  wire net_ncout;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[10] = net_ncout;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_nb9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b2 (net_nb2, net_b2);
  not inv_b3 (net_nb3, net_b3);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);
  not inv_b9 (net_nb9, net_b9);
  not inv_cout (net_ncout, net_cout9);

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_FADD
  (
  input a,
  input b,
  input c,
  output sum,
  output cout
  );

  wire prop;
  wire not_prop;
  wire sel_i0;
  wire sel_i1;

  xor u0 (prop, a, b);
  xor u1 (sum, prop, c);
  not u2 (not_prop, prop);
  and u3 (sel_i1, prop, c);
  and u4 (sel_i0, not_prop, a);
  or  u5 (cout, sel_i0, sel_i1);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  // synthesis translate_off
  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end
  // synthesis translate_on

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

