// Verilog netlist created by TD v5.0.19080
// Sun May 31 12:04:52 2020

`timescale 1ns / 1ps
module VGA_Demo  // source/rtl/VGA_Demo.v(2)
  (
  clk_24m,
  on_off,
  rst_n,
  vga_b,
  vga_clk,
  vga_de,
  vga_g,
  vga_hs,
  vga_r,
  vga_vs
  );

  input clk_24m;  // source/rtl/VGA_Demo.v(4)
  input [7:0] on_off;  // source/rtl/VGA_Demo.v(6)
  input rst_n;  // source/rtl/VGA_Demo.v(5)
  output [7:0] vga_b;  // source/rtl/VGA_Demo.v(17)
  output vga_clk;  // source/rtl/VGA_Demo.v(9)
  output vga_de;  // source/rtl/VGA_Demo.v(13)
  output [7:0] vga_g;  // source/rtl/VGA_Demo.v(16)
  output vga_hs;  // source/rtl/VGA_Demo.v(10)
  output [7:0] vga_r;  // source/rtl/VGA_Demo.v(15)
  output vga_vs;  // source/rtl/VGA_Demo.v(11)

  wire [23:0] lcd_data;  // source/rtl/VGA_Demo.v(23)
  wire [11:0] lcd_xpos;  // source/rtl/VGA_Demo.v(21)
  wire [11:0] lcd_ypos;  // source/rtl/VGA_Demo.v(22)
  wire [7:0] on_off_pad;  // source/rtl/VGA_Demo.v(6)
  wire [11:0] \u1_Driver/hcnt ;  // source/rtl/Driver.v(44)
  wire [11:0] \u1_Driver/n2 ;
  wire [12:0] \u1_Driver/n20 ;
  wire [12:0] \u1_Driver/n21 ;
  wire [11:0] \u1_Driver/n3 ;
  wire [11:0] \u1_Driver/n7 ;
  wire [11:0] \u1_Driver/n8 ;
  wire [11:0] \u1_Driver/vcnt ;  // source/rtl/Driver.v(45)
  wire [31:0] \u2_Display/counta ;  // source/rtl/Display.v(39)
  wire [31:0] \u2_Display/i ;  // source/rtl/Display.v(41)
  wire [31:0] \u2_Display/j ;  // source/rtl/Display.v(42)
  wire [30:0] \u2_Display/n ;  // source/rtl/Display.v(48)
  wire [31:0] \u2_Display/n1014 ;
  wire [31:0] \u2_Display/n102 ;
  wire [31:0] \u2_Display/n1049 ;
  wire [31:0] \u2_Display/n1084 ;
  wire [31:0] \u2_Display/n1119 ;
  wire [31:0] \u2_Display/n1154 ;
  wire [31:0] \u2_Display/n1189 ;
  wire [24:0] \u2_Display/n135 ;
  wire [31:0] \u2_Display/n137 ;
  wire [22:0] \u2_Display/n140 ;
  wire [31:0] \u2_Display/n143 ;
  wire [31:0] \u2_Display/n1542 ;
  wire [31:0] \u2_Display/n1577 ;
  wire [31:0] \u2_Display/n1612 ;
  wire [31:0] \u2_Display/n1647 ;
  wire [31:0] \u2_Display/n1682 ;
  wire [31:0] \u2_Display/n1717 ;
  wire [31:0] \u2_Display/n1752 ;
  wire [31:0] \u2_Display/n1787 ;
  wire [31:0] \u2_Display/n1822 ;
  wire [31:0] \u2_Display/n1857 ;
  wire [31:0] \u2_Display/n1892 ;
  wire [31:0] \u2_Display/n1927 ;
  wire [31:0] \u2_Display/n1962 ;
  wire [31:0] \u2_Display/n1997 ;
  wire [31:0] \u2_Display/n2032 ;
  wire [31:0] \u2_Display/n2067 ;
  wire [31:0] \u2_Display/n2102 ;
  wire [31:0] \u2_Display/n2137 ;
  wire [31:0] \u2_Display/n2172 ;
  wire [31:0] \u2_Display/n2207 ;
  wire [31:0] \u2_Display/n2242 ;
  wire [31:0] \u2_Display/n2277 ;
  wire [31:0] \u2_Display/n2312 ;
  wire [23:0] \u2_Display/n236 ;
  wire [31:0] \u2_Display/n238 ;
  wire [31:0] \u2_Display/n239 ;
  wire [23:0] \u2_Display/n240 ;
  wire [31:0] \u2_Display/n2665 ;
  wire [31:0] \u2_Display/n2700 ;
  wire [31:0] \u2_Display/n2735 ;
  wire [31:0] \u2_Display/n2770 ;
  wire [31:0] \u2_Display/n2805 ;
  wire [31:0] \u2_Display/n2840 ;
  wire [31:0] \u2_Display/n2875 ;
  wire [31:0] \u2_Display/n2910 ;
  wire [31:0] \u2_Display/n2945 ;
  wire [31:0] \u2_Display/n2980 ;
  wire [31:0] \u2_Display/n3015 ;
  wire [31:0] \u2_Display/n3050 ;
  wire [31:0] \u2_Display/n3085 ;
  wire [31:0] \u2_Display/n3120 ;
  wire [31:0] \u2_Display/n3155 ;
  wire [31:0] \u2_Display/n3190 ;
  wire [31:0] \u2_Display/n3225 ;
  wire [31:0] \u2_Display/n3260 ;
  wire [31:0] \u2_Display/n3295 ;
  wire [31:0] \u2_Display/n3330 ;
  wire [31:0] \u2_Display/n3365 ;
  wire [31:0] \u2_Display/n3400 ;
  wire [31:0] \u2_Display/n3435 ;
  wire [30:0] \u2_Display/n37 ;
  wire [31:0] \u2_Display/n3788 ;
  wire [31:0] \u2_Display/n3823 ;
  wire [31:0] \u2_Display/n3858 ;
  wire [31:0] \u2_Display/n3893 ;
  wire [31:0] \u2_Display/n3928 ;
  wire [31:0] \u2_Display/n3963 ;
  wire [31:0] \u2_Display/n3998 ;
  wire [31:0] \u2_Display/n4033 ;
  wire [31:0] \u2_Display/n4068 ;
  wire [31:0] \u2_Display/n41 ;
  wire [31:0] \u2_Display/n4103 ;
  wire [31:0] \u2_Display/n4138 ;
  wire [31:0] \u2_Display/n4173 ;
  wire [31:0] \u2_Display/n419 ;
  wire [31:0] \u2_Display/n4208 ;
  wire [31:0] \u2_Display/n4243 ;
  wire [31:0] \u2_Display/n4278 ;
  wire [23:0] \u2_Display/n43 ;
  wire [31:0] \u2_Display/n4313 ;
  wire [31:0] \u2_Display/n4348 ;
  wire [31:0] \u2_Display/n4383 ;
  wire [31:0] \u2_Display/n4418 ;
  wire [31:0] \u2_Display/n4453 ;
  wire [31:0] \u2_Display/n4488 ;
  wire [31:0] \u2_Display/n4523 ;
  wire [31:0] \u2_Display/n454 ;
  wire [31:0] \u2_Display/n4558 ;
  wire [31:0] \u2_Display/n489 ;
  wire [31:0] \u2_Display/n4911 ;
  wire [31:0] \u2_Display/n4946 ;
  wire [31:0] \u2_Display/n4981 ;
  wire [31:0] \u2_Display/n5016 ;
  wire [31:0] \u2_Display/n5051 ;
  wire [31:0] \u2_Display/n5086 ;
  wire [31:0] \u2_Display/n5121 ;
  wire [31:0] \u2_Display/n5156 ;
  wire [31:0] \u2_Display/n5191 ;
  wire [31:0] \u2_Display/n5226 ;
  wire [31:0] \u2_Display/n524 ;
  wire [31:0] \u2_Display/n5261 ;
  wire [31:0] \u2_Display/n5296 ;
  wire [31:0] \u2_Display/n5331 ;
  wire [31:0] \u2_Display/n5366 ;
  wire [31:0] \u2_Display/n5401 ;
  wire [31:0] \u2_Display/n5436 ;
  wire [31:0] \u2_Display/n5471 ;
  wire [31:0] \u2_Display/n5506 ;
  wire [31:0] \u2_Display/n5541 ;
  wire [31:0] \u2_Display/n5576 ;
  wire [31:0] \u2_Display/n559 ;
  wire [31:0] \u2_Display/n5611 ;
  wire [31:0] \u2_Display/n5646 ;
  wire [31:0] \u2_Display/n5681 ;
  wire [31:0] \u2_Display/n594 ;
  wire [31:0] \u2_Display/n629 ;
  wire [31:0] \u2_Display/n664 ;
  wire [31:0] \u2_Display/n699 ;
  wire [31:0] \u2_Display/n734 ;
  wire [31:0] \u2_Display/n769 ;
  wire [31:0] \u2_Display/n804 ;
  wire [31:0] \u2_Display/n839 ;
  wire [31:0] \u2_Display/n874 ;
  wire [31:0] \u2_Display/n909 ;
  wire [24:0] \u2_Display/n94 ;
  wire [31:0] \u2_Display/n944 ;
  wire [31:0] \u2_Display/n96 ;
  wire [31:0] \u2_Display/n979 ;
  wire [22:0] \u2_Display/n99 ;
  wire [7:0] vga_b_pad;  // source/rtl/VGA_Demo.v(17)
  wire _al_u1168_o;
  wire _al_u1170_o;
  wire _al_u1171_o;
  wire _al_u1345_o;
  wire _al_u1346_o;
  wire _al_u1347_o;
  wire _al_u1348_o;
  wire _al_u1349_o;
  wire _al_u1350_o;
  wire _al_u1351_o;
  wire _al_u1352_o;
  wire _al_u1353_o;
  wire _al_u3916_o;
  wire _al_u3917_o;
  wire _al_u3918_o;
  wire _al_u3920_o;
  wire _al_u3921_o;
  wire _al_u3922_o;
  wire _al_u3924_o;
  wire _al_u3925_o;
  wire _al_u3926_o;
  wire _al_u3928_o;
  wire _al_u3929_o;
  wire _al_u3930_o;
  wire _al_u3932_o;
  wire _al_u3933_o;
  wire _al_u3934_o;
  wire _al_u3936_o;
  wire _al_u3937_o;
  wire _al_u3938_o;
  wire _al_u3940_o;
  wire _al_u3941_o;
  wire _al_u3942_o;
  wire _al_u3944_o;
  wire _al_u3945_o;
  wire _al_u3946_o;
  wire _al_u3948_o;
  wire _al_u3949_o;
  wire _al_u3950_o;
  wire _al_u3952_o;
  wire _al_u3953_o;
  wire _al_u3954_o;
  wire _al_u3956_o;
  wire _al_u3957_o;
  wire _al_u3958_o;
  wire _al_u3960_o;
  wire _al_u3961_o;
  wire _al_u3962_o;
  wire _al_u3963_o;
  wire _al_u3965_o;
  wire _al_u3966_o;
  wire _al_u3967_o;
  wire _al_u3969_o;
  wire _al_u3970_o;
  wire _al_u3971_o;
  wire _al_u3972_o;
  wire _al_u3974_o;
  wire _al_u3975_o;
  wire _al_u3976_o;
  wire _al_u3978_o;
  wire _al_u3979_o;
  wire _al_u3980_o;
  wire _al_u3981_o;
  wire _al_u3983_o;
  wire _al_u3984_o;
  wire _al_u3985_o;
  wire _al_u3987_o;
  wire _al_u3988_o;
  wire _al_u3989_o;
  wire _al_u3991_o;
  wire _al_u3992_o;
  wire _al_u3993_o;
  wire _al_u3995_o;
  wire _al_u3996_o;
  wire _al_u3997_o;
  wire _al_u997_o;
  wire _al_u998_o;
  wire clk_24m_pad;  // source/rtl/VGA_Demo.v(4)
  wire clk_vga;  // source/rtl/VGA_Demo.v(20)
  wire rst_n_pad;  // source/rtl/VGA_Demo.v(5)
  wire \u0_PLL/n0 ;
  wire \u0_PLL/uut/clk0_buf ;  // al_ip/PLL.v(32)
  wire \u1_Driver/add0/c0 ;
  wire \u1_Driver/add0/c1 ;
  wire \u1_Driver/add0/c10 ;
  wire \u1_Driver/add0/c11 ;
  wire \u1_Driver/add0/c2 ;
  wire \u1_Driver/add0/c3 ;
  wire \u1_Driver/add0/c4 ;
  wire \u1_Driver/add0/c5 ;
  wire \u1_Driver/add0/c6 ;
  wire \u1_Driver/add0/c7 ;
  wire \u1_Driver/add0/c8 ;
  wire \u1_Driver/add0/c9 ;
  wire \u1_Driver/add1/c0 ;
  wire \u1_Driver/add1/c1 ;
  wire \u1_Driver/add1/c10 ;
  wire \u1_Driver/add1/c11 ;
  wire \u1_Driver/add1/c2 ;
  wire \u1_Driver/add1/c3 ;
  wire \u1_Driver/add1/c4 ;
  wire \u1_Driver/add1/c5 ;
  wire \u1_Driver/add1/c6 ;
  wire \u1_Driver/add1/c7 ;
  wire \u1_Driver/add1/c8 ;
  wire \u1_Driver/add1/c9 ;
  wire \u1_Driver/lcd_request ;  // source/rtl/Driver.v(46)
  wire \u1_Driver/lt0_c0 ;
  wire \u1_Driver/lt0_c1 ;
  wire \u1_Driver/lt0_c10 ;
  wire \u1_Driver/lt0_c11 ;
  wire \u1_Driver/lt0_c12 ;
  wire \u1_Driver/lt0_c2 ;
  wire \u1_Driver/lt0_c3 ;
  wire \u1_Driver/lt0_c4 ;
  wire \u1_Driver/lt0_c5 ;
  wire \u1_Driver/lt0_c6 ;
  wire \u1_Driver/lt0_c7 ;
  wire \u1_Driver/lt0_c8 ;
  wire \u1_Driver/lt0_c9 ;
  wire \u1_Driver/lt1_c0 ;
  wire \u1_Driver/lt1_c1 ;
  wire \u1_Driver/lt1_c10 ;
  wire \u1_Driver/lt1_c11 ;
  wire \u1_Driver/lt1_c12 ;
  wire \u1_Driver/lt1_c2 ;
  wire \u1_Driver/lt1_c3 ;
  wire \u1_Driver/lt1_c4 ;
  wire \u1_Driver/lt1_c5 ;
  wire \u1_Driver/lt1_c6 ;
  wire \u1_Driver/lt1_c7 ;
  wire \u1_Driver/lt1_c8 ;
  wire \u1_Driver/lt1_c9 ;
  wire \u1_Driver/lt2_c0 ;
  wire \u1_Driver/lt2_c1 ;
  wire \u1_Driver/lt2_c10 ;
  wire \u1_Driver/lt2_c11 ;
  wire \u1_Driver/lt2_c12 ;
  wire \u1_Driver/lt2_c2 ;
  wire \u1_Driver/lt2_c3 ;
  wire \u1_Driver/lt2_c4 ;
  wire \u1_Driver/lt2_c5 ;
  wire \u1_Driver/lt2_c6 ;
  wire \u1_Driver/lt2_c7 ;
  wire \u1_Driver/lt2_c8 ;
  wire \u1_Driver/lt2_c9 ;
  wire \u1_Driver/lt3_c0 ;
  wire \u1_Driver/lt3_c1 ;
  wire \u1_Driver/lt3_c10 ;
  wire \u1_Driver/lt3_c11 ;
  wire \u1_Driver/lt3_c12 ;
  wire \u1_Driver/lt3_c2 ;
  wire \u1_Driver/lt3_c3 ;
  wire \u1_Driver/lt3_c4 ;
  wire \u1_Driver/lt3_c5 ;
  wire \u1_Driver/lt3_c6 ;
  wire \u1_Driver/lt3_c7 ;
  wire \u1_Driver/lt3_c8 ;
  wire \u1_Driver/lt3_c9 ;
  wire \u1_Driver/lt4_c0 ;
  wire \u1_Driver/lt4_c1 ;
  wire \u1_Driver/lt4_c10 ;
  wire \u1_Driver/lt4_c11 ;
  wire \u1_Driver/lt4_c12 ;
  wire \u1_Driver/lt4_c2 ;
  wire \u1_Driver/lt4_c3 ;
  wire \u1_Driver/lt4_c4 ;
  wire \u1_Driver/lt4_c5 ;
  wire \u1_Driver/lt4_c6 ;
  wire \u1_Driver/lt4_c7 ;
  wire \u1_Driver/lt4_c8 ;
  wire \u1_Driver/lt4_c9 ;
  wire \u1_Driver/lt5_c0 ;
  wire \u1_Driver/lt5_c1 ;
  wire \u1_Driver/lt5_c10 ;
  wire \u1_Driver/lt5_c11 ;
  wire \u1_Driver/lt5_c12 ;
  wire \u1_Driver/lt5_c2 ;
  wire \u1_Driver/lt5_c3 ;
  wire \u1_Driver/lt5_c4 ;
  wire \u1_Driver/lt5_c5 ;
  wire \u1_Driver/lt5_c6 ;
  wire \u1_Driver/lt5_c7 ;
  wire \u1_Driver/lt5_c8 ;
  wire \u1_Driver/lt5_c9 ;
  wire \u1_Driver/lt6_c0 ;
  wire \u1_Driver/lt6_c1 ;
  wire \u1_Driver/lt6_c10 ;
  wire \u1_Driver/lt6_c11 ;
  wire \u1_Driver/lt6_c12 ;
  wire \u1_Driver/lt6_c2 ;
  wire \u1_Driver/lt6_c3 ;
  wire \u1_Driver/lt6_c4 ;
  wire \u1_Driver/lt6_c5 ;
  wire \u1_Driver/lt6_c6 ;
  wire \u1_Driver/lt6_c7 ;
  wire \u1_Driver/lt6_c8 ;
  wire \u1_Driver/lt6_c9 ;
  wire \u1_Driver/lt7_c0 ;
  wire \u1_Driver/lt7_c1 ;
  wire \u1_Driver/lt7_c10 ;
  wire \u1_Driver/lt7_c11 ;
  wire \u1_Driver/lt7_c12 ;
  wire \u1_Driver/lt7_c2 ;
  wire \u1_Driver/lt7_c3 ;
  wire \u1_Driver/lt7_c4 ;
  wire \u1_Driver/lt7_c5 ;
  wire \u1_Driver/lt7_c6 ;
  wire \u1_Driver/lt7_c7 ;
  wire \u1_Driver/lt7_c8 ;
  wire \u1_Driver/lt7_c9 ;
  wire \u1_Driver/lt8_c0 ;
  wire \u1_Driver/lt8_c1 ;
  wire \u1_Driver/lt8_c10 ;
  wire \u1_Driver/lt8_c11 ;
  wire \u1_Driver/lt8_c12 ;
  wire \u1_Driver/lt8_c2 ;
  wire \u1_Driver/lt8_c3 ;
  wire \u1_Driver/lt8_c4 ;
  wire \u1_Driver/lt8_c5 ;
  wire \u1_Driver/lt8_c6 ;
  wire \u1_Driver/lt8_c7 ;
  wire \u1_Driver/lt8_c8 ;
  wire \u1_Driver/lt8_c9 ;
  wire \u1_Driver/n1 ;
  wire \u1_Driver/n10 ;
  wire \u1_Driver/n11 ;
  wire \u1_Driver/n12 ;
  wire \u1_Driver/n14 ;
  wire \u1_Driver/n15 ;
  wire \u1_Driver/n17 ;
  wire \u1_Driver/n18 ;
  wire \u1_Driver/n4 ;
  wire \u1_Driver/n5 ;
  wire \u1_Driver/n6_lutinv ;
  wire \u1_Driver/sub0/c0 ;
  wire \u1_Driver/sub0/c1 ;
  wire \u1_Driver/sub0/c10 ;
  wire \u1_Driver/sub0/c11 ;
  wire \u1_Driver/sub0/c2 ;
  wire \u1_Driver/sub0/c3 ;
  wire \u1_Driver/sub0/c4 ;
  wire \u1_Driver/sub0/c5 ;
  wire \u1_Driver/sub0/c6 ;
  wire \u1_Driver/sub0/c7 ;
  wire \u1_Driver/sub0/c8 ;
  wire \u1_Driver/sub0/c9 ;
  wire \u1_Driver/sub1/c0 ;
  wire \u1_Driver/sub1/c1 ;
  wire \u1_Driver/sub1/c10 ;
  wire \u1_Driver/sub1/c11 ;
  wire \u1_Driver/sub1/c2 ;
  wire \u1_Driver/sub1/c3 ;
  wire \u1_Driver/sub1/c4 ;
  wire \u1_Driver/sub1/c5 ;
  wire \u1_Driver/sub1/c6 ;
  wire \u1_Driver/sub1/c7 ;
  wire \u1_Driver/sub1/c8 ;
  wire \u1_Driver/sub1/c9 ;
  wire \u2_Display/add0/c0 ;
  wire \u2_Display/add0/c1 ;
  wire \u2_Display/add0/c10 ;
  wire \u2_Display/add0/c11 ;
  wire \u2_Display/add0/c12 ;
  wire \u2_Display/add0/c13 ;
  wire \u2_Display/add0/c14 ;
  wire \u2_Display/add0/c15 ;
  wire \u2_Display/add0/c16 ;
  wire \u2_Display/add0/c17 ;
  wire \u2_Display/add0/c18 ;
  wire \u2_Display/add0/c19 ;
  wire \u2_Display/add0/c2 ;
  wire \u2_Display/add0/c20 ;
  wire \u2_Display/add0/c21 ;
  wire \u2_Display/add0/c22 ;
  wire \u2_Display/add0/c23 ;
  wire \u2_Display/add0/c24 ;
  wire \u2_Display/add0/c25 ;
  wire \u2_Display/add0/c26 ;
  wire \u2_Display/add0/c27 ;
  wire \u2_Display/add0/c28 ;
  wire \u2_Display/add0/c29 ;
  wire \u2_Display/add0/c3 ;
  wire \u2_Display/add0/c30 ;
  wire \u2_Display/add0/c4 ;
  wire \u2_Display/add0/c5 ;
  wire \u2_Display/add0/c6 ;
  wire \u2_Display/add0/c7 ;
  wire \u2_Display/add0/c8 ;
  wire \u2_Display/add0/c9 ;
  wire \u2_Display/add1/c0 ;
  wire \u2_Display/add1/c1 ;
  wire \u2_Display/add1/c10 ;
  wire \u2_Display/add1/c11 ;
  wire \u2_Display/add1/c12 ;
  wire \u2_Display/add1/c13 ;
  wire \u2_Display/add1/c14 ;
  wire \u2_Display/add1/c15 ;
  wire \u2_Display/add1/c16 ;
  wire \u2_Display/add1/c17 ;
  wire \u2_Display/add1/c18 ;
  wire \u2_Display/add1/c19 ;
  wire \u2_Display/add1/c2 ;
  wire \u2_Display/add1/c20 ;
  wire \u2_Display/add1/c21 ;
  wire \u2_Display/add1/c22 ;
  wire \u2_Display/add1/c23 ;
  wire \u2_Display/add1/c24 ;
  wire \u2_Display/add1/c25 ;
  wire \u2_Display/add1/c26 ;
  wire \u2_Display/add1/c27 ;
  wire \u2_Display/add1/c28 ;
  wire \u2_Display/add1/c29 ;
  wire \u2_Display/add1/c3 ;
  wire \u2_Display/add1/c30 ;
  wire \u2_Display/add1/c31 ;
  wire \u2_Display/add1/c4 ;
  wire \u2_Display/add1/c5 ;
  wire \u2_Display/add1/c6 ;
  wire \u2_Display/add1/c7 ;
  wire \u2_Display/add1/c8 ;
  wire \u2_Display/add1/c9 ;
  wire \u2_Display/add100/c0 ;
  wire \u2_Display/add100/c1 ;
  wire \u2_Display/add100/c10 ;
  wire \u2_Display/add100/c11 ;
  wire \u2_Display/add100/c12 ;
  wire \u2_Display/add100/c13 ;
  wire \u2_Display/add100/c14 ;
  wire \u2_Display/add100/c15 ;
  wire \u2_Display/add100/c16 ;
  wire \u2_Display/add100/c17 ;
  wire \u2_Display/add100/c18 ;
  wire \u2_Display/add100/c19 ;
  wire \u2_Display/add100/c2 ;
  wire \u2_Display/add100/c20 ;
  wire \u2_Display/add100/c21 ;
  wire \u2_Display/add100/c22 ;
  wire \u2_Display/add100/c23 ;
  wire \u2_Display/add100/c24 ;
  wire \u2_Display/add100/c25 ;
  wire \u2_Display/add100/c26 ;
  wire \u2_Display/add100/c27 ;
  wire \u2_Display/add100/c28 ;
  wire \u2_Display/add100/c29 ;
  wire \u2_Display/add100/c3 ;
  wire \u2_Display/add100/c30 ;
  wire \u2_Display/add100/c31 ;
  wire \u2_Display/add100/c4 ;
  wire \u2_Display/add100/c5 ;
  wire \u2_Display/add100/c6 ;
  wire \u2_Display/add100/c7 ;
  wire \u2_Display/add100/c8 ;
  wire \u2_Display/add100/c9 ;
  wire \u2_Display/add101/c0 ;
  wire \u2_Display/add101/c1 ;
  wire \u2_Display/add101/c10 ;
  wire \u2_Display/add101/c11 ;
  wire \u2_Display/add101/c12 ;
  wire \u2_Display/add101/c13 ;
  wire \u2_Display/add101/c14 ;
  wire \u2_Display/add101/c15 ;
  wire \u2_Display/add101/c16 ;
  wire \u2_Display/add101/c17 ;
  wire \u2_Display/add101/c18 ;
  wire \u2_Display/add101/c19 ;
  wire \u2_Display/add101/c2 ;
  wire \u2_Display/add101/c20 ;
  wire \u2_Display/add101/c21 ;
  wire \u2_Display/add101/c22 ;
  wire \u2_Display/add101/c23 ;
  wire \u2_Display/add101/c24 ;
  wire \u2_Display/add101/c25 ;
  wire \u2_Display/add101/c26 ;
  wire \u2_Display/add101/c27 ;
  wire \u2_Display/add101/c28 ;
  wire \u2_Display/add101/c29 ;
  wire \u2_Display/add101/c3 ;
  wire \u2_Display/add101/c30 ;
  wire \u2_Display/add101/c31 ;
  wire \u2_Display/add101/c4 ;
  wire \u2_Display/add101/c5 ;
  wire \u2_Display/add101/c6 ;
  wire \u2_Display/add101/c7 ;
  wire \u2_Display/add101/c8 ;
  wire \u2_Display/add101/c9 ;
  wire \u2_Display/add102/c0 ;
  wire \u2_Display/add102/c1 ;
  wire \u2_Display/add102/c10 ;
  wire \u2_Display/add102/c11 ;
  wire \u2_Display/add102/c12 ;
  wire \u2_Display/add102/c13 ;
  wire \u2_Display/add102/c14 ;
  wire \u2_Display/add102/c15 ;
  wire \u2_Display/add102/c16 ;
  wire \u2_Display/add102/c17 ;
  wire \u2_Display/add102/c18 ;
  wire \u2_Display/add102/c19 ;
  wire \u2_Display/add102/c2 ;
  wire \u2_Display/add102/c20 ;
  wire \u2_Display/add102/c21 ;
  wire \u2_Display/add102/c22 ;
  wire \u2_Display/add102/c23 ;
  wire \u2_Display/add102/c24 ;
  wire \u2_Display/add102/c25 ;
  wire \u2_Display/add102/c26 ;
  wire \u2_Display/add102/c27 ;
  wire \u2_Display/add102/c28 ;
  wire \u2_Display/add102/c29 ;
  wire \u2_Display/add102/c3 ;
  wire \u2_Display/add102/c30 ;
  wire \u2_Display/add102/c31 ;
  wire \u2_Display/add102/c4 ;
  wire \u2_Display/add102/c5 ;
  wire \u2_Display/add102/c6 ;
  wire \u2_Display/add102/c7 ;
  wire \u2_Display/add102/c8 ;
  wire \u2_Display/add102/c9 ;
  wire \u2_Display/add103/c0 ;
  wire \u2_Display/add103/c1 ;
  wire \u2_Display/add103/c10 ;
  wire \u2_Display/add103/c11 ;
  wire \u2_Display/add103/c12 ;
  wire \u2_Display/add103/c13 ;
  wire \u2_Display/add103/c14 ;
  wire \u2_Display/add103/c15 ;
  wire \u2_Display/add103/c16 ;
  wire \u2_Display/add103/c17 ;
  wire \u2_Display/add103/c18 ;
  wire \u2_Display/add103/c19 ;
  wire \u2_Display/add103/c2 ;
  wire \u2_Display/add103/c20 ;
  wire \u2_Display/add103/c21 ;
  wire \u2_Display/add103/c22 ;
  wire \u2_Display/add103/c23 ;
  wire \u2_Display/add103/c24 ;
  wire \u2_Display/add103/c25 ;
  wire \u2_Display/add103/c26 ;
  wire \u2_Display/add103/c27 ;
  wire \u2_Display/add103/c28 ;
  wire \u2_Display/add103/c29 ;
  wire \u2_Display/add103/c3 ;
  wire \u2_Display/add103/c30 ;
  wire \u2_Display/add103/c31 ;
  wire \u2_Display/add103/c4 ;
  wire \u2_Display/add103/c5 ;
  wire \u2_Display/add103/c6 ;
  wire \u2_Display/add103/c7 ;
  wire \u2_Display/add103/c8 ;
  wire \u2_Display/add103/c9 ;
  wire \u2_Display/add104/c0 ;
  wire \u2_Display/add104/c1 ;
  wire \u2_Display/add104/c10 ;
  wire \u2_Display/add104/c11 ;
  wire \u2_Display/add104/c12 ;
  wire \u2_Display/add104/c13 ;
  wire \u2_Display/add104/c14 ;
  wire \u2_Display/add104/c15 ;
  wire \u2_Display/add104/c16 ;
  wire \u2_Display/add104/c17 ;
  wire \u2_Display/add104/c18 ;
  wire \u2_Display/add104/c19 ;
  wire \u2_Display/add104/c2 ;
  wire \u2_Display/add104/c20 ;
  wire \u2_Display/add104/c21 ;
  wire \u2_Display/add104/c22 ;
  wire \u2_Display/add104/c23 ;
  wire \u2_Display/add104/c24 ;
  wire \u2_Display/add104/c25 ;
  wire \u2_Display/add104/c26 ;
  wire \u2_Display/add104/c27 ;
  wire \u2_Display/add104/c28 ;
  wire \u2_Display/add104/c29 ;
  wire \u2_Display/add104/c3 ;
  wire \u2_Display/add104/c30 ;
  wire \u2_Display/add104/c31 ;
  wire \u2_Display/add104/c4 ;
  wire \u2_Display/add104/c5 ;
  wire \u2_Display/add104/c6 ;
  wire \u2_Display/add104/c7 ;
  wire \u2_Display/add104/c8 ;
  wire \u2_Display/add104/c9 ;
  wire \u2_Display/add105/c0 ;
  wire \u2_Display/add105/c1 ;
  wire \u2_Display/add105/c10 ;
  wire \u2_Display/add105/c11 ;
  wire \u2_Display/add105/c12 ;
  wire \u2_Display/add105/c13 ;
  wire \u2_Display/add105/c14 ;
  wire \u2_Display/add105/c15 ;
  wire \u2_Display/add105/c16 ;
  wire \u2_Display/add105/c17 ;
  wire \u2_Display/add105/c18 ;
  wire \u2_Display/add105/c19 ;
  wire \u2_Display/add105/c2 ;
  wire \u2_Display/add105/c20 ;
  wire \u2_Display/add105/c21 ;
  wire \u2_Display/add105/c22 ;
  wire \u2_Display/add105/c23 ;
  wire \u2_Display/add105/c24 ;
  wire \u2_Display/add105/c25 ;
  wire \u2_Display/add105/c26 ;
  wire \u2_Display/add105/c27 ;
  wire \u2_Display/add105/c28 ;
  wire \u2_Display/add105/c29 ;
  wire \u2_Display/add105/c3 ;
  wire \u2_Display/add105/c30 ;
  wire \u2_Display/add105/c31 ;
  wire \u2_Display/add105/c4 ;
  wire \u2_Display/add105/c5 ;
  wire \u2_Display/add105/c6 ;
  wire \u2_Display/add105/c7 ;
  wire \u2_Display/add105/c8 ;
  wire \u2_Display/add105/c9 ;
  wire \u2_Display/add106/c0 ;
  wire \u2_Display/add106/c1 ;
  wire \u2_Display/add106/c2 ;
  wire \u2_Display/add106/c3 ;
  wire \u2_Display/add106/c4 ;
  wire \u2_Display/add106/c5 ;
  wire \u2_Display/add106/c6 ;
  wire \u2_Display/add106/c7 ;
  wire \u2_Display/add106/c8 ;
  wire \u2_Display/add106/c9 ;
  wire \u2_Display/add117/c0 ;
  wire \u2_Display/add117/c1 ;
  wire \u2_Display/add117/c10 ;
  wire \u2_Display/add117/c11 ;
  wire \u2_Display/add117/c12 ;
  wire \u2_Display/add117/c13 ;
  wire \u2_Display/add117/c14 ;
  wire \u2_Display/add117/c15 ;
  wire \u2_Display/add117/c16 ;
  wire \u2_Display/add117/c17 ;
  wire \u2_Display/add117/c18 ;
  wire \u2_Display/add117/c19 ;
  wire \u2_Display/add117/c2 ;
  wire \u2_Display/add117/c20 ;
  wire \u2_Display/add117/c21 ;
  wire \u2_Display/add117/c22 ;
  wire \u2_Display/add117/c23 ;
  wire \u2_Display/add117/c24 ;
  wire \u2_Display/add117/c25 ;
  wire \u2_Display/add117/c26 ;
  wire \u2_Display/add117/c27 ;
  wire \u2_Display/add117/c28 ;
  wire \u2_Display/add117/c29 ;
  wire \u2_Display/add117/c3 ;
  wire \u2_Display/add117/c30 ;
  wire \u2_Display/add117/c31 ;
  wire \u2_Display/add117/c4 ;
  wire \u2_Display/add117/c5 ;
  wire \u2_Display/add117/c6 ;
  wire \u2_Display/add117/c7 ;
  wire \u2_Display/add117/c8 ;
  wire \u2_Display/add117/c9 ;
  wire \u2_Display/add118/c0 ;
  wire \u2_Display/add118/c1 ;
  wire \u2_Display/add118/c10 ;
  wire \u2_Display/add118/c11 ;
  wire \u2_Display/add118/c12 ;
  wire \u2_Display/add118/c13 ;
  wire \u2_Display/add118/c14 ;
  wire \u2_Display/add118/c15 ;
  wire \u2_Display/add118/c16 ;
  wire \u2_Display/add118/c17 ;
  wire \u2_Display/add118/c18 ;
  wire \u2_Display/add118/c19 ;
  wire \u2_Display/add118/c2 ;
  wire \u2_Display/add118/c20 ;
  wire \u2_Display/add118/c21 ;
  wire \u2_Display/add118/c22 ;
  wire \u2_Display/add118/c23 ;
  wire \u2_Display/add118/c24 ;
  wire \u2_Display/add118/c25 ;
  wire \u2_Display/add118/c26 ;
  wire \u2_Display/add118/c27 ;
  wire \u2_Display/add118/c28 ;
  wire \u2_Display/add118/c29 ;
  wire \u2_Display/add118/c3 ;
  wire \u2_Display/add118/c30 ;
  wire \u2_Display/add118/c31 ;
  wire \u2_Display/add118/c4 ;
  wire \u2_Display/add118/c5 ;
  wire \u2_Display/add118/c6 ;
  wire \u2_Display/add118/c7 ;
  wire \u2_Display/add118/c8 ;
  wire \u2_Display/add118/c9 ;
  wire \u2_Display/add119/c0 ;
  wire \u2_Display/add119/c1 ;
  wire \u2_Display/add119/c10 ;
  wire \u2_Display/add119/c11 ;
  wire \u2_Display/add119/c12 ;
  wire \u2_Display/add119/c13 ;
  wire \u2_Display/add119/c14 ;
  wire \u2_Display/add119/c15 ;
  wire \u2_Display/add119/c16 ;
  wire \u2_Display/add119/c17 ;
  wire \u2_Display/add119/c18 ;
  wire \u2_Display/add119/c19 ;
  wire \u2_Display/add119/c2 ;
  wire \u2_Display/add119/c20 ;
  wire \u2_Display/add119/c21 ;
  wire \u2_Display/add119/c22 ;
  wire \u2_Display/add119/c23 ;
  wire \u2_Display/add119/c24 ;
  wire \u2_Display/add119/c25 ;
  wire \u2_Display/add119/c26 ;
  wire \u2_Display/add119/c27 ;
  wire \u2_Display/add119/c28 ;
  wire \u2_Display/add119/c29 ;
  wire \u2_Display/add119/c3 ;
  wire \u2_Display/add119/c30 ;
  wire \u2_Display/add119/c31 ;
  wire \u2_Display/add119/c4 ;
  wire \u2_Display/add119/c5 ;
  wire \u2_Display/add119/c6 ;
  wire \u2_Display/add119/c7 ;
  wire \u2_Display/add119/c8 ;
  wire \u2_Display/add119/c9 ;
  wire \u2_Display/add120/c0 ;
  wire \u2_Display/add120/c1 ;
  wire \u2_Display/add120/c10 ;
  wire \u2_Display/add120/c11 ;
  wire \u2_Display/add120/c12 ;
  wire \u2_Display/add120/c13 ;
  wire \u2_Display/add120/c14 ;
  wire \u2_Display/add120/c15 ;
  wire \u2_Display/add120/c16 ;
  wire \u2_Display/add120/c17 ;
  wire \u2_Display/add120/c18 ;
  wire \u2_Display/add120/c19 ;
  wire \u2_Display/add120/c2 ;
  wire \u2_Display/add120/c20 ;
  wire \u2_Display/add120/c21 ;
  wire \u2_Display/add120/c22 ;
  wire \u2_Display/add120/c23 ;
  wire \u2_Display/add120/c24 ;
  wire \u2_Display/add120/c25 ;
  wire \u2_Display/add120/c26 ;
  wire \u2_Display/add120/c27 ;
  wire \u2_Display/add120/c28 ;
  wire \u2_Display/add120/c29 ;
  wire \u2_Display/add120/c3 ;
  wire \u2_Display/add120/c30 ;
  wire \u2_Display/add120/c31 ;
  wire \u2_Display/add120/c4 ;
  wire \u2_Display/add120/c5 ;
  wire \u2_Display/add120/c6 ;
  wire \u2_Display/add120/c7 ;
  wire \u2_Display/add120/c8 ;
  wire \u2_Display/add120/c9 ;
  wire \u2_Display/add121/c0 ;
  wire \u2_Display/add121/c1 ;
  wire \u2_Display/add121/c10 ;
  wire \u2_Display/add121/c11 ;
  wire \u2_Display/add121/c12 ;
  wire \u2_Display/add121/c13 ;
  wire \u2_Display/add121/c14 ;
  wire \u2_Display/add121/c15 ;
  wire \u2_Display/add121/c16 ;
  wire \u2_Display/add121/c17 ;
  wire \u2_Display/add121/c18 ;
  wire \u2_Display/add121/c19 ;
  wire \u2_Display/add121/c2 ;
  wire \u2_Display/add121/c20 ;
  wire \u2_Display/add121/c21 ;
  wire \u2_Display/add121/c22 ;
  wire \u2_Display/add121/c23 ;
  wire \u2_Display/add121/c24 ;
  wire \u2_Display/add121/c25 ;
  wire \u2_Display/add121/c26 ;
  wire \u2_Display/add121/c27 ;
  wire \u2_Display/add121/c28 ;
  wire \u2_Display/add121/c29 ;
  wire \u2_Display/add121/c3 ;
  wire \u2_Display/add121/c30 ;
  wire \u2_Display/add121/c31 ;
  wire \u2_Display/add121/c4 ;
  wire \u2_Display/add121/c5 ;
  wire \u2_Display/add121/c6 ;
  wire \u2_Display/add121/c7 ;
  wire \u2_Display/add121/c8 ;
  wire \u2_Display/add121/c9 ;
  wire \u2_Display/add122/c0 ;
  wire \u2_Display/add122/c1 ;
  wire \u2_Display/add122/c10 ;
  wire \u2_Display/add122/c11 ;
  wire \u2_Display/add122/c12 ;
  wire \u2_Display/add122/c13 ;
  wire \u2_Display/add122/c14 ;
  wire \u2_Display/add122/c15 ;
  wire \u2_Display/add122/c16 ;
  wire \u2_Display/add122/c17 ;
  wire \u2_Display/add122/c18 ;
  wire \u2_Display/add122/c19 ;
  wire \u2_Display/add122/c2 ;
  wire \u2_Display/add122/c20 ;
  wire \u2_Display/add122/c21 ;
  wire \u2_Display/add122/c22 ;
  wire \u2_Display/add122/c23 ;
  wire \u2_Display/add122/c24 ;
  wire \u2_Display/add122/c25 ;
  wire \u2_Display/add122/c26 ;
  wire \u2_Display/add122/c27 ;
  wire \u2_Display/add122/c28 ;
  wire \u2_Display/add122/c29 ;
  wire \u2_Display/add122/c3 ;
  wire \u2_Display/add122/c30 ;
  wire \u2_Display/add122/c31 ;
  wire \u2_Display/add122/c4 ;
  wire \u2_Display/add122/c5 ;
  wire \u2_Display/add122/c6 ;
  wire \u2_Display/add122/c7 ;
  wire \u2_Display/add122/c8 ;
  wire \u2_Display/add122/c9 ;
  wire \u2_Display/add123/c0 ;
  wire \u2_Display/add123/c1 ;
  wire \u2_Display/add123/c10 ;
  wire \u2_Display/add123/c11 ;
  wire \u2_Display/add123/c12 ;
  wire \u2_Display/add123/c13 ;
  wire \u2_Display/add123/c14 ;
  wire \u2_Display/add123/c15 ;
  wire \u2_Display/add123/c16 ;
  wire \u2_Display/add123/c17 ;
  wire \u2_Display/add123/c18 ;
  wire \u2_Display/add123/c19 ;
  wire \u2_Display/add123/c2 ;
  wire \u2_Display/add123/c20 ;
  wire \u2_Display/add123/c21 ;
  wire \u2_Display/add123/c22 ;
  wire \u2_Display/add123/c23 ;
  wire \u2_Display/add123/c24 ;
  wire \u2_Display/add123/c25 ;
  wire \u2_Display/add123/c26 ;
  wire \u2_Display/add123/c27 ;
  wire \u2_Display/add123/c28 ;
  wire \u2_Display/add123/c29 ;
  wire \u2_Display/add123/c3 ;
  wire \u2_Display/add123/c30 ;
  wire \u2_Display/add123/c31 ;
  wire \u2_Display/add123/c4 ;
  wire \u2_Display/add123/c5 ;
  wire \u2_Display/add123/c6 ;
  wire \u2_Display/add123/c7 ;
  wire \u2_Display/add123/c8 ;
  wire \u2_Display/add123/c9 ;
  wire \u2_Display/add124/c0 ;
  wire \u2_Display/add124/c1 ;
  wire \u2_Display/add124/c10 ;
  wire \u2_Display/add124/c11 ;
  wire \u2_Display/add124/c12 ;
  wire \u2_Display/add124/c13 ;
  wire \u2_Display/add124/c14 ;
  wire \u2_Display/add124/c15 ;
  wire \u2_Display/add124/c16 ;
  wire \u2_Display/add124/c17 ;
  wire \u2_Display/add124/c18 ;
  wire \u2_Display/add124/c19 ;
  wire \u2_Display/add124/c2 ;
  wire \u2_Display/add124/c20 ;
  wire \u2_Display/add124/c21 ;
  wire \u2_Display/add124/c22 ;
  wire \u2_Display/add124/c23 ;
  wire \u2_Display/add124/c24 ;
  wire \u2_Display/add124/c25 ;
  wire \u2_Display/add124/c26 ;
  wire \u2_Display/add124/c27 ;
  wire \u2_Display/add124/c28 ;
  wire \u2_Display/add124/c29 ;
  wire \u2_Display/add124/c3 ;
  wire \u2_Display/add124/c30 ;
  wire \u2_Display/add124/c31 ;
  wire \u2_Display/add124/c4 ;
  wire \u2_Display/add124/c5 ;
  wire \u2_Display/add124/c6 ;
  wire \u2_Display/add124/c7 ;
  wire \u2_Display/add124/c8 ;
  wire \u2_Display/add124/c9 ;
  wire \u2_Display/add125/c0 ;
  wire \u2_Display/add125/c1 ;
  wire \u2_Display/add125/c10 ;
  wire \u2_Display/add125/c11 ;
  wire \u2_Display/add125/c12 ;
  wire \u2_Display/add125/c13 ;
  wire \u2_Display/add125/c14 ;
  wire \u2_Display/add125/c15 ;
  wire \u2_Display/add125/c16 ;
  wire \u2_Display/add125/c17 ;
  wire \u2_Display/add125/c18 ;
  wire \u2_Display/add125/c19 ;
  wire \u2_Display/add125/c2 ;
  wire \u2_Display/add125/c20 ;
  wire \u2_Display/add125/c21 ;
  wire \u2_Display/add125/c22 ;
  wire \u2_Display/add125/c23 ;
  wire \u2_Display/add125/c24 ;
  wire \u2_Display/add125/c25 ;
  wire \u2_Display/add125/c26 ;
  wire \u2_Display/add125/c27 ;
  wire \u2_Display/add125/c28 ;
  wire \u2_Display/add125/c29 ;
  wire \u2_Display/add125/c3 ;
  wire \u2_Display/add125/c30 ;
  wire \u2_Display/add125/c31 ;
  wire \u2_Display/add125/c4 ;
  wire \u2_Display/add125/c5 ;
  wire \u2_Display/add125/c6 ;
  wire \u2_Display/add125/c7 ;
  wire \u2_Display/add125/c8 ;
  wire \u2_Display/add125/c9 ;
  wire \u2_Display/add126/c0 ;
  wire \u2_Display/add126/c1 ;
  wire \u2_Display/add126/c10 ;
  wire \u2_Display/add126/c11 ;
  wire \u2_Display/add126/c12 ;
  wire \u2_Display/add126/c13 ;
  wire \u2_Display/add126/c14 ;
  wire \u2_Display/add126/c15 ;
  wire \u2_Display/add126/c16 ;
  wire \u2_Display/add126/c17 ;
  wire \u2_Display/add126/c18 ;
  wire \u2_Display/add126/c19 ;
  wire \u2_Display/add126/c2 ;
  wire \u2_Display/add126/c20 ;
  wire \u2_Display/add126/c21 ;
  wire \u2_Display/add126/c22 ;
  wire \u2_Display/add126/c23 ;
  wire \u2_Display/add126/c24 ;
  wire \u2_Display/add126/c25 ;
  wire \u2_Display/add126/c26 ;
  wire \u2_Display/add126/c27 ;
  wire \u2_Display/add126/c28 ;
  wire \u2_Display/add126/c29 ;
  wire \u2_Display/add126/c3 ;
  wire \u2_Display/add126/c30 ;
  wire \u2_Display/add126/c31 ;
  wire \u2_Display/add126/c4 ;
  wire \u2_Display/add126/c5 ;
  wire \u2_Display/add126/c6 ;
  wire \u2_Display/add126/c7 ;
  wire \u2_Display/add126/c8 ;
  wire \u2_Display/add126/c9 ;
  wire \u2_Display/add127/c0 ;
  wire \u2_Display/add127/c1 ;
  wire \u2_Display/add127/c10 ;
  wire \u2_Display/add127/c11 ;
  wire \u2_Display/add127/c12 ;
  wire \u2_Display/add127/c13 ;
  wire \u2_Display/add127/c14 ;
  wire \u2_Display/add127/c15 ;
  wire \u2_Display/add127/c16 ;
  wire \u2_Display/add127/c17 ;
  wire \u2_Display/add127/c18 ;
  wire \u2_Display/add127/c19 ;
  wire \u2_Display/add127/c2 ;
  wire \u2_Display/add127/c20 ;
  wire \u2_Display/add127/c21 ;
  wire \u2_Display/add127/c22 ;
  wire \u2_Display/add127/c23 ;
  wire \u2_Display/add127/c24 ;
  wire \u2_Display/add127/c25 ;
  wire \u2_Display/add127/c26 ;
  wire \u2_Display/add127/c27 ;
  wire \u2_Display/add127/c28 ;
  wire \u2_Display/add127/c29 ;
  wire \u2_Display/add127/c3 ;
  wire \u2_Display/add127/c30 ;
  wire \u2_Display/add127/c31 ;
  wire \u2_Display/add127/c4 ;
  wire \u2_Display/add127/c5 ;
  wire \u2_Display/add127/c6 ;
  wire \u2_Display/add127/c7 ;
  wire \u2_Display/add127/c8 ;
  wire \u2_Display/add127/c9 ;
  wire \u2_Display/add128/c0 ;
  wire \u2_Display/add128/c1 ;
  wire \u2_Display/add128/c10 ;
  wire \u2_Display/add128/c11 ;
  wire \u2_Display/add128/c12 ;
  wire \u2_Display/add128/c13 ;
  wire \u2_Display/add128/c14 ;
  wire \u2_Display/add128/c15 ;
  wire \u2_Display/add128/c16 ;
  wire \u2_Display/add128/c17 ;
  wire \u2_Display/add128/c18 ;
  wire \u2_Display/add128/c19 ;
  wire \u2_Display/add128/c2 ;
  wire \u2_Display/add128/c20 ;
  wire \u2_Display/add128/c21 ;
  wire \u2_Display/add128/c22 ;
  wire \u2_Display/add128/c23 ;
  wire \u2_Display/add128/c24 ;
  wire \u2_Display/add128/c25 ;
  wire \u2_Display/add128/c26 ;
  wire \u2_Display/add128/c27 ;
  wire \u2_Display/add128/c28 ;
  wire \u2_Display/add128/c29 ;
  wire \u2_Display/add128/c3 ;
  wire \u2_Display/add128/c30 ;
  wire \u2_Display/add128/c31 ;
  wire \u2_Display/add128/c4 ;
  wire \u2_Display/add128/c5 ;
  wire \u2_Display/add128/c6 ;
  wire \u2_Display/add128/c7 ;
  wire \u2_Display/add128/c8 ;
  wire \u2_Display/add128/c9 ;
  wire \u2_Display/add129/c0 ;
  wire \u2_Display/add129/c1 ;
  wire \u2_Display/add129/c10 ;
  wire \u2_Display/add129/c11 ;
  wire \u2_Display/add129/c12 ;
  wire \u2_Display/add129/c13 ;
  wire \u2_Display/add129/c14 ;
  wire \u2_Display/add129/c15 ;
  wire \u2_Display/add129/c16 ;
  wire \u2_Display/add129/c17 ;
  wire \u2_Display/add129/c18 ;
  wire \u2_Display/add129/c19 ;
  wire \u2_Display/add129/c2 ;
  wire \u2_Display/add129/c20 ;
  wire \u2_Display/add129/c21 ;
  wire \u2_Display/add129/c22 ;
  wire \u2_Display/add129/c23 ;
  wire \u2_Display/add129/c24 ;
  wire \u2_Display/add129/c25 ;
  wire \u2_Display/add129/c26 ;
  wire \u2_Display/add129/c27 ;
  wire \u2_Display/add129/c28 ;
  wire \u2_Display/add129/c29 ;
  wire \u2_Display/add129/c3 ;
  wire \u2_Display/add129/c30 ;
  wire \u2_Display/add129/c31 ;
  wire \u2_Display/add129/c4 ;
  wire \u2_Display/add129/c5 ;
  wire \u2_Display/add129/c6 ;
  wire \u2_Display/add129/c7 ;
  wire \u2_Display/add129/c8 ;
  wire \u2_Display/add129/c9 ;
  wire \u2_Display/add130/c0 ;
  wire \u2_Display/add130/c1 ;
  wire \u2_Display/add130/c10 ;
  wire \u2_Display/add130/c11 ;
  wire \u2_Display/add130/c12 ;
  wire \u2_Display/add130/c13 ;
  wire \u2_Display/add130/c14 ;
  wire \u2_Display/add130/c15 ;
  wire \u2_Display/add130/c16 ;
  wire \u2_Display/add130/c17 ;
  wire \u2_Display/add130/c18 ;
  wire \u2_Display/add130/c19 ;
  wire \u2_Display/add130/c2 ;
  wire \u2_Display/add130/c20 ;
  wire \u2_Display/add130/c21 ;
  wire \u2_Display/add130/c22 ;
  wire \u2_Display/add130/c23 ;
  wire \u2_Display/add130/c24 ;
  wire \u2_Display/add130/c25 ;
  wire \u2_Display/add130/c26 ;
  wire \u2_Display/add130/c27 ;
  wire \u2_Display/add130/c28 ;
  wire \u2_Display/add130/c29 ;
  wire \u2_Display/add130/c3 ;
  wire \u2_Display/add130/c30 ;
  wire \u2_Display/add130/c31 ;
  wire \u2_Display/add130/c4 ;
  wire \u2_Display/add130/c5 ;
  wire \u2_Display/add130/c6 ;
  wire \u2_Display/add130/c7 ;
  wire \u2_Display/add130/c8 ;
  wire \u2_Display/add130/c9 ;
  wire \u2_Display/add131/c0 ;
  wire \u2_Display/add131/c1 ;
  wire \u2_Display/add131/c10 ;
  wire \u2_Display/add131/c11 ;
  wire \u2_Display/add131/c12 ;
  wire \u2_Display/add131/c13 ;
  wire \u2_Display/add131/c14 ;
  wire \u2_Display/add131/c15 ;
  wire \u2_Display/add131/c16 ;
  wire \u2_Display/add131/c17 ;
  wire \u2_Display/add131/c18 ;
  wire \u2_Display/add131/c19 ;
  wire \u2_Display/add131/c2 ;
  wire \u2_Display/add131/c20 ;
  wire \u2_Display/add131/c21 ;
  wire \u2_Display/add131/c22 ;
  wire \u2_Display/add131/c23 ;
  wire \u2_Display/add131/c24 ;
  wire \u2_Display/add131/c25 ;
  wire \u2_Display/add131/c26 ;
  wire \u2_Display/add131/c27 ;
  wire \u2_Display/add131/c28 ;
  wire \u2_Display/add131/c29 ;
  wire \u2_Display/add131/c3 ;
  wire \u2_Display/add131/c30 ;
  wire \u2_Display/add131/c31 ;
  wire \u2_Display/add131/c4 ;
  wire \u2_Display/add131/c5 ;
  wire \u2_Display/add131/c6 ;
  wire \u2_Display/add131/c7 ;
  wire \u2_Display/add131/c8 ;
  wire \u2_Display/add131/c9 ;
  wire \u2_Display/add132/c0 ;
  wire \u2_Display/add132/c1 ;
  wire \u2_Display/add132/c10 ;
  wire \u2_Display/add132/c11 ;
  wire \u2_Display/add132/c12 ;
  wire \u2_Display/add132/c13 ;
  wire \u2_Display/add132/c14 ;
  wire \u2_Display/add132/c15 ;
  wire \u2_Display/add132/c16 ;
  wire \u2_Display/add132/c17 ;
  wire \u2_Display/add132/c18 ;
  wire \u2_Display/add132/c19 ;
  wire \u2_Display/add132/c2 ;
  wire \u2_Display/add132/c20 ;
  wire \u2_Display/add132/c21 ;
  wire \u2_Display/add132/c22 ;
  wire \u2_Display/add132/c23 ;
  wire \u2_Display/add132/c24 ;
  wire \u2_Display/add132/c25 ;
  wire \u2_Display/add132/c26 ;
  wire \u2_Display/add132/c27 ;
  wire \u2_Display/add132/c28 ;
  wire \u2_Display/add132/c29 ;
  wire \u2_Display/add132/c3 ;
  wire \u2_Display/add132/c30 ;
  wire \u2_Display/add132/c31 ;
  wire \u2_Display/add132/c4 ;
  wire \u2_Display/add132/c5 ;
  wire \u2_Display/add132/c6 ;
  wire \u2_Display/add132/c7 ;
  wire \u2_Display/add132/c8 ;
  wire \u2_Display/add132/c9 ;
  wire \u2_Display/add133/c0 ;
  wire \u2_Display/add133/c1 ;
  wire \u2_Display/add133/c10 ;
  wire \u2_Display/add133/c11 ;
  wire \u2_Display/add133/c12 ;
  wire \u2_Display/add133/c13 ;
  wire \u2_Display/add133/c14 ;
  wire \u2_Display/add133/c15 ;
  wire \u2_Display/add133/c16 ;
  wire \u2_Display/add133/c17 ;
  wire \u2_Display/add133/c18 ;
  wire \u2_Display/add133/c19 ;
  wire \u2_Display/add133/c2 ;
  wire \u2_Display/add133/c20 ;
  wire \u2_Display/add133/c21 ;
  wire \u2_Display/add133/c22 ;
  wire \u2_Display/add133/c23 ;
  wire \u2_Display/add133/c24 ;
  wire \u2_Display/add133/c25 ;
  wire \u2_Display/add133/c26 ;
  wire \u2_Display/add133/c27 ;
  wire \u2_Display/add133/c28 ;
  wire \u2_Display/add133/c29 ;
  wire \u2_Display/add133/c3 ;
  wire \u2_Display/add133/c30 ;
  wire \u2_Display/add133/c31 ;
  wire \u2_Display/add133/c4 ;
  wire \u2_Display/add133/c5 ;
  wire \u2_Display/add133/c6 ;
  wire \u2_Display/add133/c7 ;
  wire \u2_Display/add133/c8 ;
  wire \u2_Display/add133/c9 ;
  wire \u2_Display/add134/c0 ;
  wire \u2_Display/add134/c1 ;
  wire \u2_Display/add134/c10 ;
  wire \u2_Display/add134/c11 ;
  wire \u2_Display/add134/c12 ;
  wire \u2_Display/add134/c13 ;
  wire \u2_Display/add134/c14 ;
  wire \u2_Display/add134/c15 ;
  wire \u2_Display/add134/c16 ;
  wire \u2_Display/add134/c17 ;
  wire \u2_Display/add134/c18 ;
  wire \u2_Display/add134/c19 ;
  wire \u2_Display/add134/c2 ;
  wire \u2_Display/add134/c20 ;
  wire \u2_Display/add134/c21 ;
  wire \u2_Display/add134/c22 ;
  wire \u2_Display/add134/c23 ;
  wire \u2_Display/add134/c24 ;
  wire \u2_Display/add134/c25 ;
  wire \u2_Display/add134/c26 ;
  wire \u2_Display/add134/c27 ;
  wire \u2_Display/add134/c28 ;
  wire \u2_Display/add134/c29 ;
  wire \u2_Display/add134/c3 ;
  wire \u2_Display/add134/c30 ;
  wire \u2_Display/add134/c31 ;
  wire \u2_Display/add134/c4 ;
  wire \u2_Display/add134/c5 ;
  wire \u2_Display/add134/c6 ;
  wire \u2_Display/add134/c7 ;
  wire \u2_Display/add134/c8 ;
  wire \u2_Display/add134/c9 ;
  wire \u2_Display/add135/c0 ;
  wire \u2_Display/add135/c1 ;
  wire \u2_Display/add135/c10 ;
  wire \u2_Display/add135/c11 ;
  wire \u2_Display/add135/c12 ;
  wire \u2_Display/add135/c13 ;
  wire \u2_Display/add135/c14 ;
  wire \u2_Display/add135/c15 ;
  wire \u2_Display/add135/c16 ;
  wire \u2_Display/add135/c17 ;
  wire \u2_Display/add135/c18 ;
  wire \u2_Display/add135/c19 ;
  wire \u2_Display/add135/c2 ;
  wire \u2_Display/add135/c20 ;
  wire \u2_Display/add135/c21 ;
  wire \u2_Display/add135/c22 ;
  wire \u2_Display/add135/c23 ;
  wire \u2_Display/add135/c24 ;
  wire \u2_Display/add135/c25 ;
  wire \u2_Display/add135/c26 ;
  wire \u2_Display/add135/c27 ;
  wire \u2_Display/add135/c28 ;
  wire \u2_Display/add135/c29 ;
  wire \u2_Display/add135/c3 ;
  wire \u2_Display/add135/c30 ;
  wire \u2_Display/add135/c31 ;
  wire \u2_Display/add135/c4 ;
  wire \u2_Display/add135/c5 ;
  wire \u2_Display/add135/c6 ;
  wire \u2_Display/add135/c7 ;
  wire \u2_Display/add135/c8 ;
  wire \u2_Display/add135/c9 ;
  wire \u2_Display/add136/c0 ;
  wire \u2_Display/add136/c1 ;
  wire \u2_Display/add136/c10 ;
  wire \u2_Display/add136/c11 ;
  wire \u2_Display/add136/c12 ;
  wire \u2_Display/add136/c13 ;
  wire \u2_Display/add136/c14 ;
  wire \u2_Display/add136/c15 ;
  wire \u2_Display/add136/c16 ;
  wire \u2_Display/add136/c17 ;
  wire \u2_Display/add136/c18 ;
  wire \u2_Display/add136/c19 ;
  wire \u2_Display/add136/c2 ;
  wire \u2_Display/add136/c20 ;
  wire \u2_Display/add136/c21 ;
  wire \u2_Display/add136/c22 ;
  wire \u2_Display/add136/c23 ;
  wire \u2_Display/add136/c24 ;
  wire \u2_Display/add136/c25 ;
  wire \u2_Display/add136/c26 ;
  wire \u2_Display/add136/c27 ;
  wire \u2_Display/add136/c28 ;
  wire \u2_Display/add136/c29 ;
  wire \u2_Display/add136/c3 ;
  wire \u2_Display/add136/c30 ;
  wire \u2_Display/add136/c31 ;
  wire \u2_Display/add136/c4 ;
  wire \u2_Display/add136/c5 ;
  wire \u2_Display/add136/c6 ;
  wire \u2_Display/add136/c7 ;
  wire \u2_Display/add136/c8 ;
  wire \u2_Display/add136/c9 ;
  wire \u2_Display/add137/c0 ;
  wire \u2_Display/add137/c1 ;
  wire \u2_Display/add137/c10 ;
  wire \u2_Display/add137/c11 ;
  wire \u2_Display/add137/c12 ;
  wire \u2_Display/add137/c13 ;
  wire \u2_Display/add137/c14 ;
  wire \u2_Display/add137/c15 ;
  wire \u2_Display/add137/c16 ;
  wire \u2_Display/add137/c17 ;
  wire \u2_Display/add137/c18 ;
  wire \u2_Display/add137/c19 ;
  wire \u2_Display/add137/c2 ;
  wire \u2_Display/add137/c20 ;
  wire \u2_Display/add137/c21 ;
  wire \u2_Display/add137/c22 ;
  wire \u2_Display/add137/c23 ;
  wire \u2_Display/add137/c24 ;
  wire \u2_Display/add137/c25 ;
  wire \u2_Display/add137/c26 ;
  wire \u2_Display/add137/c27 ;
  wire \u2_Display/add137/c28 ;
  wire \u2_Display/add137/c29 ;
  wire \u2_Display/add137/c3 ;
  wire \u2_Display/add137/c30 ;
  wire \u2_Display/add137/c31 ;
  wire \u2_Display/add137/c4 ;
  wire \u2_Display/add137/c5 ;
  wire \u2_Display/add137/c6 ;
  wire \u2_Display/add137/c7 ;
  wire \u2_Display/add137/c8 ;
  wire \u2_Display/add137/c9 ;
  wire \u2_Display/add138/c0 ;
  wire \u2_Display/add138/c1 ;
  wire \u2_Display/add138/c10 ;
  wire \u2_Display/add138/c11 ;
  wire \u2_Display/add138/c12 ;
  wire \u2_Display/add138/c13 ;
  wire \u2_Display/add138/c14 ;
  wire \u2_Display/add138/c15 ;
  wire \u2_Display/add138/c16 ;
  wire \u2_Display/add138/c17 ;
  wire \u2_Display/add138/c18 ;
  wire \u2_Display/add138/c19 ;
  wire \u2_Display/add138/c2 ;
  wire \u2_Display/add138/c20 ;
  wire \u2_Display/add138/c21 ;
  wire \u2_Display/add138/c22 ;
  wire \u2_Display/add138/c23 ;
  wire \u2_Display/add138/c24 ;
  wire \u2_Display/add138/c25 ;
  wire \u2_Display/add138/c26 ;
  wire \u2_Display/add138/c27 ;
  wire \u2_Display/add138/c28 ;
  wire \u2_Display/add138/c29 ;
  wire \u2_Display/add138/c3 ;
  wire \u2_Display/add138/c30 ;
  wire \u2_Display/add138/c31 ;
  wire \u2_Display/add138/c4 ;
  wire \u2_Display/add138/c5 ;
  wire \u2_Display/add138/c6 ;
  wire \u2_Display/add138/c7 ;
  wire \u2_Display/add138/c8 ;
  wire \u2_Display/add138/c9 ;
  wire \u2_Display/add139/c0 ;
  wire \u2_Display/add139/c1 ;
  wire \u2_Display/add139/c2 ;
  wire \u2_Display/add139/c3 ;
  wire \u2_Display/add139/c4 ;
  wire \u2_Display/add139/c5 ;
  wire \u2_Display/add139/c6 ;
  wire \u2_Display/add139/c7 ;
  wire \u2_Display/add139/c8 ;
  wire \u2_Display/add139/c9 ;
  wire \u2_Display/add14/c0 ;
  wire \u2_Display/add14/c1 ;
  wire \u2_Display/add14/c10 ;
  wire \u2_Display/add14/c11 ;
  wire \u2_Display/add14/c12 ;
  wire \u2_Display/add14/c13 ;
  wire \u2_Display/add14/c14 ;
  wire \u2_Display/add14/c15 ;
  wire \u2_Display/add14/c16 ;
  wire \u2_Display/add14/c17 ;
  wire \u2_Display/add14/c18 ;
  wire \u2_Display/add14/c19 ;
  wire \u2_Display/add14/c2 ;
  wire \u2_Display/add14/c20 ;
  wire \u2_Display/add14/c21 ;
  wire \u2_Display/add14/c22 ;
  wire \u2_Display/add14/c23 ;
  wire \u2_Display/add14/c24 ;
  wire \u2_Display/add14/c25 ;
  wire \u2_Display/add14/c26 ;
  wire \u2_Display/add14/c27 ;
  wire \u2_Display/add14/c28 ;
  wire \u2_Display/add14/c29 ;
  wire \u2_Display/add14/c3 ;
  wire \u2_Display/add14/c30 ;
  wire \u2_Display/add14/c31 ;
  wire \u2_Display/add14/c4 ;
  wire \u2_Display/add14/c5 ;
  wire \u2_Display/add14/c6 ;
  wire \u2_Display/add14/c7 ;
  wire \u2_Display/add14/c8 ;
  wire \u2_Display/add14/c9 ;
  wire \u2_Display/add151/c0 ;
  wire \u2_Display/add151/c1 ;
  wire \u2_Display/add151/c10 ;
  wire \u2_Display/add151/c11 ;
  wire \u2_Display/add151/c12 ;
  wire \u2_Display/add151/c13 ;
  wire \u2_Display/add151/c14 ;
  wire \u2_Display/add151/c15 ;
  wire \u2_Display/add151/c16 ;
  wire \u2_Display/add151/c17 ;
  wire \u2_Display/add151/c18 ;
  wire \u2_Display/add151/c19 ;
  wire \u2_Display/add151/c2 ;
  wire \u2_Display/add151/c20 ;
  wire \u2_Display/add151/c21 ;
  wire \u2_Display/add151/c22 ;
  wire \u2_Display/add151/c23 ;
  wire \u2_Display/add151/c24 ;
  wire \u2_Display/add151/c25 ;
  wire \u2_Display/add151/c26 ;
  wire \u2_Display/add151/c27 ;
  wire \u2_Display/add151/c28 ;
  wire \u2_Display/add151/c29 ;
  wire \u2_Display/add151/c3 ;
  wire \u2_Display/add151/c30 ;
  wire \u2_Display/add151/c31 ;
  wire \u2_Display/add151/c4 ;
  wire \u2_Display/add151/c5 ;
  wire \u2_Display/add151/c6 ;
  wire \u2_Display/add151/c7 ;
  wire \u2_Display/add151/c8 ;
  wire \u2_Display/add151/c9 ;
  wire \u2_Display/add152/c0 ;
  wire \u2_Display/add152/c1 ;
  wire \u2_Display/add152/c10 ;
  wire \u2_Display/add152/c11 ;
  wire \u2_Display/add152/c12 ;
  wire \u2_Display/add152/c13 ;
  wire \u2_Display/add152/c14 ;
  wire \u2_Display/add152/c15 ;
  wire \u2_Display/add152/c16 ;
  wire \u2_Display/add152/c17 ;
  wire \u2_Display/add152/c18 ;
  wire \u2_Display/add152/c19 ;
  wire \u2_Display/add152/c2 ;
  wire \u2_Display/add152/c20 ;
  wire \u2_Display/add152/c21 ;
  wire \u2_Display/add152/c22 ;
  wire \u2_Display/add152/c23 ;
  wire \u2_Display/add152/c24 ;
  wire \u2_Display/add152/c25 ;
  wire \u2_Display/add152/c26 ;
  wire \u2_Display/add152/c27 ;
  wire \u2_Display/add152/c28 ;
  wire \u2_Display/add152/c29 ;
  wire \u2_Display/add152/c3 ;
  wire \u2_Display/add152/c30 ;
  wire \u2_Display/add152/c31 ;
  wire \u2_Display/add152/c4 ;
  wire \u2_Display/add152/c5 ;
  wire \u2_Display/add152/c6 ;
  wire \u2_Display/add152/c7 ;
  wire \u2_Display/add152/c8 ;
  wire \u2_Display/add152/c9 ;
  wire \u2_Display/add153/c0 ;
  wire \u2_Display/add153/c1 ;
  wire \u2_Display/add153/c10 ;
  wire \u2_Display/add153/c11 ;
  wire \u2_Display/add153/c12 ;
  wire \u2_Display/add153/c13 ;
  wire \u2_Display/add153/c14 ;
  wire \u2_Display/add153/c15 ;
  wire \u2_Display/add153/c16 ;
  wire \u2_Display/add153/c17 ;
  wire \u2_Display/add153/c18 ;
  wire \u2_Display/add153/c19 ;
  wire \u2_Display/add153/c2 ;
  wire \u2_Display/add153/c20 ;
  wire \u2_Display/add153/c21 ;
  wire \u2_Display/add153/c22 ;
  wire \u2_Display/add153/c23 ;
  wire \u2_Display/add153/c24 ;
  wire \u2_Display/add153/c25 ;
  wire \u2_Display/add153/c26 ;
  wire \u2_Display/add153/c27 ;
  wire \u2_Display/add153/c28 ;
  wire \u2_Display/add153/c29 ;
  wire \u2_Display/add153/c3 ;
  wire \u2_Display/add153/c30 ;
  wire \u2_Display/add153/c31 ;
  wire \u2_Display/add153/c4 ;
  wire \u2_Display/add153/c5 ;
  wire \u2_Display/add153/c6 ;
  wire \u2_Display/add153/c7 ;
  wire \u2_Display/add153/c8 ;
  wire \u2_Display/add153/c9 ;
  wire \u2_Display/add154/c0 ;
  wire \u2_Display/add154/c1 ;
  wire \u2_Display/add154/c10 ;
  wire \u2_Display/add154/c11 ;
  wire \u2_Display/add154/c12 ;
  wire \u2_Display/add154/c13 ;
  wire \u2_Display/add154/c14 ;
  wire \u2_Display/add154/c15 ;
  wire \u2_Display/add154/c16 ;
  wire \u2_Display/add154/c17 ;
  wire \u2_Display/add154/c18 ;
  wire \u2_Display/add154/c19 ;
  wire \u2_Display/add154/c2 ;
  wire \u2_Display/add154/c20 ;
  wire \u2_Display/add154/c21 ;
  wire \u2_Display/add154/c22 ;
  wire \u2_Display/add154/c23 ;
  wire \u2_Display/add154/c24 ;
  wire \u2_Display/add154/c25 ;
  wire \u2_Display/add154/c26 ;
  wire \u2_Display/add154/c27 ;
  wire \u2_Display/add154/c28 ;
  wire \u2_Display/add154/c29 ;
  wire \u2_Display/add154/c3 ;
  wire \u2_Display/add154/c30 ;
  wire \u2_Display/add154/c31 ;
  wire \u2_Display/add154/c4 ;
  wire \u2_Display/add154/c5 ;
  wire \u2_Display/add154/c6 ;
  wire \u2_Display/add154/c7 ;
  wire \u2_Display/add154/c8 ;
  wire \u2_Display/add154/c9 ;
  wire \u2_Display/add155/c0 ;
  wire \u2_Display/add155/c1 ;
  wire \u2_Display/add155/c10 ;
  wire \u2_Display/add155/c11 ;
  wire \u2_Display/add155/c12 ;
  wire \u2_Display/add155/c13 ;
  wire \u2_Display/add155/c14 ;
  wire \u2_Display/add155/c15 ;
  wire \u2_Display/add155/c16 ;
  wire \u2_Display/add155/c17 ;
  wire \u2_Display/add155/c18 ;
  wire \u2_Display/add155/c19 ;
  wire \u2_Display/add155/c2 ;
  wire \u2_Display/add155/c20 ;
  wire \u2_Display/add155/c21 ;
  wire \u2_Display/add155/c22 ;
  wire \u2_Display/add155/c23 ;
  wire \u2_Display/add155/c24 ;
  wire \u2_Display/add155/c25 ;
  wire \u2_Display/add155/c26 ;
  wire \u2_Display/add155/c27 ;
  wire \u2_Display/add155/c28 ;
  wire \u2_Display/add155/c29 ;
  wire \u2_Display/add155/c3 ;
  wire \u2_Display/add155/c30 ;
  wire \u2_Display/add155/c31 ;
  wire \u2_Display/add155/c4 ;
  wire \u2_Display/add155/c5 ;
  wire \u2_Display/add155/c6 ;
  wire \u2_Display/add155/c7 ;
  wire \u2_Display/add155/c8 ;
  wire \u2_Display/add155/c9 ;
  wire \u2_Display/add156/c0 ;
  wire \u2_Display/add156/c1 ;
  wire \u2_Display/add156/c10 ;
  wire \u2_Display/add156/c11 ;
  wire \u2_Display/add156/c12 ;
  wire \u2_Display/add156/c13 ;
  wire \u2_Display/add156/c14 ;
  wire \u2_Display/add156/c15 ;
  wire \u2_Display/add156/c16 ;
  wire \u2_Display/add156/c17 ;
  wire \u2_Display/add156/c18 ;
  wire \u2_Display/add156/c19 ;
  wire \u2_Display/add156/c2 ;
  wire \u2_Display/add156/c20 ;
  wire \u2_Display/add156/c21 ;
  wire \u2_Display/add156/c22 ;
  wire \u2_Display/add156/c23 ;
  wire \u2_Display/add156/c24 ;
  wire \u2_Display/add156/c25 ;
  wire \u2_Display/add156/c26 ;
  wire \u2_Display/add156/c27 ;
  wire \u2_Display/add156/c28 ;
  wire \u2_Display/add156/c29 ;
  wire \u2_Display/add156/c3 ;
  wire \u2_Display/add156/c30 ;
  wire \u2_Display/add156/c31 ;
  wire \u2_Display/add156/c4 ;
  wire \u2_Display/add156/c5 ;
  wire \u2_Display/add156/c6 ;
  wire \u2_Display/add156/c7 ;
  wire \u2_Display/add156/c8 ;
  wire \u2_Display/add156/c9 ;
  wire \u2_Display/add157/c0 ;
  wire \u2_Display/add157/c1 ;
  wire \u2_Display/add157/c10 ;
  wire \u2_Display/add157/c11 ;
  wire \u2_Display/add157/c12 ;
  wire \u2_Display/add157/c13 ;
  wire \u2_Display/add157/c14 ;
  wire \u2_Display/add157/c15 ;
  wire \u2_Display/add157/c16 ;
  wire \u2_Display/add157/c17 ;
  wire \u2_Display/add157/c18 ;
  wire \u2_Display/add157/c19 ;
  wire \u2_Display/add157/c2 ;
  wire \u2_Display/add157/c20 ;
  wire \u2_Display/add157/c21 ;
  wire \u2_Display/add157/c22 ;
  wire \u2_Display/add157/c23 ;
  wire \u2_Display/add157/c24 ;
  wire \u2_Display/add157/c25 ;
  wire \u2_Display/add157/c26 ;
  wire \u2_Display/add157/c27 ;
  wire \u2_Display/add157/c28 ;
  wire \u2_Display/add157/c29 ;
  wire \u2_Display/add157/c3 ;
  wire \u2_Display/add157/c30 ;
  wire \u2_Display/add157/c31 ;
  wire \u2_Display/add157/c4 ;
  wire \u2_Display/add157/c5 ;
  wire \u2_Display/add157/c6 ;
  wire \u2_Display/add157/c7 ;
  wire \u2_Display/add157/c8 ;
  wire \u2_Display/add157/c9 ;
  wire \u2_Display/add158/c0 ;
  wire \u2_Display/add158/c1 ;
  wire \u2_Display/add158/c10 ;
  wire \u2_Display/add158/c11 ;
  wire \u2_Display/add158/c12 ;
  wire \u2_Display/add158/c13 ;
  wire \u2_Display/add158/c14 ;
  wire \u2_Display/add158/c15 ;
  wire \u2_Display/add158/c16 ;
  wire \u2_Display/add158/c17 ;
  wire \u2_Display/add158/c18 ;
  wire \u2_Display/add158/c19 ;
  wire \u2_Display/add158/c2 ;
  wire \u2_Display/add158/c20 ;
  wire \u2_Display/add158/c21 ;
  wire \u2_Display/add158/c22 ;
  wire \u2_Display/add158/c23 ;
  wire \u2_Display/add158/c24 ;
  wire \u2_Display/add158/c25 ;
  wire \u2_Display/add158/c26 ;
  wire \u2_Display/add158/c27 ;
  wire \u2_Display/add158/c28 ;
  wire \u2_Display/add158/c29 ;
  wire \u2_Display/add158/c3 ;
  wire \u2_Display/add158/c30 ;
  wire \u2_Display/add158/c31 ;
  wire \u2_Display/add158/c4 ;
  wire \u2_Display/add158/c5 ;
  wire \u2_Display/add158/c6 ;
  wire \u2_Display/add158/c7 ;
  wire \u2_Display/add158/c8 ;
  wire \u2_Display/add158/c9 ;
  wire \u2_Display/add159/c0 ;
  wire \u2_Display/add159/c1 ;
  wire \u2_Display/add159/c10 ;
  wire \u2_Display/add159/c11 ;
  wire \u2_Display/add159/c12 ;
  wire \u2_Display/add159/c13 ;
  wire \u2_Display/add159/c14 ;
  wire \u2_Display/add159/c15 ;
  wire \u2_Display/add159/c16 ;
  wire \u2_Display/add159/c17 ;
  wire \u2_Display/add159/c18 ;
  wire \u2_Display/add159/c19 ;
  wire \u2_Display/add159/c2 ;
  wire \u2_Display/add159/c20 ;
  wire \u2_Display/add159/c21 ;
  wire \u2_Display/add159/c22 ;
  wire \u2_Display/add159/c23 ;
  wire \u2_Display/add159/c24 ;
  wire \u2_Display/add159/c25 ;
  wire \u2_Display/add159/c26 ;
  wire \u2_Display/add159/c27 ;
  wire \u2_Display/add159/c28 ;
  wire \u2_Display/add159/c29 ;
  wire \u2_Display/add159/c3 ;
  wire \u2_Display/add159/c30 ;
  wire \u2_Display/add159/c31 ;
  wire \u2_Display/add159/c4 ;
  wire \u2_Display/add159/c5 ;
  wire \u2_Display/add159/c6 ;
  wire \u2_Display/add159/c7 ;
  wire \u2_Display/add159/c8 ;
  wire \u2_Display/add159/c9 ;
  wire \u2_Display/add160/c0 ;
  wire \u2_Display/add160/c1 ;
  wire \u2_Display/add160/c10 ;
  wire \u2_Display/add160/c11 ;
  wire \u2_Display/add160/c12 ;
  wire \u2_Display/add160/c13 ;
  wire \u2_Display/add160/c14 ;
  wire \u2_Display/add160/c15 ;
  wire \u2_Display/add160/c16 ;
  wire \u2_Display/add160/c17 ;
  wire \u2_Display/add160/c18 ;
  wire \u2_Display/add160/c19 ;
  wire \u2_Display/add160/c2 ;
  wire \u2_Display/add160/c20 ;
  wire \u2_Display/add160/c21 ;
  wire \u2_Display/add160/c22 ;
  wire \u2_Display/add160/c23 ;
  wire \u2_Display/add160/c24 ;
  wire \u2_Display/add160/c25 ;
  wire \u2_Display/add160/c26 ;
  wire \u2_Display/add160/c27 ;
  wire \u2_Display/add160/c28 ;
  wire \u2_Display/add160/c29 ;
  wire \u2_Display/add160/c3 ;
  wire \u2_Display/add160/c30 ;
  wire \u2_Display/add160/c31 ;
  wire \u2_Display/add160/c4 ;
  wire \u2_Display/add160/c5 ;
  wire \u2_Display/add160/c6 ;
  wire \u2_Display/add160/c7 ;
  wire \u2_Display/add160/c8 ;
  wire \u2_Display/add160/c9 ;
  wire \u2_Display/add161/c0 ;
  wire \u2_Display/add161/c1 ;
  wire \u2_Display/add161/c10 ;
  wire \u2_Display/add161/c11 ;
  wire \u2_Display/add161/c12 ;
  wire \u2_Display/add161/c13 ;
  wire \u2_Display/add161/c14 ;
  wire \u2_Display/add161/c15 ;
  wire \u2_Display/add161/c16 ;
  wire \u2_Display/add161/c17 ;
  wire \u2_Display/add161/c18 ;
  wire \u2_Display/add161/c19 ;
  wire \u2_Display/add161/c2 ;
  wire \u2_Display/add161/c20 ;
  wire \u2_Display/add161/c21 ;
  wire \u2_Display/add161/c22 ;
  wire \u2_Display/add161/c23 ;
  wire \u2_Display/add161/c24 ;
  wire \u2_Display/add161/c25 ;
  wire \u2_Display/add161/c26 ;
  wire \u2_Display/add161/c27 ;
  wire \u2_Display/add161/c28 ;
  wire \u2_Display/add161/c29 ;
  wire \u2_Display/add161/c3 ;
  wire \u2_Display/add161/c30 ;
  wire \u2_Display/add161/c31 ;
  wire \u2_Display/add161/c4 ;
  wire \u2_Display/add161/c5 ;
  wire \u2_Display/add161/c6 ;
  wire \u2_Display/add161/c7 ;
  wire \u2_Display/add161/c8 ;
  wire \u2_Display/add161/c9 ;
  wire \u2_Display/add162/c0 ;
  wire \u2_Display/add162/c1 ;
  wire \u2_Display/add162/c10 ;
  wire \u2_Display/add162/c11 ;
  wire \u2_Display/add162/c12 ;
  wire \u2_Display/add162/c13 ;
  wire \u2_Display/add162/c14 ;
  wire \u2_Display/add162/c15 ;
  wire \u2_Display/add162/c16 ;
  wire \u2_Display/add162/c17 ;
  wire \u2_Display/add162/c18 ;
  wire \u2_Display/add162/c19 ;
  wire \u2_Display/add162/c2 ;
  wire \u2_Display/add162/c20 ;
  wire \u2_Display/add162/c21 ;
  wire \u2_Display/add162/c22 ;
  wire \u2_Display/add162/c23 ;
  wire \u2_Display/add162/c24 ;
  wire \u2_Display/add162/c25 ;
  wire \u2_Display/add162/c26 ;
  wire \u2_Display/add162/c27 ;
  wire \u2_Display/add162/c28 ;
  wire \u2_Display/add162/c29 ;
  wire \u2_Display/add162/c3 ;
  wire \u2_Display/add162/c30 ;
  wire \u2_Display/add162/c31 ;
  wire \u2_Display/add162/c4 ;
  wire \u2_Display/add162/c5 ;
  wire \u2_Display/add162/c6 ;
  wire \u2_Display/add162/c7 ;
  wire \u2_Display/add162/c8 ;
  wire \u2_Display/add162/c9 ;
  wire \u2_Display/add163/c0 ;
  wire \u2_Display/add163/c1 ;
  wire \u2_Display/add163/c10 ;
  wire \u2_Display/add163/c11 ;
  wire \u2_Display/add163/c12 ;
  wire \u2_Display/add163/c13 ;
  wire \u2_Display/add163/c14 ;
  wire \u2_Display/add163/c15 ;
  wire \u2_Display/add163/c16 ;
  wire \u2_Display/add163/c17 ;
  wire \u2_Display/add163/c18 ;
  wire \u2_Display/add163/c19 ;
  wire \u2_Display/add163/c2 ;
  wire \u2_Display/add163/c20 ;
  wire \u2_Display/add163/c21 ;
  wire \u2_Display/add163/c22 ;
  wire \u2_Display/add163/c23 ;
  wire \u2_Display/add163/c24 ;
  wire \u2_Display/add163/c25 ;
  wire \u2_Display/add163/c26 ;
  wire \u2_Display/add163/c27 ;
  wire \u2_Display/add163/c28 ;
  wire \u2_Display/add163/c29 ;
  wire \u2_Display/add163/c3 ;
  wire \u2_Display/add163/c30 ;
  wire \u2_Display/add163/c31 ;
  wire \u2_Display/add163/c4 ;
  wire \u2_Display/add163/c5 ;
  wire \u2_Display/add163/c6 ;
  wire \u2_Display/add163/c7 ;
  wire \u2_Display/add163/c8 ;
  wire \u2_Display/add163/c9 ;
  wire \u2_Display/add164/c0 ;
  wire \u2_Display/add164/c1 ;
  wire \u2_Display/add164/c10 ;
  wire \u2_Display/add164/c11 ;
  wire \u2_Display/add164/c12 ;
  wire \u2_Display/add164/c13 ;
  wire \u2_Display/add164/c14 ;
  wire \u2_Display/add164/c15 ;
  wire \u2_Display/add164/c16 ;
  wire \u2_Display/add164/c17 ;
  wire \u2_Display/add164/c18 ;
  wire \u2_Display/add164/c19 ;
  wire \u2_Display/add164/c2 ;
  wire \u2_Display/add164/c20 ;
  wire \u2_Display/add164/c21 ;
  wire \u2_Display/add164/c22 ;
  wire \u2_Display/add164/c23 ;
  wire \u2_Display/add164/c24 ;
  wire \u2_Display/add164/c25 ;
  wire \u2_Display/add164/c26 ;
  wire \u2_Display/add164/c27 ;
  wire \u2_Display/add164/c28 ;
  wire \u2_Display/add164/c29 ;
  wire \u2_Display/add164/c3 ;
  wire \u2_Display/add164/c30 ;
  wire \u2_Display/add164/c31 ;
  wire \u2_Display/add164/c4 ;
  wire \u2_Display/add164/c5 ;
  wire \u2_Display/add164/c6 ;
  wire \u2_Display/add164/c7 ;
  wire \u2_Display/add164/c8 ;
  wire \u2_Display/add164/c9 ;
  wire \u2_Display/add165/c0 ;
  wire \u2_Display/add165/c1 ;
  wire \u2_Display/add165/c10 ;
  wire \u2_Display/add165/c11 ;
  wire \u2_Display/add165/c12 ;
  wire \u2_Display/add165/c13 ;
  wire \u2_Display/add165/c14 ;
  wire \u2_Display/add165/c15 ;
  wire \u2_Display/add165/c16 ;
  wire \u2_Display/add165/c17 ;
  wire \u2_Display/add165/c18 ;
  wire \u2_Display/add165/c19 ;
  wire \u2_Display/add165/c2 ;
  wire \u2_Display/add165/c20 ;
  wire \u2_Display/add165/c21 ;
  wire \u2_Display/add165/c22 ;
  wire \u2_Display/add165/c23 ;
  wire \u2_Display/add165/c24 ;
  wire \u2_Display/add165/c25 ;
  wire \u2_Display/add165/c26 ;
  wire \u2_Display/add165/c27 ;
  wire \u2_Display/add165/c28 ;
  wire \u2_Display/add165/c29 ;
  wire \u2_Display/add165/c3 ;
  wire \u2_Display/add165/c30 ;
  wire \u2_Display/add165/c31 ;
  wire \u2_Display/add165/c4 ;
  wire \u2_Display/add165/c5 ;
  wire \u2_Display/add165/c6 ;
  wire \u2_Display/add165/c7 ;
  wire \u2_Display/add165/c8 ;
  wire \u2_Display/add165/c9 ;
  wire \u2_Display/add166/c0 ;
  wire \u2_Display/add166/c1 ;
  wire \u2_Display/add166/c10 ;
  wire \u2_Display/add166/c11 ;
  wire \u2_Display/add166/c12 ;
  wire \u2_Display/add166/c13 ;
  wire \u2_Display/add166/c14 ;
  wire \u2_Display/add166/c15 ;
  wire \u2_Display/add166/c16 ;
  wire \u2_Display/add166/c17 ;
  wire \u2_Display/add166/c18 ;
  wire \u2_Display/add166/c19 ;
  wire \u2_Display/add166/c2 ;
  wire \u2_Display/add166/c20 ;
  wire \u2_Display/add166/c21 ;
  wire \u2_Display/add166/c22 ;
  wire \u2_Display/add166/c23 ;
  wire \u2_Display/add166/c24 ;
  wire \u2_Display/add166/c25 ;
  wire \u2_Display/add166/c26 ;
  wire \u2_Display/add166/c27 ;
  wire \u2_Display/add166/c28 ;
  wire \u2_Display/add166/c29 ;
  wire \u2_Display/add166/c3 ;
  wire \u2_Display/add166/c30 ;
  wire \u2_Display/add166/c31 ;
  wire \u2_Display/add166/c4 ;
  wire \u2_Display/add166/c5 ;
  wire \u2_Display/add166/c6 ;
  wire \u2_Display/add166/c7 ;
  wire \u2_Display/add166/c8 ;
  wire \u2_Display/add166/c9 ;
  wire \u2_Display/add167/c0 ;
  wire \u2_Display/add167/c1 ;
  wire \u2_Display/add167/c10 ;
  wire \u2_Display/add167/c11 ;
  wire \u2_Display/add167/c12 ;
  wire \u2_Display/add167/c13 ;
  wire \u2_Display/add167/c14 ;
  wire \u2_Display/add167/c15 ;
  wire \u2_Display/add167/c16 ;
  wire \u2_Display/add167/c17 ;
  wire \u2_Display/add167/c18 ;
  wire \u2_Display/add167/c19 ;
  wire \u2_Display/add167/c2 ;
  wire \u2_Display/add167/c20 ;
  wire \u2_Display/add167/c21 ;
  wire \u2_Display/add167/c22 ;
  wire \u2_Display/add167/c23 ;
  wire \u2_Display/add167/c24 ;
  wire \u2_Display/add167/c25 ;
  wire \u2_Display/add167/c26 ;
  wire \u2_Display/add167/c27 ;
  wire \u2_Display/add167/c28 ;
  wire \u2_Display/add167/c29 ;
  wire \u2_Display/add167/c3 ;
  wire \u2_Display/add167/c30 ;
  wire \u2_Display/add167/c31 ;
  wire \u2_Display/add167/c4 ;
  wire \u2_Display/add167/c5 ;
  wire \u2_Display/add167/c6 ;
  wire \u2_Display/add167/c7 ;
  wire \u2_Display/add167/c8 ;
  wire \u2_Display/add167/c9 ;
  wire \u2_Display/add168/c0 ;
  wire \u2_Display/add168/c1 ;
  wire \u2_Display/add168/c10 ;
  wire \u2_Display/add168/c11 ;
  wire \u2_Display/add168/c12 ;
  wire \u2_Display/add168/c13 ;
  wire \u2_Display/add168/c14 ;
  wire \u2_Display/add168/c15 ;
  wire \u2_Display/add168/c16 ;
  wire \u2_Display/add168/c17 ;
  wire \u2_Display/add168/c18 ;
  wire \u2_Display/add168/c19 ;
  wire \u2_Display/add168/c2 ;
  wire \u2_Display/add168/c20 ;
  wire \u2_Display/add168/c21 ;
  wire \u2_Display/add168/c22 ;
  wire \u2_Display/add168/c23 ;
  wire \u2_Display/add168/c24 ;
  wire \u2_Display/add168/c25 ;
  wire \u2_Display/add168/c26 ;
  wire \u2_Display/add168/c27 ;
  wire \u2_Display/add168/c28 ;
  wire \u2_Display/add168/c29 ;
  wire \u2_Display/add168/c3 ;
  wire \u2_Display/add168/c30 ;
  wire \u2_Display/add168/c31 ;
  wire \u2_Display/add168/c4 ;
  wire \u2_Display/add168/c5 ;
  wire \u2_Display/add168/c6 ;
  wire \u2_Display/add168/c7 ;
  wire \u2_Display/add168/c8 ;
  wire \u2_Display/add168/c9 ;
  wire \u2_Display/add169/c0 ;
  wire \u2_Display/add169/c1 ;
  wire \u2_Display/add169/c10 ;
  wire \u2_Display/add169/c11 ;
  wire \u2_Display/add169/c12 ;
  wire \u2_Display/add169/c13 ;
  wire \u2_Display/add169/c14 ;
  wire \u2_Display/add169/c15 ;
  wire \u2_Display/add169/c16 ;
  wire \u2_Display/add169/c17 ;
  wire \u2_Display/add169/c18 ;
  wire \u2_Display/add169/c19 ;
  wire \u2_Display/add169/c2 ;
  wire \u2_Display/add169/c20 ;
  wire \u2_Display/add169/c21 ;
  wire \u2_Display/add169/c22 ;
  wire \u2_Display/add169/c23 ;
  wire \u2_Display/add169/c24 ;
  wire \u2_Display/add169/c25 ;
  wire \u2_Display/add169/c26 ;
  wire \u2_Display/add169/c27 ;
  wire \u2_Display/add169/c28 ;
  wire \u2_Display/add169/c29 ;
  wire \u2_Display/add169/c3 ;
  wire \u2_Display/add169/c30 ;
  wire \u2_Display/add169/c31 ;
  wire \u2_Display/add169/c4 ;
  wire \u2_Display/add169/c5 ;
  wire \u2_Display/add169/c6 ;
  wire \u2_Display/add169/c7 ;
  wire \u2_Display/add169/c8 ;
  wire \u2_Display/add169/c9 ;
  wire \u2_Display/add170/c0 ;
  wire \u2_Display/add170/c1 ;
  wire \u2_Display/add170/c10 ;
  wire \u2_Display/add170/c11 ;
  wire \u2_Display/add170/c12 ;
  wire \u2_Display/add170/c13 ;
  wire \u2_Display/add170/c14 ;
  wire \u2_Display/add170/c15 ;
  wire \u2_Display/add170/c16 ;
  wire \u2_Display/add170/c17 ;
  wire \u2_Display/add170/c18 ;
  wire \u2_Display/add170/c19 ;
  wire \u2_Display/add170/c2 ;
  wire \u2_Display/add170/c20 ;
  wire \u2_Display/add170/c21 ;
  wire \u2_Display/add170/c22 ;
  wire \u2_Display/add170/c23 ;
  wire \u2_Display/add170/c24 ;
  wire \u2_Display/add170/c25 ;
  wire \u2_Display/add170/c26 ;
  wire \u2_Display/add170/c27 ;
  wire \u2_Display/add170/c28 ;
  wire \u2_Display/add170/c29 ;
  wire \u2_Display/add170/c3 ;
  wire \u2_Display/add170/c30 ;
  wire \u2_Display/add170/c31 ;
  wire \u2_Display/add170/c4 ;
  wire \u2_Display/add170/c5 ;
  wire \u2_Display/add170/c6 ;
  wire \u2_Display/add170/c7 ;
  wire \u2_Display/add170/c8 ;
  wire \u2_Display/add170/c9 ;
  wire \u2_Display/add171/c0 ;
  wire \u2_Display/add171/c1 ;
  wire \u2_Display/add171/c10 ;
  wire \u2_Display/add171/c11 ;
  wire \u2_Display/add171/c12 ;
  wire \u2_Display/add171/c13 ;
  wire \u2_Display/add171/c14 ;
  wire \u2_Display/add171/c15 ;
  wire \u2_Display/add171/c16 ;
  wire \u2_Display/add171/c17 ;
  wire \u2_Display/add171/c18 ;
  wire \u2_Display/add171/c19 ;
  wire \u2_Display/add171/c2 ;
  wire \u2_Display/add171/c20 ;
  wire \u2_Display/add171/c21 ;
  wire \u2_Display/add171/c22 ;
  wire \u2_Display/add171/c23 ;
  wire \u2_Display/add171/c24 ;
  wire \u2_Display/add171/c25 ;
  wire \u2_Display/add171/c26 ;
  wire \u2_Display/add171/c27 ;
  wire \u2_Display/add171/c28 ;
  wire \u2_Display/add171/c29 ;
  wire \u2_Display/add171/c3 ;
  wire \u2_Display/add171/c30 ;
  wire \u2_Display/add171/c31 ;
  wire \u2_Display/add171/c4 ;
  wire \u2_Display/add171/c5 ;
  wire \u2_Display/add171/c6 ;
  wire \u2_Display/add171/c7 ;
  wire \u2_Display/add171/c8 ;
  wire \u2_Display/add171/c9 ;
  wire \u2_Display/add172/c0 ;
  wire \u2_Display/add172/c1 ;
  wire \u2_Display/add172/c2 ;
  wire \u2_Display/add172/c3 ;
  wire \u2_Display/add172/c4 ;
  wire \u2_Display/add172/c5 ;
  wire \u2_Display/add172/c6 ;
  wire \u2_Display/add172/c7 ;
  wire \u2_Display/add172/c8 ;
  wire \u2_Display/add172/c9 ;
  wire \u2_Display/add18/c0 ;
  wire \u2_Display/add18/c1 ;
  wire \u2_Display/add18/c10 ;
  wire \u2_Display/add18/c11 ;
  wire \u2_Display/add18/c12 ;
  wire \u2_Display/add18/c13 ;
  wire \u2_Display/add18/c14 ;
  wire \u2_Display/add18/c15 ;
  wire \u2_Display/add18/c16 ;
  wire \u2_Display/add18/c17 ;
  wire \u2_Display/add18/c18 ;
  wire \u2_Display/add18/c19 ;
  wire \u2_Display/add18/c2 ;
  wire \u2_Display/add18/c20 ;
  wire \u2_Display/add18/c21 ;
  wire \u2_Display/add18/c22 ;
  wire \u2_Display/add18/c23 ;
  wire \u2_Display/add18/c24 ;
  wire \u2_Display/add18/c25 ;
  wire \u2_Display/add18/c26 ;
  wire \u2_Display/add18/c27 ;
  wire \u2_Display/add18/c28 ;
  wire \u2_Display/add18/c29 ;
  wire \u2_Display/add18/c3 ;
  wire \u2_Display/add18/c30 ;
  wire \u2_Display/add18/c31 ;
  wire \u2_Display/add18/c4 ;
  wire \u2_Display/add18/c5 ;
  wire \u2_Display/add18/c6 ;
  wire \u2_Display/add18/c7 ;
  wire \u2_Display/add18/c8 ;
  wire \u2_Display/add18/c9 ;
  wire \u2_Display/add19/c0 ;
  wire \u2_Display/add19/c1 ;
  wire \u2_Display/add19/c10 ;
  wire \u2_Display/add19/c11 ;
  wire \u2_Display/add19/c12 ;
  wire \u2_Display/add19/c13 ;
  wire \u2_Display/add19/c14 ;
  wire \u2_Display/add19/c15 ;
  wire \u2_Display/add19/c16 ;
  wire \u2_Display/add19/c17 ;
  wire \u2_Display/add19/c18 ;
  wire \u2_Display/add19/c19 ;
  wire \u2_Display/add19/c2 ;
  wire \u2_Display/add19/c20 ;
  wire \u2_Display/add19/c21 ;
  wire \u2_Display/add19/c22 ;
  wire \u2_Display/add19/c23 ;
  wire \u2_Display/add19/c24 ;
  wire \u2_Display/add19/c25 ;
  wire \u2_Display/add19/c26 ;
  wire \u2_Display/add19/c27 ;
  wire \u2_Display/add19/c28 ;
  wire \u2_Display/add19/c29 ;
  wire \u2_Display/add19/c3 ;
  wire \u2_Display/add19/c30 ;
  wire \u2_Display/add19/c31 ;
  wire \u2_Display/add19/c4 ;
  wire \u2_Display/add19/c5 ;
  wire \u2_Display/add19/c6 ;
  wire \u2_Display/add19/c7 ;
  wire \u2_Display/add19/c8 ;
  wire \u2_Display/add19/c9 ;
  wire \u2_Display/add20/c0 ;
  wire \u2_Display/add20/c1 ;
  wire \u2_Display/add20/c10 ;
  wire \u2_Display/add20/c11 ;
  wire \u2_Display/add20/c12 ;
  wire \u2_Display/add20/c13 ;
  wire \u2_Display/add20/c14 ;
  wire \u2_Display/add20/c15 ;
  wire \u2_Display/add20/c16 ;
  wire \u2_Display/add20/c17 ;
  wire \u2_Display/add20/c18 ;
  wire \u2_Display/add20/c19 ;
  wire \u2_Display/add20/c2 ;
  wire \u2_Display/add20/c20 ;
  wire \u2_Display/add20/c21 ;
  wire \u2_Display/add20/c22 ;
  wire \u2_Display/add20/c23 ;
  wire \u2_Display/add20/c24 ;
  wire \u2_Display/add20/c25 ;
  wire \u2_Display/add20/c26 ;
  wire \u2_Display/add20/c27 ;
  wire \u2_Display/add20/c28 ;
  wire \u2_Display/add20/c29 ;
  wire \u2_Display/add20/c3 ;
  wire \u2_Display/add20/c30 ;
  wire \u2_Display/add20/c31 ;
  wire \u2_Display/add20/c4 ;
  wire \u2_Display/add20/c5 ;
  wire \u2_Display/add20/c6 ;
  wire \u2_Display/add20/c7 ;
  wire \u2_Display/add20/c8 ;
  wire \u2_Display/add20/c9 ;
  wire \u2_Display/add21/c0 ;
  wire \u2_Display/add21/c1 ;
  wire \u2_Display/add21/c10 ;
  wire \u2_Display/add21/c11 ;
  wire \u2_Display/add21/c12 ;
  wire \u2_Display/add21/c13 ;
  wire \u2_Display/add21/c14 ;
  wire \u2_Display/add21/c15 ;
  wire \u2_Display/add21/c16 ;
  wire \u2_Display/add21/c17 ;
  wire \u2_Display/add21/c18 ;
  wire \u2_Display/add21/c19 ;
  wire \u2_Display/add21/c2 ;
  wire \u2_Display/add21/c20 ;
  wire \u2_Display/add21/c21 ;
  wire \u2_Display/add21/c22 ;
  wire \u2_Display/add21/c23 ;
  wire \u2_Display/add21/c24 ;
  wire \u2_Display/add21/c25 ;
  wire \u2_Display/add21/c26 ;
  wire \u2_Display/add21/c27 ;
  wire \u2_Display/add21/c28 ;
  wire \u2_Display/add21/c29 ;
  wire \u2_Display/add21/c3 ;
  wire \u2_Display/add21/c30 ;
  wire \u2_Display/add21/c31 ;
  wire \u2_Display/add21/c4 ;
  wire \u2_Display/add21/c5 ;
  wire \u2_Display/add21/c6 ;
  wire \u2_Display/add21/c7 ;
  wire \u2_Display/add21/c8 ;
  wire \u2_Display/add21/c9 ;
  wire \u2_Display/add22/c0 ;
  wire \u2_Display/add22/c1 ;
  wire \u2_Display/add22/c10 ;
  wire \u2_Display/add22/c11 ;
  wire \u2_Display/add22/c12 ;
  wire \u2_Display/add22/c13 ;
  wire \u2_Display/add22/c14 ;
  wire \u2_Display/add22/c15 ;
  wire \u2_Display/add22/c16 ;
  wire \u2_Display/add22/c17 ;
  wire \u2_Display/add22/c18 ;
  wire \u2_Display/add22/c19 ;
  wire \u2_Display/add22/c2 ;
  wire \u2_Display/add22/c20 ;
  wire \u2_Display/add22/c21 ;
  wire \u2_Display/add22/c22 ;
  wire \u2_Display/add22/c23 ;
  wire \u2_Display/add22/c24 ;
  wire \u2_Display/add22/c25 ;
  wire \u2_Display/add22/c26 ;
  wire \u2_Display/add22/c27 ;
  wire \u2_Display/add22/c28 ;
  wire \u2_Display/add22/c29 ;
  wire \u2_Display/add22/c3 ;
  wire \u2_Display/add22/c30 ;
  wire \u2_Display/add22/c31 ;
  wire \u2_Display/add22/c4 ;
  wire \u2_Display/add22/c5 ;
  wire \u2_Display/add22/c6 ;
  wire \u2_Display/add22/c7 ;
  wire \u2_Display/add22/c8 ;
  wire \u2_Display/add22/c9 ;
  wire \u2_Display/add23/c0 ;
  wire \u2_Display/add23/c1 ;
  wire \u2_Display/add23/c10 ;
  wire \u2_Display/add23/c11 ;
  wire \u2_Display/add23/c12 ;
  wire \u2_Display/add23/c13 ;
  wire \u2_Display/add23/c14 ;
  wire \u2_Display/add23/c15 ;
  wire \u2_Display/add23/c16 ;
  wire \u2_Display/add23/c17 ;
  wire \u2_Display/add23/c18 ;
  wire \u2_Display/add23/c19 ;
  wire \u2_Display/add23/c2 ;
  wire \u2_Display/add23/c20 ;
  wire \u2_Display/add23/c21 ;
  wire \u2_Display/add23/c22 ;
  wire \u2_Display/add23/c23 ;
  wire \u2_Display/add23/c24 ;
  wire \u2_Display/add23/c25 ;
  wire \u2_Display/add23/c26 ;
  wire \u2_Display/add23/c27 ;
  wire \u2_Display/add23/c28 ;
  wire \u2_Display/add23/c29 ;
  wire \u2_Display/add23/c3 ;
  wire \u2_Display/add23/c30 ;
  wire \u2_Display/add23/c31 ;
  wire \u2_Display/add23/c4 ;
  wire \u2_Display/add23/c5 ;
  wire \u2_Display/add23/c6 ;
  wire \u2_Display/add23/c7 ;
  wire \u2_Display/add23/c8 ;
  wire \u2_Display/add23/c9 ;
  wire \u2_Display/add24/c0 ;
  wire \u2_Display/add24/c1 ;
  wire \u2_Display/add24/c10 ;
  wire \u2_Display/add24/c11 ;
  wire \u2_Display/add24/c12 ;
  wire \u2_Display/add24/c13 ;
  wire \u2_Display/add24/c14 ;
  wire \u2_Display/add24/c15 ;
  wire \u2_Display/add24/c16 ;
  wire \u2_Display/add24/c17 ;
  wire \u2_Display/add24/c18 ;
  wire \u2_Display/add24/c19 ;
  wire \u2_Display/add24/c2 ;
  wire \u2_Display/add24/c20 ;
  wire \u2_Display/add24/c21 ;
  wire \u2_Display/add24/c22 ;
  wire \u2_Display/add24/c23 ;
  wire \u2_Display/add24/c24 ;
  wire \u2_Display/add24/c25 ;
  wire \u2_Display/add24/c26 ;
  wire \u2_Display/add24/c27 ;
  wire \u2_Display/add24/c28 ;
  wire \u2_Display/add24/c29 ;
  wire \u2_Display/add24/c3 ;
  wire \u2_Display/add24/c30 ;
  wire \u2_Display/add24/c31 ;
  wire \u2_Display/add24/c4 ;
  wire \u2_Display/add24/c5 ;
  wire \u2_Display/add24/c6 ;
  wire \u2_Display/add24/c7 ;
  wire \u2_Display/add24/c8 ;
  wire \u2_Display/add24/c9 ;
  wire \u2_Display/add25/c0 ;
  wire \u2_Display/add25/c1 ;
  wire \u2_Display/add25/c10 ;
  wire \u2_Display/add25/c11 ;
  wire \u2_Display/add25/c12 ;
  wire \u2_Display/add25/c13 ;
  wire \u2_Display/add25/c14 ;
  wire \u2_Display/add25/c15 ;
  wire \u2_Display/add25/c16 ;
  wire \u2_Display/add25/c17 ;
  wire \u2_Display/add25/c18 ;
  wire \u2_Display/add25/c19 ;
  wire \u2_Display/add25/c2 ;
  wire \u2_Display/add25/c20 ;
  wire \u2_Display/add25/c21 ;
  wire \u2_Display/add25/c22 ;
  wire \u2_Display/add25/c23 ;
  wire \u2_Display/add25/c24 ;
  wire \u2_Display/add25/c25 ;
  wire \u2_Display/add25/c26 ;
  wire \u2_Display/add25/c27 ;
  wire \u2_Display/add25/c28 ;
  wire \u2_Display/add25/c29 ;
  wire \u2_Display/add25/c3 ;
  wire \u2_Display/add25/c30 ;
  wire \u2_Display/add25/c31 ;
  wire \u2_Display/add25/c4 ;
  wire \u2_Display/add25/c5 ;
  wire \u2_Display/add25/c6 ;
  wire \u2_Display/add25/c7 ;
  wire \u2_Display/add25/c8 ;
  wire \u2_Display/add25/c9 ;
  wire \u2_Display/add26/c0 ;
  wire \u2_Display/add26/c1 ;
  wire \u2_Display/add26/c10 ;
  wire \u2_Display/add26/c11 ;
  wire \u2_Display/add26/c12 ;
  wire \u2_Display/add26/c13 ;
  wire \u2_Display/add26/c14 ;
  wire \u2_Display/add26/c15 ;
  wire \u2_Display/add26/c16 ;
  wire \u2_Display/add26/c17 ;
  wire \u2_Display/add26/c18 ;
  wire \u2_Display/add26/c19 ;
  wire \u2_Display/add26/c2 ;
  wire \u2_Display/add26/c20 ;
  wire \u2_Display/add26/c21 ;
  wire \u2_Display/add26/c22 ;
  wire \u2_Display/add26/c23 ;
  wire \u2_Display/add26/c24 ;
  wire \u2_Display/add26/c25 ;
  wire \u2_Display/add26/c26 ;
  wire \u2_Display/add26/c27 ;
  wire \u2_Display/add26/c28 ;
  wire \u2_Display/add26/c29 ;
  wire \u2_Display/add26/c3 ;
  wire \u2_Display/add26/c30 ;
  wire \u2_Display/add26/c31 ;
  wire \u2_Display/add26/c4 ;
  wire \u2_Display/add26/c5 ;
  wire \u2_Display/add26/c6 ;
  wire \u2_Display/add26/c7 ;
  wire \u2_Display/add26/c8 ;
  wire \u2_Display/add26/c9 ;
  wire \u2_Display/add27/c0 ;
  wire \u2_Display/add27/c1 ;
  wire \u2_Display/add27/c10 ;
  wire \u2_Display/add27/c11 ;
  wire \u2_Display/add27/c12 ;
  wire \u2_Display/add27/c13 ;
  wire \u2_Display/add27/c14 ;
  wire \u2_Display/add27/c15 ;
  wire \u2_Display/add27/c16 ;
  wire \u2_Display/add27/c17 ;
  wire \u2_Display/add27/c18 ;
  wire \u2_Display/add27/c19 ;
  wire \u2_Display/add27/c2 ;
  wire \u2_Display/add27/c20 ;
  wire \u2_Display/add27/c21 ;
  wire \u2_Display/add27/c22 ;
  wire \u2_Display/add27/c23 ;
  wire \u2_Display/add27/c24 ;
  wire \u2_Display/add27/c25 ;
  wire \u2_Display/add27/c26 ;
  wire \u2_Display/add27/c27 ;
  wire \u2_Display/add27/c28 ;
  wire \u2_Display/add27/c29 ;
  wire \u2_Display/add27/c3 ;
  wire \u2_Display/add27/c30 ;
  wire \u2_Display/add27/c31 ;
  wire \u2_Display/add27/c4 ;
  wire \u2_Display/add27/c5 ;
  wire \u2_Display/add27/c6 ;
  wire \u2_Display/add27/c7 ;
  wire \u2_Display/add27/c8 ;
  wire \u2_Display/add27/c9 ;
  wire \u2_Display/add28/c0 ;
  wire \u2_Display/add28/c1 ;
  wire \u2_Display/add28/c10 ;
  wire \u2_Display/add28/c11 ;
  wire \u2_Display/add28/c12 ;
  wire \u2_Display/add28/c13 ;
  wire \u2_Display/add28/c14 ;
  wire \u2_Display/add28/c15 ;
  wire \u2_Display/add28/c16 ;
  wire \u2_Display/add28/c17 ;
  wire \u2_Display/add28/c18 ;
  wire \u2_Display/add28/c19 ;
  wire \u2_Display/add28/c2 ;
  wire \u2_Display/add28/c20 ;
  wire \u2_Display/add28/c21 ;
  wire \u2_Display/add28/c22 ;
  wire \u2_Display/add28/c23 ;
  wire \u2_Display/add28/c24 ;
  wire \u2_Display/add28/c25 ;
  wire \u2_Display/add28/c26 ;
  wire \u2_Display/add28/c27 ;
  wire \u2_Display/add28/c28 ;
  wire \u2_Display/add28/c29 ;
  wire \u2_Display/add28/c3 ;
  wire \u2_Display/add28/c30 ;
  wire \u2_Display/add28/c31 ;
  wire \u2_Display/add28/c4 ;
  wire \u2_Display/add28/c5 ;
  wire \u2_Display/add28/c6 ;
  wire \u2_Display/add28/c7 ;
  wire \u2_Display/add28/c8 ;
  wire \u2_Display/add28/c9 ;
  wire \u2_Display/add29/c0 ;
  wire \u2_Display/add29/c1 ;
  wire \u2_Display/add29/c10 ;
  wire \u2_Display/add29/c11 ;
  wire \u2_Display/add29/c12 ;
  wire \u2_Display/add29/c13 ;
  wire \u2_Display/add29/c14 ;
  wire \u2_Display/add29/c15 ;
  wire \u2_Display/add29/c16 ;
  wire \u2_Display/add29/c17 ;
  wire \u2_Display/add29/c18 ;
  wire \u2_Display/add29/c19 ;
  wire \u2_Display/add29/c2 ;
  wire \u2_Display/add29/c20 ;
  wire \u2_Display/add29/c21 ;
  wire \u2_Display/add29/c22 ;
  wire \u2_Display/add29/c23 ;
  wire \u2_Display/add29/c24 ;
  wire \u2_Display/add29/c25 ;
  wire \u2_Display/add29/c26 ;
  wire \u2_Display/add29/c27 ;
  wire \u2_Display/add29/c28 ;
  wire \u2_Display/add29/c29 ;
  wire \u2_Display/add29/c3 ;
  wire \u2_Display/add29/c30 ;
  wire \u2_Display/add29/c31 ;
  wire \u2_Display/add29/c4 ;
  wire \u2_Display/add29/c5 ;
  wire \u2_Display/add29/c6 ;
  wire \u2_Display/add29/c7 ;
  wire \u2_Display/add29/c8 ;
  wire \u2_Display/add29/c9 ;
  wire \u2_Display/add2_2/c0 ;
  wire \u2_Display/add2_2/c1 ;
  wire \u2_Display/add2_2/c2 ;
  wire \u2_Display/add2_2/c3 ;
  wire \u2_Display/add2_2_co ;
  wire \u2_Display/add30/c0 ;
  wire \u2_Display/add30/c1 ;
  wire \u2_Display/add30/c10 ;
  wire \u2_Display/add30/c11 ;
  wire \u2_Display/add30/c12 ;
  wire \u2_Display/add30/c13 ;
  wire \u2_Display/add30/c14 ;
  wire \u2_Display/add30/c15 ;
  wire \u2_Display/add30/c16 ;
  wire \u2_Display/add30/c17 ;
  wire \u2_Display/add30/c18 ;
  wire \u2_Display/add30/c19 ;
  wire \u2_Display/add30/c2 ;
  wire \u2_Display/add30/c20 ;
  wire \u2_Display/add30/c21 ;
  wire \u2_Display/add30/c22 ;
  wire \u2_Display/add30/c23 ;
  wire \u2_Display/add30/c24 ;
  wire \u2_Display/add30/c25 ;
  wire \u2_Display/add30/c26 ;
  wire \u2_Display/add30/c27 ;
  wire \u2_Display/add30/c28 ;
  wire \u2_Display/add30/c29 ;
  wire \u2_Display/add30/c3 ;
  wire \u2_Display/add30/c30 ;
  wire \u2_Display/add30/c31 ;
  wire \u2_Display/add30/c4 ;
  wire \u2_Display/add30/c5 ;
  wire \u2_Display/add30/c6 ;
  wire \u2_Display/add30/c7 ;
  wire \u2_Display/add30/c8 ;
  wire \u2_Display/add30/c9 ;
  wire \u2_Display/add31/c0 ;
  wire \u2_Display/add31/c1 ;
  wire \u2_Display/add31/c10 ;
  wire \u2_Display/add31/c11 ;
  wire \u2_Display/add31/c12 ;
  wire \u2_Display/add31/c13 ;
  wire \u2_Display/add31/c14 ;
  wire \u2_Display/add31/c15 ;
  wire \u2_Display/add31/c16 ;
  wire \u2_Display/add31/c17 ;
  wire \u2_Display/add31/c18 ;
  wire \u2_Display/add31/c19 ;
  wire \u2_Display/add31/c2 ;
  wire \u2_Display/add31/c20 ;
  wire \u2_Display/add31/c21 ;
  wire \u2_Display/add31/c22 ;
  wire \u2_Display/add31/c23 ;
  wire \u2_Display/add31/c24 ;
  wire \u2_Display/add31/c25 ;
  wire \u2_Display/add31/c26 ;
  wire \u2_Display/add31/c27 ;
  wire \u2_Display/add31/c28 ;
  wire \u2_Display/add31/c29 ;
  wire \u2_Display/add31/c3 ;
  wire \u2_Display/add31/c30 ;
  wire \u2_Display/add31/c31 ;
  wire \u2_Display/add31/c4 ;
  wire \u2_Display/add31/c5 ;
  wire \u2_Display/add31/c6 ;
  wire \u2_Display/add31/c7 ;
  wire \u2_Display/add31/c8 ;
  wire \u2_Display/add31/c9 ;
  wire \u2_Display/add32/c0 ;
  wire \u2_Display/add32/c1 ;
  wire \u2_Display/add32/c10 ;
  wire \u2_Display/add32/c11 ;
  wire \u2_Display/add32/c12 ;
  wire \u2_Display/add32/c13 ;
  wire \u2_Display/add32/c14 ;
  wire \u2_Display/add32/c15 ;
  wire \u2_Display/add32/c16 ;
  wire \u2_Display/add32/c17 ;
  wire \u2_Display/add32/c18 ;
  wire \u2_Display/add32/c19 ;
  wire \u2_Display/add32/c2 ;
  wire \u2_Display/add32/c20 ;
  wire \u2_Display/add32/c21 ;
  wire \u2_Display/add32/c22 ;
  wire \u2_Display/add32/c23 ;
  wire \u2_Display/add32/c24 ;
  wire \u2_Display/add32/c25 ;
  wire \u2_Display/add32/c26 ;
  wire \u2_Display/add32/c27 ;
  wire \u2_Display/add32/c28 ;
  wire \u2_Display/add32/c29 ;
  wire \u2_Display/add32/c3 ;
  wire \u2_Display/add32/c30 ;
  wire \u2_Display/add32/c31 ;
  wire \u2_Display/add32/c4 ;
  wire \u2_Display/add32/c5 ;
  wire \u2_Display/add32/c6 ;
  wire \u2_Display/add32/c7 ;
  wire \u2_Display/add32/c8 ;
  wire \u2_Display/add32/c9 ;
  wire \u2_Display/add33/c0 ;
  wire \u2_Display/add33/c1 ;
  wire \u2_Display/add33/c10 ;
  wire \u2_Display/add33/c11 ;
  wire \u2_Display/add33/c12 ;
  wire \u2_Display/add33/c13 ;
  wire \u2_Display/add33/c14 ;
  wire \u2_Display/add33/c15 ;
  wire \u2_Display/add33/c16 ;
  wire \u2_Display/add33/c17 ;
  wire \u2_Display/add33/c18 ;
  wire \u2_Display/add33/c19 ;
  wire \u2_Display/add33/c2 ;
  wire \u2_Display/add33/c20 ;
  wire \u2_Display/add33/c21 ;
  wire \u2_Display/add33/c22 ;
  wire \u2_Display/add33/c23 ;
  wire \u2_Display/add33/c24 ;
  wire \u2_Display/add33/c25 ;
  wire \u2_Display/add33/c26 ;
  wire \u2_Display/add33/c27 ;
  wire \u2_Display/add33/c28 ;
  wire \u2_Display/add33/c29 ;
  wire \u2_Display/add33/c3 ;
  wire \u2_Display/add33/c30 ;
  wire \u2_Display/add33/c31 ;
  wire \u2_Display/add33/c4 ;
  wire \u2_Display/add33/c5 ;
  wire \u2_Display/add33/c6 ;
  wire \u2_Display/add33/c7 ;
  wire \u2_Display/add33/c8 ;
  wire \u2_Display/add33/c9 ;
  wire \u2_Display/add34/c0 ;
  wire \u2_Display/add34/c1 ;
  wire \u2_Display/add34/c10 ;
  wire \u2_Display/add34/c11 ;
  wire \u2_Display/add34/c12 ;
  wire \u2_Display/add34/c13 ;
  wire \u2_Display/add34/c14 ;
  wire \u2_Display/add34/c15 ;
  wire \u2_Display/add34/c16 ;
  wire \u2_Display/add34/c17 ;
  wire \u2_Display/add34/c18 ;
  wire \u2_Display/add34/c19 ;
  wire \u2_Display/add34/c2 ;
  wire \u2_Display/add34/c20 ;
  wire \u2_Display/add34/c21 ;
  wire \u2_Display/add34/c22 ;
  wire \u2_Display/add34/c23 ;
  wire \u2_Display/add34/c24 ;
  wire \u2_Display/add34/c25 ;
  wire \u2_Display/add34/c26 ;
  wire \u2_Display/add34/c27 ;
  wire \u2_Display/add34/c28 ;
  wire \u2_Display/add34/c29 ;
  wire \u2_Display/add34/c3 ;
  wire \u2_Display/add34/c30 ;
  wire \u2_Display/add34/c31 ;
  wire \u2_Display/add34/c4 ;
  wire \u2_Display/add34/c5 ;
  wire \u2_Display/add34/c6 ;
  wire \u2_Display/add34/c7 ;
  wire \u2_Display/add34/c8 ;
  wire \u2_Display/add34/c9 ;
  wire \u2_Display/add35/c0 ;
  wire \u2_Display/add35/c1 ;
  wire \u2_Display/add35/c10 ;
  wire \u2_Display/add35/c11 ;
  wire \u2_Display/add35/c12 ;
  wire \u2_Display/add35/c13 ;
  wire \u2_Display/add35/c14 ;
  wire \u2_Display/add35/c15 ;
  wire \u2_Display/add35/c16 ;
  wire \u2_Display/add35/c17 ;
  wire \u2_Display/add35/c18 ;
  wire \u2_Display/add35/c19 ;
  wire \u2_Display/add35/c2 ;
  wire \u2_Display/add35/c20 ;
  wire \u2_Display/add35/c21 ;
  wire \u2_Display/add35/c22 ;
  wire \u2_Display/add35/c23 ;
  wire \u2_Display/add35/c24 ;
  wire \u2_Display/add35/c25 ;
  wire \u2_Display/add35/c26 ;
  wire \u2_Display/add35/c27 ;
  wire \u2_Display/add35/c28 ;
  wire \u2_Display/add35/c29 ;
  wire \u2_Display/add35/c3 ;
  wire \u2_Display/add35/c30 ;
  wire \u2_Display/add35/c31 ;
  wire \u2_Display/add35/c4 ;
  wire \u2_Display/add35/c5 ;
  wire \u2_Display/add35/c6 ;
  wire \u2_Display/add35/c7 ;
  wire \u2_Display/add35/c8 ;
  wire \u2_Display/add35/c9 ;
  wire \u2_Display/add36/c0 ;
  wire \u2_Display/add36/c1 ;
  wire \u2_Display/add36/c10 ;
  wire \u2_Display/add36/c11 ;
  wire \u2_Display/add36/c12 ;
  wire \u2_Display/add36/c13 ;
  wire \u2_Display/add36/c14 ;
  wire \u2_Display/add36/c15 ;
  wire \u2_Display/add36/c16 ;
  wire \u2_Display/add36/c17 ;
  wire \u2_Display/add36/c18 ;
  wire \u2_Display/add36/c19 ;
  wire \u2_Display/add36/c2 ;
  wire \u2_Display/add36/c20 ;
  wire \u2_Display/add36/c21 ;
  wire \u2_Display/add36/c22 ;
  wire \u2_Display/add36/c23 ;
  wire \u2_Display/add36/c24 ;
  wire \u2_Display/add36/c25 ;
  wire \u2_Display/add36/c26 ;
  wire \u2_Display/add36/c27 ;
  wire \u2_Display/add36/c28 ;
  wire \u2_Display/add36/c29 ;
  wire \u2_Display/add36/c3 ;
  wire \u2_Display/add36/c30 ;
  wire \u2_Display/add36/c31 ;
  wire \u2_Display/add36/c4 ;
  wire \u2_Display/add36/c5 ;
  wire \u2_Display/add36/c6 ;
  wire \u2_Display/add36/c7 ;
  wire \u2_Display/add36/c8 ;
  wire \u2_Display/add36/c9 ;
  wire \u2_Display/add37/c0 ;
  wire \u2_Display/add37/c1 ;
  wire \u2_Display/add37/c10 ;
  wire \u2_Display/add37/c11 ;
  wire \u2_Display/add37/c12 ;
  wire \u2_Display/add37/c13 ;
  wire \u2_Display/add37/c14 ;
  wire \u2_Display/add37/c15 ;
  wire \u2_Display/add37/c16 ;
  wire \u2_Display/add37/c17 ;
  wire \u2_Display/add37/c18 ;
  wire \u2_Display/add37/c19 ;
  wire \u2_Display/add37/c2 ;
  wire \u2_Display/add37/c20 ;
  wire \u2_Display/add37/c21 ;
  wire \u2_Display/add37/c22 ;
  wire \u2_Display/add37/c23 ;
  wire \u2_Display/add37/c24 ;
  wire \u2_Display/add37/c25 ;
  wire \u2_Display/add37/c26 ;
  wire \u2_Display/add37/c27 ;
  wire \u2_Display/add37/c28 ;
  wire \u2_Display/add37/c29 ;
  wire \u2_Display/add37/c3 ;
  wire \u2_Display/add37/c30 ;
  wire \u2_Display/add37/c31 ;
  wire \u2_Display/add37/c4 ;
  wire \u2_Display/add37/c5 ;
  wire \u2_Display/add37/c6 ;
  wire \u2_Display/add37/c7 ;
  wire \u2_Display/add37/c8 ;
  wire \u2_Display/add37/c9 ;
  wire \u2_Display/add38/c0 ;
  wire \u2_Display/add38/c1 ;
  wire \u2_Display/add38/c10 ;
  wire \u2_Display/add38/c11 ;
  wire \u2_Display/add38/c12 ;
  wire \u2_Display/add38/c13 ;
  wire \u2_Display/add38/c14 ;
  wire \u2_Display/add38/c15 ;
  wire \u2_Display/add38/c16 ;
  wire \u2_Display/add38/c17 ;
  wire \u2_Display/add38/c18 ;
  wire \u2_Display/add38/c19 ;
  wire \u2_Display/add38/c2 ;
  wire \u2_Display/add38/c20 ;
  wire \u2_Display/add38/c21 ;
  wire \u2_Display/add38/c22 ;
  wire \u2_Display/add38/c23 ;
  wire \u2_Display/add38/c24 ;
  wire \u2_Display/add38/c25 ;
  wire \u2_Display/add38/c26 ;
  wire \u2_Display/add38/c27 ;
  wire \u2_Display/add38/c28 ;
  wire \u2_Display/add38/c29 ;
  wire \u2_Display/add38/c3 ;
  wire \u2_Display/add38/c30 ;
  wire \u2_Display/add38/c31 ;
  wire \u2_Display/add38/c4 ;
  wire \u2_Display/add38/c5 ;
  wire \u2_Display/add38/c6 ;
  wire \u2_Display/add38/c7 ;
  wire \u2_Display/add38/c8 ;
  wire \u2_Display/add38/c9 ;
  wire \u2_Display/add39/c0 ;
  wire \u2_Display/add39/c1 ;
  wire \u2_Display/add39/c10 ;
  wire \u2_Display/add39/c11 ;
  wire \u2_Display/add39/c12 ;
  wire \u2_Display/add39/c13 ;
  wire \u2_Display/add39/c14 ;
  wire \u2_Display/add39/c15 ;
  wire \u2_Display/add39/c16 ;
  wire \u2_Display/add39/c17 ;
  wire \u2_Display/add39/c18 ;
  wire \u2_Display/add39/c19 ;
  wire \u2_Display/add39/c2 ;
  wire \u2_Display/add39/c20 ;
  wire \u2_Display/add39/c21 ;
  wire \u2_Display/add39/c22 ;
  wire \u2_Display/add39/c23 ;
  wire \u2_Display/add39/c24 ;
  wire \u2_Display/add39/c25 ;
  wire \u2_Display/add39/c26 ;
  wire \u2_Display/add39/c27 ;
  wire \u2_Display/add39/c28 ;
  wire \u2_Display/add39/c29 ;
  wire \u2_Display/add39/c3 ;
  wire \u2_Display/add39/c30 ;
  wire \u2_Display/add39/c31 ;
  wire \u2_Display/add39/c4 ;
  wire \u2_Display/add39/c5 ;
  wire \u2_Display/add39/c6 ;
  wire \u2_Display/add39/c7 ;
  wire \u2_Display/add39/c8 ;
  wire \u2_Display/add39/c9 ;
  wire \u2_Display/add40/c0 ;
  wire \u2_Display/add40/c1 ;
  wire \u2_Display/add40/c2 ;
  wire \u2_Display/add40/c3 ;
  wire \u2_Display/add40/c4 ;
  wire \u2_Display/add40/c5 ;
  wire \u2_Display/add40/c6 ;
  wire \u2_Display/add40/c7 ;
  wire \u2_Display/add40/c8 ;
  wire \u2_Display/add40/c9 ;
  wire \u2_Display/add4_2/c0 ;
  wire \u2_Display/add4_2/c1 ;
  wire \u2_Display/add4_2/c2 ;
  wire \u2_Display/add4_2/c3 ;
  wire \u2_Display/add4_2/c4 ;
  wire \u2_Display/add4_2_co ;
  wire \u2_Display/add51/c0 ;
  wire \u2_Display/add51/c1 ;
  wire \u2_Display/add51/c10 ;
  wire \u2_Display/add51/c11 ;
  wire \u2_Display/add51/c12 ;
  wire \u2_Display/add51/c13 ;
  wire \u2_Display/add51/c14 ;
  wire \u2_Display/add51/c15 ;
  wire \u2_Display/add51/c16 ;
  wire \u2_Display/add51/c17 ;
  wire \u2_Display/add51/c18 ;
  wire \u2_Display/add51/c19 ;
  wire \u2_Display/add51/c2 ;
  wire \u2_Display/add51/c20 ;
  wire \u2_Display/add51/c21 ;
  wire \u2_Display/add51/c22 ;
  wire \u2_Display/add51/c23 ;
  wire \u2_Display/add51/c24 ;
  wire \u2_Display/add51/c25 ;
  wire \u2_Display/add51/c26 ;
  wire \u2_Display/add51/c27 ;
  wire \u2_Display/add51/c28 ;
  wire \u2_Display/add51/c29 ;
  wire \u2_Display/add51/c3 ;
  wire \u2_Display/add51/c30 ;
  wire \u2_Display/add51/c31 ;
  wire \u2_Display/add51/c4 ;
  wire \u2_Display/add51/c5 ;
  wire \u2_Display/add51/c6 ;
  wire \u2_Display/add51/c7 ;
  wire \u2_Display/add51/c8 ;
  wire \u2_Display/add51/c9 ;
  wire \u2_Display/add52/c0 ;
  wire \u2_Display/add52/c1 ;
  wire \u2_Display/add52/c10 ;
  wire \u2_Display/add52/c11 ;
  wire \u2_Display/add52/c12 ;
  wire \u2_Display/add52/c13 ;
  wire \u2_Display/add52/c14 ;
  wire \u2_Display/add52/c15 ;
  wire \u2_Display/add52/c16 ;
  wire \u2_Display/add52/c17 ;
  wire \u2_Display/add52/c18 ;
  wire \u2_Display/add52/c19 ;
  wire \u2_Display/add52/c2 ;
  wire \u2_Display/add52/c20 ;
  wire \u2_Display/add52/c21 ;
  wire \u2_Display/add52/c22 ;
  wire \u2_Display/add52/c23 ;
  wire \u2_Display/add52/c24 ;
  wire \u2_Display/add52/c25 ;
  wire \u2_Display/add52/c26 ;
  wire \u2_Display/add52/c27 ;
  wire \u2_Display/add52/c28 ;
  wire \u2_Display/add52/c29 ;
  wire \u2_Display/add52/c3 ;
  wire \u2_Display/add52/c30 ;
  wire \u2_Display/add52/c31 ;
  wire \u2_Display/add52/c4 ;
  wire \u2_Display/add52/c5 ;
  wire \u2_Display/add52/c6 ;
  wire \u2_Display/add52/c7 ;
  wire \u2_Display/add52/c8 ;
  wire \u2_Display/add52/c9 ;
  wire \u2_Display/add53/c0 ;
  wire \u2_Display/add53/c1 ;
  wire \u2_Display/add53/c10 ;
  wire \u2_Display/add53/c11 ;
  wire \u2_Display/add53/c12 ;
  wire \u2_Display/add53/c13 ;
  wire \u2_Display/add53/c14 ;
  wire \u2_Display/add53/c15 ;
  wire \u2_Display/add53/c16 ;
  wire \u2_Display/add53/c17 ;
  wire \u2_Display/add53/c18 ;
  wire \u2_Display/add53/c19 ;
  wire \u2_Display/add53/c2 ;
  wire \u2_Display/add53/c20 ;
  wire \u2_Display/add53/c21 ;
  wire \u2_Display/add53/c22 ;
  wire \u2_Display/add53/c23 ;
  wire \u2_Display/add53/c24 ;
  wire \u2_Display/add53/c25 ;
  wire \u2_Display/add53/c26 ;
  wire \u2_Display/add53/c27 ;
  wire \u2_Display/add53/c28 ;
  wire \u2_Display/add53/c29 ;
  wire \u2_Display/add53/c3 ;
  wire \u2_Display/add53/c30 ;
  wire \u2_Display/add53/c31 ;
  wire \u2_Display/add53/c4 ;
  wire \u2_Display/add53/c5 ;
  wire \u2_Display/add53/c6 ;
  wire \u2_Display/add53/c7 ;
  wire \u2_Display/add53/c8 ;
  wire \u2_Display/add53/c9 ;
  wire \u2_Display/add54/c0 ;
  wire \u2_Display/add54/c1 ;
  wire \u2_Display/add54/c10 ;
  wire \u2_Display/add54/c11 ;
  wire \u2_Display/add54/c12 ;
  wire \u2_Display/add54/c13 ;
  wire \u2_Display/add54/c14 ;
  wire \u2_Display/add54/c15 ;
  wire \u2_Display/add54/c16 ;
  wire \u2_Display/add54/c17 ;
  wire \u2_Display/add54/c18 ;
  wire \u2_Display/add54/c19 ;
  wire \u2_Display/add54/c2 ;
  wire \u2_Display/add54/c20 ;
  wire \u2_Display/add54/c21 ;
  wire \u2_Display/add54/c22 ;
  wire \u2_Display/add54/c23 ;
  wire \u2_Display/add54/c24 ;
  wire \u2_Display/add54/c25 ;
  wire \u2_Display/add54/c26 ;
  wire \u2_Display/add54/c27 ;
  wire \u2_Display/add54/c28 ;
  wire \u2_Display/add54/c29 ;
  wire \u2_Display/add54/c3 ;
  wire \u2_Display/add54/c30 ;
  wire \u2_Display/add54/c31 ;
  wire \u2_Display/add54/c4 ;
  wire \u2_Display/add54/c5 ;
  wire \u2_Display/add54/c6 ;
  wire \u2_Display/add54/c7 ;
  wire \u2_Display/add54/c8 ;
  wire \u2_Display/add54/c9 ;
  wire \u2_Display/add55/c0 ;
  wire \u2_Display/add55/c1 ;
  wire \u2_Display/add55/c10 ;
  wire \u2_Display/add55/c11 ;
  wire \u2_Display/add55/c12 ;
  wire \u2_Display/add55/c13 ;
  wire \u2_Display/add55/c14 ;
  wire \u2_Display/add55/c15 ;
  wire \u2_Display/add55/c16 ;
  wire \u2_Display/add55/c17 ;
  wire \u2_Display/add55/c18 ;
  wire \u2_Display/add55/c19 ;
  wire \u2_Display/add55/c2 ;
  wire \u2_Display/add55/c20 ;
  wire \u2_Display/add55/c21 ;
  wire \u2_Display/add55/c22 ;
  wire \u2_Display/add55/c23 ;
  wire \u2_Display/add55/c24 ;
  wire \u2_Display/add55/c25 ;
  wire \u2_Display/add55/c26 ;
  wire \u2_Display/add55/c27 ;
  wire \u2_Display/add55/c28 ;
  wire \u2_Display/add55/c29 ;
  wire \u2_Display/add55/c3 ;
  wire \u2_Display/add55/c30 ;
  wire \u2_Display/add55/c31 ;
  wire \u2_Display/add55/c4 ;
  wire \u2_Display/add55/c5 ;
  wire \u2_Display/add55/c6 ;
  wire \u2_Display/add55/c7 ;
  wire \u2_Display/add55/c8 ;
  wire \u2_Display/add55/c9 ;
  wire \u2_Display/add56/c0 ;
  wire \u2_Display/add56/c1 ;
  wire \u2_Display/add56/c10 ;
  wire \u2_Display/add56/c11 ;
  wire \u2_Display/add56/c12 ;
  wire \u2_Display/add56/c13 ;
  wire \u2_Display/add56/c14 ;
  wire \u2_Display/add56/c15 ;
  wire \u2_Display/add56/c16 ;
  wire \u2_Display/add56/c17 ;
  wire \u2_Display/add56/c18 ;
  wire \u2_Display/add56/c19 ;
  wire \u2_Display/add56/c2 ;
  wire \u2_Display/add56/c20 ;
  wire \u2_Display/add56/c21 ;
  wire \u2_Display/add56/c22 ;
  wire \u2_Display/add56/c23 ;
  wire \u2_Display/add56/c24 ;
  wire \u2_Display/add56/c25 ;
  wire \u2_Display/add56/c26 ;
  wire \u2_Display/add56/c27 ;
  wire \u2_Display/add56/c28 ;
  wire \u2_Display/add56/c29 ;
  wire \u2_Display/add56/c3 ;
  wire \u2_Display/add56/c30 ;
  wire \u2_Display/add56/c31 ;
  wire \u2_Display/add56/c4 ;
  wire \u2_Display/add56/c5 ;
  wire \u2_Display/add56/c6 ;
  wire \u2_Display/add56/c7 ;
  wire \u2_Display/add56/c8 ;
  wire \u2_Display/add56/c9 ;
  wire \u2_Display/add57/c0 ;
  wire \u2_Display/add57/c1 ;
  wire \u2_Display/add57/c10 ;
  wire \u2_Display/add57/c11 ;
  wire \u2_Display/add57/c12 ;
  wire \u2_Display/add57/c13 ;
  wire \u2_Display/add57/c14 ;
  wire \u2_Display/add57/c15 ;
  wire \u2_Display/add57/c16 ;
  wire \u2_Display/add57/c17 ;
  wire \u2_Display/add57/c18 ;
  wire \u2_Display/add57/c19 ;
  wire \u2_Display/add57/c2 ;
  wire \u2_Display/add57/c20 ;
  wire \u2_Display/add57/c21 ;
  wire \u2_Display/add57/c22 ;
  wire \u2_Display/add57/c23 ;
  wire \u2_Display/add57/c24 ;
  wire \u2_Display/add57/c25 ;
  wire \u2_Display/add57/c26 ;
  wire \u2_Display/add57/c27 ;
  wire \u2_Display/add57/c28 ;
  wire \u2_Display/add57/c29 ;
  wire \u2_Display/add57/c3 ;
  wire \u2_Display/add57/c30 ;
  wire \u2_Display/add57/c31 ;
  wire \u2_Display/add57/c4 ;
  wire \u2_Display/add57/c5 ;
  wire \u2_Display/add57/c6 ;
  wire \u2_Display/add57/c7 ;
  wire \u2_Display/add57/c8 ;
  wire \u2_Display/add57/c9 ;
  wire \u2_Display/add58/c0 ;
  wire \u2_Display/add58/c1 ;
  wire \u2_Display/add58/c10 ;
  wire \u2_Display/add58/c11 ;
  wire \u2_Display/add58/c12 ;
  wire \u2_Display/add58/c13 ;
  wire \u2_Display/add58/c14 ;
  wire \u2_Display/add58/c15 ;
  wire \u2_Display/add58/c16 ;
  wire \u2_Display/add58/c17 ;
  wire \u2_Display/add58/c18 ;
  wire \u2_Display/add58/c19 ;
  wire \u2_Display/add58/c2 ;
  wire \u2_Display/add58/c20 ;
  wire \u2_Display/add58/c21 ;
  wire \u2_Display/add58/c22 ;
  wire \u2_Display/add58/c23 ;
  wire \u2_Display/add58/c24 ;
  wire \u2_Display/add58/c25 ;
  wire \u2_Display/add58/c26 ;
  wire \u2_Display/add58/c27 ;
  wire \u2_Display/add58/c28 ;
  wire \u2_Display/add58/c29 ;
  wire \u2_Display/add58/c3 ;
  wire \u2_Display/add58/c30 ;
  wire \u2_Display/add58/c31 ;
  wire \u2_Display/add58/c4 ;
  wire \u2_Display/add58/c5 ;
  wire \u2_Display/add58/c6 ;
  wire \u2_Display/add58/c7 ;
  wire \u2_Display/add58/c8 ;
  wire \u2_Display/add58/c9 ;
  wire \u2_Display/add59/c0 ;
  wire \u2_Display/add59/c1 ;
  wire \u2_Display/add59/c10 ;
  wire \u2_Display/add59/c11 ;
  wire \u2_Display/add59/c12 ;
  wire \u2_Display/add59/c13 ;
  wire \u2_Display/add59/c14 ;
  wire \u2_Display/add59/c15 ;
  wire \u2_Display/add59/c16 ;
  wire \u2_Display/add59/c17 ;
  wire \u2_Display/add59/c18 ;
  wire \u2_Display/add59/c19 ;
  wire \u2_Display/add59/c2 ;
  wire \u2_Display/add59/c20 ;
  wire \u2_Display/add59/c21 ;
  wire \u2_Display/add59/c22 ;
  wire \u2_Display/add59/c23 ;
  wire \u2_Display/add59/c24 ;
  wire \u2_Display/add59/c25 ;
  wire \u2_Display/add59/c26 ;
  wire \u2_Display/add59/c27 ;
  wire \u2_Display/add59/c28 ;
  wire \u2_Display/add59/c29 ;
  wire \u2_Display/add59/c3 ;
  wire \u2_Display/add59/c30 ;
  wire \u2_Display/add59/c31 ;
  wire \u2_Display/add59/c4 ;
  wire \u2_Display/add59/c5 ;
  wire \u2_Display/add59/c6 ;
  wire \u2_Display/add59/c7 ;
  wire \u2_Display/add59/c8 ;
  wire \u2_Display/add59/c9 ;
  wire \u2_Display/add60/c0 ;
  wire \u2_Display/add60/c1 ;
  wire \u2_Display/add60/c10 ;
  wire \u2_Display/add60/c11 ;
  wire \u2_Display/add60/c12 ;
  wire \u2_Display/add60/c13 ;
  wire \u2_Display/add60/c14 ;
  wire \u2_Display/add60/c15 ;
  wire \u2_Display/add60/c16 ;
  wire \u2_Display/add60/c17 ;
  wire \u2_Display/add60/c18 ;
  wire \u2_Display/add60/c19 ;
  wire \u2_Display/add60/c2 ;
  wire \u2_Display/add60/c20 ;
  wire \u2_Display/add60/c21 ;
  wire \u2_Display/add60/c22 ;
  wire \u2_Display/add60/c23 ;
  wire \u2_Display/add60/c24 ;
  wire \u2_Display/add60/c25 ;
  wire \u2_Display/add60/c26 ;
  wire \u2_Display/add60/c27 ;
  wire \u2_Display/add60/c28 ;
  wire \u2_Display/add60/c29 ;
  wire \u2_Display/add60/c3 ;
  wire \u2_Display/add60/c30 ;
  wire \u2_Display/add60/c31 ;
  wire \u2_Display/add60/c4 ;
  wire \u2_Display/add60/c5 ;
  wire \u2_Display/add60/c6 ;
  wire \u2_Display/add60/c7 ;
  wire \u2_Display/add60/c8 ;
  wire \u2_Display/add60/c9 ;
  wire \u2_Display/add61/c0 ;
  wire \u2_Display/add61/c1 ;
  wire \u2_Display/add61/c10 ;
  wire \u2_Display/add61/c11 ;
  wire \u2_Display/add61/c12 ;
  wire \u2_Display/add61/c13 ;
  wire \u2_Display/add61/c14 ;
  wire \u2_Display/add61/c15 ;
  wire \u2_Display/add61/c16 ;
  wire \u2_Display/add61/c17 ;
  wire \u2_Display/add61/c18 ;
  wire \u2_Display/add61/c19 ;
  wire \u2_Display/add61/c2 ;
  wire \u2_Display/add61/c20 ;
  wire \u2_Display/add61/c21 ;
  wire \u2_Display/add61/c22 ;
  wire \u2_Display/add61/c23 ;
  wire \u2_Display/add61/c24 ;
  wire \u2_Display/add61/c25 ;
  wire \u2_Display/add61/c26 ;
  wire \u2_Display/add61/c27 ;
  wire \u2_Display/add61/c28 ;
  wire \u2_Display/add61/c29 ;
  wire \u2_Display/add61/c3 ;
  wire \u2_Display/add61/c30 ;
  wire \u2_Display/add61/c31 ;
  wire \u2_Display/add61/c4 ;
  wire \u2_Display/add61/c5 ;
  wire \u2_Display/add61/c6 ;
  wire \u2_Display/add61/c7 ;
  wire \u2_Display/add61/c8 ;
  wire \u2_Display/add61/c9 ;
  wire \u2_Display/add62/c0 ;
  wire \u2_Display/add62/c1 ;
  wire \u2_Display/add62/c10 ;
  wire \u2_Display/add62/c11 ;
  wire \u2_Display/add62/c12 ;
  wire \u2_Display/add62/c13 ;
  wire \u2_Display/add62/c14 ;
  wire \u2_Display/add62/c15 ;
  wire \u2_Display/add62/c16 ;
  wire \u2_Display/add62/c17 ;
  wire \u2_Display/add62/c18 ;
  wire \u2_Display/add62/c19 ;
  wire \u2_Display/add62/c2 ;
  wire \u2_Display/add62/c20 ;
  wire \u2_Display/add62/c21 ;
  wire \u2_Display/add62/c22 ;
  wire \u2_Display/add62/c23 ;
  wire \u2_Display/add62/c24 ;
  wire \u2_Display/add62/c25 ;
  wire \u2_Display/add62/c26 ;
  wire \u2_Display/add62/c27 ;
  wire \u2_Display/add62/c28 ;
  wire \u2_Display/add62/c29 ;
  wire \u2_Display/add62/c3 ;
  wire \u2_Display/add62/c30 ;
  wire \u2_Display/add62/c31 ;
  wire \u2_Display/add62/c4 ;
  wire \u2_Display/add62/c5 ;
  wire \u2_Display/add62/c6 ;
  wire \u2_Display/add62/c7 ;
  wire \u2_Display/add62/c8 ;
  wire \u2_Display/add62/c9 ;
  wire \u2_Display/add63/c0 ;
  wire \u2_Display/add63/c1 ;
  wire \u2_Display/add63/c10 ;
  wire \u2_Display/add63/c11 ;
  wire \u2_Display/add63/c12 ;
  wire \u2_Display/add63/c13 ;
  wire \u2_Display/add63/c14 ;
  wire \u2_Display/add63/c15 ;
  wire \u2_Display/add63/c16 ;
  wire \u2_Display/add63/c17 ;
  wire \u2_Display/add63/c18 ;
  wire \u2_Display/add63/c19 ;
  wire \u2_Display/add63/c2 ;
  wire \u2_Display/add63/c20 ;
  wire \u2_Display/add63/c21 ;
  wire \u2_Display/add63/c22 ;
  wire \u2_Display/add63/c23 ;
  wire \u2_Display/add63/c24 ;
  wire \u2_Display/add63/c25 ;
  wire \u2_Display/add63/c26 ;
  wire \u2_Display/add63/c27 ;
  wire \u2_Display/add63/c28 ;
  wire \u2_Display/add63/c29 ;
  wire \u2_Display/add63/c3 ;
  wire \u2_Display/add63/c30 ;
  wire \u2_Display/add63/c31 ;
  wire \u2_Display/add63/c4 ;
  wire \u2_Display/add63/c5 ;
  wire \u2_Display/add63/c6 ;
  wire \u2_Display/add63/c7 ;
  wire \u2_Display/add63/c8 ;
  wire \u2_Display/add63/c9 ;
  wire \u2_Display/add64/c0 ;
  wire \u2_Display/add64/c1 ;
  wire \u2_Display/add64/c10 ;
  wire \u2_Display/add64/c11 ;
  wire \u2_Display/add64/c12 ;
  wire \u2_Display/add64/c13 ;
  wire \u2_Display/add64/c14 ;
  wire \u2_Display/add64/c15 ;
  wire \u2_Display/add64/c16 ;
  wire \u2_Display/add64/c17 ;
  wire \u2_Display/add64/c18 ;
  wire \u2_Display/add64/c19 ;
  wire \u2_Display/add64/c2 ;
  wire \u2_Display/add64/c20 ;
  wire \u2_Display/add64/c21 ;
  wire \u2_Display/add64/c22 ;
  wire \u2_Display/add64/c23 ;
  wire \u2_Display/add64/c24 ;
  wire \u2_Display/add64/c25 ;
  wire \u2_Display/add64/c26 ;
  wire \u2_Display/add64/c27 ;
  wire \u2_Display/add64/c28 ;
  wire \u2_Display/add64/c29 ;
  wire \u2_Display/add64/c3 ;
  wire \u2_Display/add64/c30 ;
  wire \u2_Display/add64/c31 ;
  wire \u2_Display/add64/c4 ;
  wire \u2_Display/add64/c5 ;
  wire \u2_Display/add64/c6 ;
  wire \u2_Display/add64/c7 ;
  wire \u2_Display/add64/c8 ;
  wire \u2_Display/add64/c9 ;
  wire \u2_Display/add65/c0 ;
  wire \u2_Display/add65/c1 ;
  wire \u2_Display/add65/c10 ;
  wire \u2_Display/add65/c11 ;
  wire \u2_Display/add65/c12 ;
  wire \u2_Display/add65/c13 ;
  wire \u2_Display/add65/c14 ;
  wire \u2_Display/add65/c15 ;
  wire \u2_Display/add65/c16 ;
  wire \u2_Display/add65/c17 ;
  wire \u2_Display/add65/c18 ;
  wire \u2_Display/add65/c19 ;
  wire \u2_Display/add65/c2 ;
  wire \u2_Display/add65/c20 ;
  wire \u2_Display/add65/c21 ;
  wire \u2_Display/add65/c22 ;
  wire \u2_Display/add65/c23 ;
  wire \u2_Display/add65/c24 ;
  wire \u2_Display/add65/c25 ;
  wire \u2_Display/add65/c26 ;
  wire \u2_Display/add65/c27 ;
  wire \u2_Display/add65/c28 ;
  wire \u2_Display/add65/c29 ;
  wire \u2_Display/add65/c3 ;
  wire \u2_Display/add65/c30 ;
  wire \u2_Display/add65/c31 ;
  wire \u2_Display/add65/c4 ;
  wire \u2_Display/add65/c5 ;
  wire \u2_Display/add65/c6 ;
  wire \u2_Display/add65/c7 ;
  wire \u2_Display/add65/c8 ;
  wire \u2_Display/add65/c9 ;
  wire \u2_Display/add66/c0 ;
  wire \u2_Display/add66/c1 ;
  wire \u2_Display/add66/c10 ;
  wire \u2_Display/add66/c11 ;
  wire \u2_Display/add66/c12 ;
  wire \u2_Display/add66/c13 ;
  wire \u2_Display/add66/c14 ;
  wire \u2_Display/add66/c15 ;
  wire \u2_Display/add66/c16 ;
  wire \u2_Display/add66/c17 ;
  wire \u2_Display/add66/c18 ;
  wire \u2_Display/add66/c19 ;
  wire \u2_Display/add66/c2 ;
  wire \u2_Display/add66/c20 ;
  wire \u2_Display/add66/c21 ;
  wire \u2_Display/add66/c22 ;
  wire \u2_Display/add66/c23 ;
  wire \u2_Display/add66/c24 ;
  wire \u2_Display/add66/c25 ;
  wire \u2_Display/add66/c26 ;
  wire \u2_Display/add66/c27 ;
  wire \u2_Display/add66/c28 ;
  wire \u2_Display/add66/c29 ;
  wire \u2_Display/add66/c3 ;
  wire \u2_Display/add66/c30 ;
  wire \u2_Display/add66/c31 ;
  wire \u2_Display/add66/c4 ;
  wire \u2_Display/add66/c5 ;
  wire \u2_Display/add66/c6 ;
  wire \u2_Display/add66/c7 ;
  wire \u2_Display/add66/c8 ;
  wire \u2_Display/add66/c9 ;
  wire \u2_Display/add67/c0 ;
  wire \u2_Display/add67/c1 ;
  wire \u2_Display/add67/c10 ;
  wire \u2_Display/add67/c11 ;
  wire \u2_Display/add67/c12 ;
  wire \u2_Display/add67/c13 ;
  wire \u2_Display/add67/c14 ;
  wire \u2_Display/add67/c15 ;
  wire \u2_Display/add67/c16 ;
  wire \u2_Display/add67/c17 ;
  wire \u2_Display/add67/c18 ;
  wire \u2_Display/add67/c19 ;
  wire \u2_Display/add67/c2 ;
  wire \u2_Display/add67/c20 ;
  wire \u2_Display/add67/c21 ;
  wire \u2_Display/add67/c22 ;
  wire \u2_Display/add67/c23 ;
  wire \u2_Display/add67/c24 ;
  wire \u2_Display/add67/c25 ;
  wire \u2_Display/add67/c26 ;
  wire \u2_Display/add67/c27 ;
  wire \u2_Display/add67/c28 ;
  wire \u2_Display/add67/c29 ;
  wire \u2_Display/add67/c3 ;
  wire \u2_Display/add67/c30 ;
  wire \u2_Display/add67/c31 ;
  wire \u2_Display/add67/c4 ;
  wire \u2_Display/add67/c5 ;
  wire \u2_Display/add67/c6 ;
  wire \u2_Display/add67/c7 ;
  wire \u2_Display/add67/c8 ;
  wire \u2_Display/add67/c9 ;
  wire \u2_Display/add68/c0 ;
  wire \u2_Display/add68/c1 ;
  wire \u2_Display/add68/c10 ;
  wire \u2_Display/add68/c11 ;
  wire \u2_Display/add68/c12 ;
  wire \u2_Display/add68/c13 ;
  wire \u2_Display/add68/c14 ;
  wire \u2_Display/add68/c15 ;
  wire \u2_Display/add68/c16 ;
  wire \u2_Display/add68/c17 ;
  wire \u2_Display/add68/c18 ;
  wire \u2_Display/add68/c19 ;
  wire \u2_Display/add68/c2 ;
  wire \u2_Display/add68/c20 ;
  wire \u2_Display/add68/c21 ;
  wire \u2_Display/add68/c22 ;
  wire \u2_Display/add68/c23 ;
  wire \u2_Display/add68/c24 ;
  wire \u2_Display/add68/c25 ;
  wire \u2_Display/add68/c26 ;
  wire \u2_Display/add68/c27 ;
  wire \u2_Display/add68/c28 ;
  wire \u2_Display/add68/c29 ;
  wire \u2_Display/add68/c3 ;
  wire \u2_Display/add68/c30 ;
  wire \u2_Display/add68/c31 ;
  wire \u2_Display/add68/c4 ;
  wire \u2_Display/add68/c5 ;
  wire \u2_Display/add68/c6 ;
  wire \u2_Display/add68/c7 ;
  wire \u2_Display/add68/c8 ;
  wire \u2_Display/add68/c9 ;
  wire \u2_Display/add69/c0 ;
  wire \u2_Display/add69/c1 ;
  wire \u2_Display/add69/c10 ;
  wire \u2_Display/add69/c11 ;
  wire \u2_Display/add69/c12 ;
  wire \u2_Display/add69/c13 ;
  wire \u2_Display/add69/c14 ;
  wire \u2_Display/add69/c15 ;
  wire \u2_Display/add69/c16 ;
  wire \u2_Display/add69/c17 ;
  wire \u2_Display/add69/c18 ;
  wire \u2_Display/add69/c19 ;
  wire \u2_Display/add69/c2 ;
  wire \u2_Display/add69/c20 ;
  wire \u2_Display/add69/c21 ;
  wire \u2_Display/add69/c22 ;
  wire \u2_Display/add69/c23 ;
  wire \u2_Display/add69/c24 ;
  wire \u2_Display/add69/c25 ;
  wire \u2_Display/add69/c26 ;
  wire \u2_Display/add69/c27 ;
  wire \u2_Display/add69/c28 ;
  wire \u2_Display/add69/c29 ;
  wire \u2_Display/add69/c3 ;
  wire \u2_Display/add69/c30 ;
  wire \u2_Display/add69/c31 ;
  wire \u2_Display/add69/c4 ;
  wire \u2_Display/add69/c5 ;
  wire \u2_Display/add69/c6 ;
  wire \u2_Display/add69/c7 ;
  wire \u2_Display/add69/c8 ;
  wire \u2_Display/add69/c9 ;
  wire \u2_Display/add6_2/c0 ;
  wire \u2_Display/add6_2/c1 ;
  wire \u2_Display/add6_2/c2 ;
  wire \u2_Display/add6_2/c3 ;
  wire \u2_Display/add6_2_co ;
  wire \u2_Display/add70/c0 ;
  wire \u2_Display/add70/c1 ;
  wire \u2_Display/add70/c10 ;
  wire \u2_Display/add70/c11 ;
  wire \u2_Display/add70/c12 ;
  wire \u2_Display/add70/c13 ;
  wire \u2_Display/add70/c14 ;
  wire \u2_Display/add70/c15 ;
  wire \u2_Display/add70/c16 ;
  wire \u2_Display/add70/c17 ;
  wire \u2_Display/add70/c18 ;
  wire \u2_Display/add70/c19 ;
  wire \u2_Display/add70/c2 ;
  wire \u2_Display/add70/c20 ;
  wire \u2_Display/add70/c21 ;
  wire \u2_Display/add70/c22 ;
  wire \u2_Display/add70/c23 ;
  wire \u2_Display/add70/c24 ;
  wire \u2_Display/add70/c25 ;
  wire \u2_Display/add70/c26 ;
  wire \u2_Display/add70/c27 ;
  wire \u2_Display/add70/c28 ;
  wire \u2_Display/add70/c29 ;
  wire \u2_Display/add70/c3 ;
  wire \u2_Display/add70/c30 ;
  wire \u2_Display/add70/c31 ;
  wire \u2_Display/add70/c4 ;
  wire \u2_Display/add70/c5 ;
  wire \u2_Display/add70/c6 ;
  wire \u2_Display/add70/c7 ;
  wire \u2_Display/add70/c8 ;
  wire \u2_Display/add70/c9 ;
  wire \u2_Display/add71/c0 ;
  wire \u2_Display/add71/c1 ;
  wire \u2_Display/add71/c10 ;
  wire \u2_Display/add71/c11 ;
  wire \u2_Display/add71/c12 ;
  wire \u2_Display/add71/c13 ;
  wire \u2_Display/add71/c14 ;
  wire \u2_Display/add71/c15 ;
  wire \u2_Display/add71/c16 ;
  wire \u2_Display/add71/c17 ;
  wire \u2_Display/add71/c18 ;
  wire \u2_Display/add71/c19 ;
  wire \u2_Display/add71/c2 ;
  wire \u2_Display/add71/c20 ;
  wire \u2_Display/add71/c21 ;
  wire \u2_Display/add71/c22 ;
  wire \u2_Display/add71/c23 ;
  wire \u2_Display/add71/c24 ;
  wire \u2_Display/add71/c25 ;
  wire \u2_Display/add71/c26 ;
  wire \u2_Display/add71/c27 ;
  wire \u2_Display/add71/c28 ;
  wire \u2_Display/add71/c29 ;
  wire \u2_Display/add71/c3 ;
  wire \u2_Display/add71/c30 ;
  wire \u2_Display/add71/c31 ;
  wire \u2_Display/add71/c4 ;
  wire \u2_Display/add71/c5 ;
  wire \u2_Display/add71/c6 ;
  wire \u2_Display/add71/c7 ;
  wire \u2_Display/add71/c8 ;
  wire \u2_Display/add71/c9 ;
  wire \u2_Display/add72/c0 ;
  wire \u2_Display/add72/c1 ;
  wire \u2_Display/add72/c10 ;
  wire \u2_Display/add72/c11 ;
  wire \u2_Display/add72/c12 ;
  wire \u2_Display/add72/c13 ;
  wire \u2_Display/add72/c14 ;
  wire \u2_Display/add72/c15 ;
  wire \u2_Display/add72/c16 ;
  wire \u2_Display/add72/c17 ;
  wire \u2_Display/add72/c18 ;
  wire \u2_Display/add72/c19 ;
  wire \u2_Display/add72/c2 ;
  wire \u2_Display/add72/c20 ;
  wire \u2_Display/add72/c21 ;
  wire \u2_Display/add72/c22 ;
  wire \u2_Display/add72/c23 ;
  wire \u2_Display/add72/c24 ;
  wire \u2_Display/add72/c25 ;
  wire \u2_Display/add72/c26 ;
  wire \u2_Display/add72/c27 ;
  wire \u2_Display/add72/c28 ;
  wire \u2_Display/add72/c29 ;
  wire \u2_Display/add72/c3 ;
  wire \u2_Display/add72/c30 ;
  wire \u2_Display/add72/c31 ;
  wire \u2_Display/add72/c4 ;
  wire \u2_Display/add72/c5 ;
  wire \u2_Display/add72/c6 ;
  wire \u2_Display/add72/c7 ;
  wire \u2_Display/add72/c8 ;
  wire \u2_Display/add72/c9 ;
  wire \u2_Display/add73/c0 ;
  wire \u2_Display/add73/c1 ;
  wire \u2_Display/add73/c2 ;
  wire \u2_Display/add73/c3 ;
  wire \u2_Display/add73/c4 ;
  wire \u2_Display/add73/c5 ;
  wire \u2_Display/add73/c6 ;
  wire \u2_Display/add73/c7 ;
  wire \u2_Display/add73/c8 ;
  wire \u2_Display/add73/c9 ;
  wire \u2_Display/add7_2_co ;
  wire \u2_Display/add84/c0 ;
  wire \u2_Display/add84/c1 ;
  wire \u2_Display/add84/c10 ;
  wire \u2_Display/add84/c11 ;
  wire \u2_Display/add84/c12 ;
  wire \u2_Display/add84/c13 ;
  wire \u2_Display/add84/c14 ;
  wire \u2_Display/add84/c15 ;
  wire \u2_Display/add84/c16 ;
  wire \u2_Display/add84/c17 ;
  wire \u2_Display/add84/c18 ;
  wire \u2_Display/add84/c19 ;
  wire \u2_Display/add84/c2 ;
  wire \u2_Display/add84/c20 ;
  wire \u2_Display/add84/c21 ;
  wire \u2_Display/add84/c22 ;
  wire \u2_Display/add84/c23 ;
  wire \u2_Display/add84/c24 ;
  wire \u2_Display/add84/c25 ;
  wire \u2_Display/add84/c26 ;
  wire \u2_Display/add84/c27 ;
  wire \u2_Display/add84/c28 ;
  wire \u2_Display/add84/c29 ;
  wire \u2_Display/add84/c3 ;
  wire \u2_Display/add84/c30 ;
  wire \u2_Display/add84/c31 ;
  wire \u2_Display/add84/c4 ;
  wire \u2_Display/add84/c5 ;
  wire \u2_Display/add84/c6 ;
  wire \u2_Display/add84/c7 ;
  wire \u2_Display/add84/c8 ;
  wire \u2_Display/add84/c9 ;
  wire \u2_Display/add85/c0 ;
  wire \u2_Display/add85/c1 ;
  wire \u2_Display/add85/c10 ;
  wire \u2_Display/add85/c11 ;
  wire \u2_Display/add85/c12 ;
  wire \u2_Display/add85/c13 ;
  wire \u2_Display/add85/c14 ;
  wire \u2_Display/add85/c15 ;
  wire \u2_Display/add85/c16 ;
  wire \u2_Display/add85/c17 ;
  wire \u2_Display/add85/c18 ;
  wire \u2_Display/add85/c19 ;
  wire \u2_Display/add85/c2 ;
  wire \u2_Display/add85/c20 ;
  wire \u2_Display/add85/c21 ;
  wire \u2_Display/add85/c22 ;
  wire \u2_Display/add85/c23 ;
  wire \u2_Display/add85/c24 ;
  wire \u2_Display/add85/c25 ;
  wire \u2_Display/add85/c26 ;
  wire \u2_Display/add85/c27 ;
  wire \u2_Display/add85/c28 ;
  wire \u2_Display/add85/c29 ;
  wire \u2_Display/add85/c3 ;
  wire \u2_Display/add85/c30 ;
  wire \u2_Display/add85/c31 ;
  wire \u2_Display/add85/c4 ;
  wire \u2_Display/add85/c5 ;
  wire \u2_Display/add85/c6 ;
  wire \u2_Display/add85/c7 ;
  wire \u2_Display/add85/c8 ;
  wire \u2_Display/add85/c9 ;
  wire \u2_Display/add86/c0 ;
  wire \u2_Display/add86/c1 ;
  wire \u2_Display/add86/c10 ;
  wire \u2_Display/add86/c11 ;
  wire \u2_Display/add86/c12 ;
  wire \u2_Display/add86/c13 ;
  wire \u2_Display/add86/c14 ;
  wire \u2_Display/add86/c15 ;
  wire \u2_Display/add86/c16 ;
  wire \u2_Display/add86/c17 ;
  wire \u2_Display/add86/c18 ;
  wire \u2_Display/add86/c19 ;
  wire \u2_Display/add86/c2 ;
  wire \u2_Display/add86/c20 ;
  wire \u2_Display/add86/c21 ;
  wire \u2_Display/add86/c22 ;
  wire \u2_Display/add86/c23 ;
  wire \u2_Display/add86/c24 ;
  wire \u2_Display/add86/c25 ;
  wire \u2_Display/add86/c26 ;
  wire \u2_Display/add86/c27 ;
  wire \u2_Display/add86/c28 ;
  wire \u2_Display/add86/c29 ;
  wire \u2_Display/add86/c3 ;
  wire \u2_Display/add86/c30 ;
  wire \u2_Display/add86/c31 ;
  wire \u2_Display/add86/c4 ;
  wire \u2_Display/add86/c5 ;
  wire \u2_Display/add86/c6 ;
  wire \u2_Display/add86/c7 ;
  wire \u2_Display/add86/c8 ;
  wire \u2_Display/add86/c9 ;
  wire \u2_Display/add87/c0 ;
  wire \u2_Display/add87/c1 ;
  wire \u2_Display/add87/c10 ;
  wire \u2_Display/add87/c11 ;
  wire \u2_Display/add87/c12 ;
  wire \u2_Display/add87/c13 ;
  wire \u2_Display/add87/c14 ;
  wire \u2_Display/add87/c15 ;
  wire \u2_Display/add87/c16 ;
  wire \u2_Display/add87/c17 ;
  wire \u2_Display/add87/c18 ;
  wire \u2_Display/add87/c19 ;
  wire \u2_Display/add87/c2 ;
  wire \u2_Display/add87/c20 ;
  wire \u2_Display/add87/c21 ;
  wire \u2_Display/add87/c22 ;
  wire \u2_Display/add87/c23 ;
  wire \u2_Display/add87/c24 ;
  wire \u2_Display/add87/c25 ;
  wire \u2_Display/add87/c26 ;
  wire \u2_Display/add87/c27 ;
  wire \u2_Display/add87/c28 ;
  wire \u2_Display/add87/c29 ;
  wire \u2_Display/add87/c3 ;
  wire \u2_Display/add87/c30 ;
  wire \u2_Display/add87/c31 ;
  wire \u2_Display/add87/c4 ;
  wire \u2_Display/add87/c5 ;
  wire \u2_Display/add87/c6 ;
  wire \u2_Display/add87/c7 ;
  wire \u2_Display/add87/c8 ;
  wire \u2_Display/add87/c9 ;
  wire \u2_Display/add88/c0 ;
  wire \u2_Display/add88/c1 ;
  wire \u2_Display/add88/c10 ;
  wire \u2_Display/add88/c11 ;
  wire \u2_Display/add88/c12 ;
  wire \u2_Display/add88/c13 ;
  wire \u2_Display/add88/c14 ;
  wire \u2_Display/add88/c15 ;
  wire \u2_Display/add88/c16 ;
  wire \u2_Display/add88/c17 ;
  wire \u2_Display/add88/c18 ;
  wire \u2_Display/add88/c19 ;
  wire \u2_Display/add88/c2 ;
  wire \u2_Display/add88/c20 ;
  wire \u2_Display/add88/c21 ;
  wire \u2_Display/add88/c22 ;
  wire \u2_Display/add88/c23 ;
  wire \u2_Display/add88/c24 ;
  wire \u2_Display/add88/c25 ;
  wire \u2_Display/add88/c26 ;
  wire \u2_Display/add88/c27 ;
  wire \u2_Display/add88/c28 ;
  wire \u2_Display/add88/c29 ;
  wire \u2_Display/add88/c3 ;
  wire \u2_Display/add88/c30 ;
  wire \u2_Display/add88/c31 ;
  wire \u2_Display/add88/c4 ;
  wire \u2_Display/add88/c5 ;
  wire \u2_Display/add88/c6 ;
  wire \u2_Display/add88/c7 ;
  wire \u2_Display/add88/c8 ;
  wire \u2_Display/add88/c9 ;
  wire \u2_Display/add89/c0 ;
  wire \u2_Display/add89/c1 ;
  wire \u2_Display/add89/c10 ;
  wire \u2_Display/add89/c11 ;
  wire \u2_Display/add89/c12 ;
  wire \u2_Display/add89/c13 ;
  wire \u2_Display/add89/c14 ;
  wire \u2_Display/add89/c15 ;
  wire \u2_Display/add89/c16 ;
  wire \u2_Display/add89/c17 ;
  wire \u2_Display/add89/c18 ;
  wire \u2_Display/add89/c19 ;
  wire \u2_Display/add89/c2 ;
  wire \u2_Display/add89/c20 ;
  wire \u2_Display/add89/c21 ;
  wire \u2_Display/add89/c22 ;
  wire \u2_Display/add89/c23 ;
  wire \u2_Display/add89/c24 ;
  wire \u2_Display/add89/c25 ;
  wire \u2_Display/add89/c26 ;
  wire \u2_Display/add89/c27 ;
  wire \u2_Display/add89/c28 ;
  wire \u2_Display/add89/c29 ;
  wire \u2_Display/add89/c3 ;
  wire \u2_Display/add89/c30 ;
  wire \u2_Display/add89/c31 ;
  wire \u2_Display/add89/c4 ;
  wire \u2_Display/add89/c5 ;
  wire \u2_Display/add89/c6 ;
  wire \u2_Display/add89/c7 ;
  wire \u2_Display/add89/c8 ;
  wire \u2_Display/add89/c9 ;
  wire \u2_Display/add90/c0 ;
  wire \u2_Display/add90/c1 ;
  wire \u2_Display/add90/c10 ;
  wire \u2_Display/add90/c11 ;
  wire \u2_Display/add90/c12 ;
  wire \u2_Display/add90/c13 ;
  wire \u2_Display/add90/c14 ;
  wire \u2_Display/add90/c15 ;
  wire \u2_Display/add90/c16 ;
  wire \u2_Display/add90/c17 ;
  wire \u2_Display/add90/c18 ;
  wire \u2_Display/add90/c19 ;
  wire \u2_Display/add90/c2 ;
  wire \u2_Display/add90/c20 ;
  wire \u2_Display/add90/c21 ;
  wire \u2_Display/add90/c22 ;
  wire \u2_Display/add90/c23 ;
  wire \u2_Display/add90/c24 ;
  wire \u2_Display/add90/c25 ;
  wire \u2_Display/add90/c26 ;
  wire \u2_Display/add90/c27 ;
  wire \u2_Display/add90/c28 ;
  wire \u2_Display/add90/c29 ;
  wire \u2_Display/add90/c3 ;
  wire \u2_Display/add90/c30 ;
  wire \u2_Display/add90/c31 ;
  wire \u2_Display/add90/c4 ;
  wire \u2_Display/add90/c5 ;
  wire \u2_Display/add90/c6 ;
  wire \u2_Display/add90/c7 ;
  wire \u2_Display/add90/c8 ;
  wire \u2_Display/add90/c9 ;
  wire \u2_Display/add91/c0 ;
  wire \u2_Display/add91/c1 ;
  wire \u2_Display/add91/c10 ;
  wire \u2_Display/add91/c11 ;
  wire \u2_Display/add91/c12 ;
  wire \u2_Display/add91/c13 ;
  wire \u2_Display/add91/c14 ;
  wire \u2_Display/add91/c15 ;
  wire \u2_Display/add91/c16 ;
  wire \u2_Display/add91/c17 ;
  wire \u2_Display/add91/c18 ;
  wire \u2_Display/add91/c19 ;
  wire \u2_Display/add91/c2 ;
  wire \u2_Display/add91/c20 ;
  wire \u2_Display/add91/c21 ;
  wire \u2_Display/add91/c22 ;
  wire \u2_Display/add91/c23 ;
  wire \u2_Display/add91/c24 ;
  wire \u2_Display/add91/c25 ;
  wire \u2_Display/add91/c26 ;
  wire \u2_Display/add91/c27 ;
  wire \u2_Display/add91/c28 ;
  wire \u2_Display/add91/c29 ;
  wire \u2_Display/add91/c3 ;
  wire \u2_Display/add91/c30 ;
  wire \u2_Display/add91/c31 ;
  wire \u2_Display/add91/c4 ;
  wire \u2_Display/add91/c5 ;
  wire \u2_Display/add91/c6 ;
  wire \u2_Display/add91/c7 ;
  wire \u2_Display/add91/c8 ;
  wire \u2_Display/add91/c9 ;
  wire \u2_Display/add92/c0 ;
  wire \u2_Display/add92/c1 ;
  wire \u2_Display/add92/c10 ;
  wire \u2_Display/add92/c11 ;
  wire \u2_Display/add92/c12 ;
  wire \u2_Display/add92/c13 ;
  wire \u2_Display/add92/c14 ;
  wire \u2_Display/add92/c15 ;
  wire \u2_Display/add92/c16 ;
  wire \u2_Display/add92/c17 ;
  wire \u2_Display/add92/c18 ;
  wire \u2_Display/add92/c19 ;
  wire \u2_Display/add92/c2 ;
  wire \u2_Display/add92/c20 ;
  wire \u2_Display/add92/c21 ;
  wire \u2_Display/add92/c22 ;
  wire \u2_Display/add92/c23 ;
  wire \u2_Display/add92/c24 ;
  wire \u2_Display/add92/c25 ;
  wire \u2_Display/add92/c26 ;
  wire \u2_Display/add92/c27 ;
  wire \u2_Display/add92/c28 ;
  wire \u2_Display/add92/c29 ;
  wire \u2_Display/add92/c3 ;
  wire \u2_Display/add92/c30 ;
  wire \u2_Display/add92/c31 ;
  wire \u2_Display/add92/c4 ;
  wire \u2_Display/add92/c5 ;
  wire \u2_Display/add92/c6 ;
  wire \u2_Display/add92/c7 ;
  wire \u2_Display/add92/c8 ;
  wire \u2_Display/add92/c9 ;
  wire \u2_Display/add93/c0 ;
  wire \u2_Display/add93/c1 ;
  wire \u2_Display/add93/c10 ;
  wire \u2_Display/add93/c11 ;
  wire \u2_Display/add93/c12 ;
  wire \u2_Display/add93/c13 ;
  wire \u2_Display/add93/c14 ;
  wire \u2_Display/add93/c15 ;
  wire \u2_Display/add93/c16 ;
  wire \u2_Display/add93/c17 ;
  wire \u2_Display/add93/c18 ;
  wire \u2_Display/add93/c19 ;
  wire \u2_Display/add93/c2 ;
  wire \u2_Display/add93/c20 ;
  wire \u2_Display/add93/c21 ;
  wire \u2_Display/add93/c22 ;
  wire \u2_Display/add93/c23 ;
  wire \u2_Display/add93/c24 ;
  wire \u2_Display/add93/c25 ;
  wire \u2_Display/add93/c26 ;
  wire \u2_Display/add93/c27 ;
  wire \u2_Display/add93/c28 ;
  wire \u2_Display/add93/c29 ;
  wire \u2_Display/add93/c3 ;
  wire \u2_Display/add93/c30 ;
  wire \u2_Display/add93/c31 ;
  wire \u2_Display/add93/c4 ;
  wire \u2_Display/add93/c5 ;
  wire \u2_Display/add93/c6 ;
  wire \u2_Display/add93/c7 ;
  wire \u2_Display/add93/c8 ;
  wire \u2_Display/add93/c9 ;
  wire \u2_Display/add94/c0 ;
  wire \u2_Display/add94/c1 ;
  wire \u2_Display/add94/c10 ;
  wire \u2_Display/add94/c11 ;
  wire \u2_Display/add94/c12 ;
  wire \u2_Display/add94/c13 ;
  wire \u2_Display/add94/c14 ;
  wire \u2_Display/add94/c15 ;
  wire \u2_Display/add94/c16 ;
  wire \u2_Display/add94/c17 ;
  wire \u2_Display/add94/c18 ;
  wire \u2_Display/add94/c19 ;
  wire \u2_Display/add94/c2 ;
  wire \u2_Display/add94/c20 ;
  wire \u2_Display/add94/c21 ;
  wire \u2_Display/add94/c22 ;
  wire \u2_Display/add94/c23 ;
  wire \u2_Display/add94/c24 ;
  wire \u2_Display/add94/c25 ;
  wire \u2_Display/add94/c26 ;
  wire \u2_Display/add94/c27 ;
  wire \u2_Display/add94/c28 ;
  wire \u2_Display/add94/c29 ;
  wire \u2_Display/add94/c3 ;
  wire \u2_Display/add94/c30 ;
  wire \u2_Display/add94/c31 ;
  wire \u2_Display/add94/c4 ;
  wire \u2_Display/add94/c5 ;
  wire \u2_Display/add94/c6 ;
  wire \u2_Display/add94/c7 ;
  wire \u2_Display/add94/c8 ;
  wire \u2_Display/add94/c9 ;
  wire \u2_Display/add95/c0 ;
  wire \u2_Display/add95/c1 ;
  wire \u2_Display/add95/c10 ;
  wire \u2_Display/add95/c11 ;
  wire \u2_Display/add95/c12 ;
  wire \u2_Display/add95/c13 ;
  wire \u2_Display/add95/c14 ;
  wire \u2_Display/add95/c15 ;
  wire \u2_Display/add95/c16 ;
  wire \u2_Display/add95/c17 ;
  wire \u2_Display/add95/c18 ;
  wire \u2_Display/add95/c19 ;
  wire \u2_Display/add95/c2 ;
  wire \u2_Display/add95/c20 ;
  wire \u2_Display/add95/c21 ;
  wire \u2_Display/add95/c22 ;
  wire \u2_Display/add95/c23 ;
  wire \u2_Display/add95/c24 ;
  wire \u2_Display/add95/c25 ;
  wire \u2_Display/add95/c26 ;
  wire \u2_Display/add95/c27 ;
  wire \u2_Display/add95/c28 ;
  wire \u2_Display/add95/c29 ;
  wire \u2_Display/add95/c3 ;
  wire \u2_Display/add95/c30 ;
  wire \u2_Display/add95/c31 ;
  wire \u2_Display/add95/c4 ;
  wire \u2_Display/add95/c5 ;
  wire \u2_Display/add95/c6 ;
  wire \u2_Display/add95/c7 ;
  wire \u2_Display/add95/c8 ;
  wire \u2_Display/add95/c9 ;
  wire \u2_Display/add96/c0 ;
  wire \u2_Display/add96/c1 ;
  wire \u2_Display/add96/c10 ;
  wire \u2_Display/add96/c11 ;
  wire \u2_Display/add96/c12 ;
  wire \u2_Display/add96/c13 ;
  wire \u2_Display/add96/c14 ;
  wire \u2_Display/add96/c15 ;
  wire \u2_Display/add96/c16 ;
  wire \u2_Display/add96/c17 ;
  wire \u2_Display/add96/c18 ;
  wire \u2_Display/add96/c19 ;
  wire \u2_Display/add96/c2 ;
  wire \u2_Display/add96/c20 ;
  wire \u2_Display/add96/c21 ;
  wire \u2_Display/add96/c22 ;
  wire \u2_Display/add96/c23 ;
  wire \u2_Display/add96/c24 ;
  wire \u2_Display/add96/c25 ;
  wire \u2_Display/add96/c26 ;
  wire \u2_Display/add96/c27 ;
  wire \u2_Display/add96/c28 ;
  wire \u2_Display/add96/c29 ;
  wire \u2_Display/add96/c3 ;
  wire \u2_Display/add96/c30 ;
  wire \u2_Display/add96/c31 ;
  wire \u2_Display/add96/c4 ;
  wire \u2_Display/add96/c5 ;
  wire \u2_Display/add96/c6 ;
  wire \u2_Display/add96/c7 ;
  wire \u2_Display/add96/c8 ;
  wire \u2_Display/add96/c9 ;
  wire \u2_Display/add97/c0 ;
  wire \u2_Display/add97/c1 ;
  wire \u2_Display/add97/c10 ;
  wire \u2_Display/add97/c11 ;
  wire \u2_Display/add97/c12 ;
  wire \u2_Display/add97/c13 ;
  wire \u2_Display/add97/c14 ;
  wire \u2_Display/add97/c15 ;
  wire \u2_Display/add97/c16 ;
  wire \u2_Display/add97/c17 ;
  wire \u2_Display/add97/c18 ;
  wire \u2_Display/add97/c19 ;
  wire \u2_Display/add97/c2 ;
  wire \u2_Display/add97/c20 ;
  wire \u2_Display/add97/c21 ;
  wire \u2_Display/add97/c22 ;
  wire \u2_Display/add97/c23 ;
  wire \u2_Display/add97/c24 ;
  wire \u2_Display/add97/c25 ;
  wire \u2_Display/add97/c26 ;
  wire \u2_Display/add97/c27 ;
  wire \u2_Display/add97/c28 ;
  wire \u2_Display/add97/c29 ;
  wire \u2_Display/add97/c3 ;
  wire \u2_Display/add97/c30 ;
  wire \u2_Display/add97/c31 ;
  wire \u2_Display/add97/c4 ;
  wire \u2_Display/add97/c5 ;
  wire \u2_Display/add97/c6 ;
  wire \u2_Display/add97/c7 ;
  wire \u2_Display/add97/c8 ;
  wire \u2_Display/add97/c9 ;
  wire \u2_Display/add98/c0 ;
  wire \u2_Display/add98/c1 ;
  wire \u2_Display/add98/c10 ;
  wire \u2_Display/add98/c11 ;
  wire \u2_Display/add98/c12 ;
  wire \u2_Display/add98/c13 ;
  wire \u2_Display/add98/c14 ;
  wire \u2_Display/add98/c15 ;
  wire \u2_Display/add98/c16 ;
  wire \u2_Display/add98/c17 ;
  wire \u2_Display/add98/c18 ;
  wire \u2_Display/add98/c19 ;
  wire \u2_Display/add98/c2 ;
  wire \u2_Display/add98/c20 ;
  wire \u2_Display/add98/c21 ;
  wire \u2_Display/add98/c22 ;
  wire \u2_Display/add98/c23 ;
  wire \u2_Display/add98/c24 ;
  wire \u2_Display/add98/c25 ;
  wire \u2_Display/add98/c26 ;
  wire \u2_Display/add98/c27 ;
  wire \u2_Display/add98/c28 ;
  wire \u2_Display/add98/c29 ;
  wire \u2_Display/add98/c3 ;
  wire \u2_Display/add98/c30 ;
  wire \u2_Display/add98/c31 ;
  wire \u2_Display/add98/c4 ;
  wire \u2_Display/add98/c5 ;
  wire \u2_Display/add98/c6 ;
  wire \u2_Display/add98/c7 ;
  wire \u2_Display/add98/c8 ;
  wire \u2_Display/add98/c9 ;
  wire \u2_Display/add99/c0 ;
  wire \u2_Display/add99/c1 ;
  wire \u2_Display/add99/c10 ;
  wire \u2_Display/add99/c11 ;
  wire \u2_Display/add99/c12 ;
  wire \u2_Display/add99/c13 ;
  wire \u2_Display/add99/c14 ;
  wire \u2_Display/add99/c15 ;
  wire \u2_Display/add99/c16 ;
  wire \u2_Display/add99/c17 ;
  wire \u2_Display/add99/c18 ;
  wire \u2_Display/add99/c19 ;
  wire \u2_Display/add99/c2 ;
  wire \u2_Display/add99/c20 ;
  wire \u2_Display/add99/c21 ;
  wire \u2_Display/add99/c22 ;
  wire \u2_Display/add99/c23 ;
  wire \u2_Display/add99/c24 ;
  wire \u2_Display/add99/c25 ;
  wire \u2_Display/add99/c26 ;
  wire \u2_Display/add99/c27 ;
  wire \u2_Display/add99/c28 ;
  wire \u2_Display/add99/c29 ;
  wire \u2_Display/add99/c3 ;
  wire \u2_Display/add99/c30 ;
  wire \u2_Display/add99/c31 ;
  wire \u2_Display/add99/c4 ;
  wire \u2_Display/add99/c5 ;
  wire \u2_Display/add99/c6 ;
  wire \u2_Display/add99/c7 ;
  wire \u2_Display/add99/c8 ;
  wire \u2_Display/add99/c9 ;
  wire \u2_Display/clk1s ;  // source/rtl/Display.v(46)
  wire \u2_Display/lt0_2_c0 ;
  wire \u2_Display/lt0_2_c1 ;
  wire \u2_Display/lt0_2_c10 ;
  wire \u2_Display/lt0_2_c11 ;
  wire \u2_Display/lt0_2_c12 ;
  wire \u2_Display/lt0_2_c2 ;
  wire \u2_Display/lt0_2_c3 ;
  wire \u2_Display/lt0_2_c4 ;
  wire \u2_Display/lt0_2_c5 ;
  wire \u2_Display/lt0_2_c6 ;
  wire \u2_Display/lt0_2_c7 ;
  wire \u2_Display/lt0_2_c8 ;
  wire \u2_Display/lt0_2_c9 ;
  wire \u2_Display/lt100_c0 ;
  wire \u2_Display/lt100_c1 ;
  wire \u2_Display/lt100_c10 ;
  wire \u2_Display/lt100_c11 ;
  wire \u2_Display/lt100_c12 ;
  wire \u2_Display/lt100_c13 ;
  wire \u2_Display/lt100_c14 ;
  wire \u2_Display/lt100_c15 ;
  wire \u2_Display/lt100_c16 ;
  wire \u2_Display/lt100_c17 ;
  wire \u2_Display/lt100_c18 ;
  wire \u2_Display/lt100_c19 ;
  wire \u2_Display/lt100_c2 ;
  wire \u2_Display/lt100_c20 ;
  wire \u2_Display/lt100_c21 ;
  wire \u2_Display/lt100_c22 ;
  wire \u2_Display/lt100_c23 ;
  wire \u2_Display/lt100_c24 ;
  wire \u2_Display/lt100_c25 ;
  wire \u2_Display/lt100_c26 ;
  wire \u2_Display/lt100_c27 ;
  wire \u2_Display/lt100_c28 ;
  wire \u2_Display/lt100_c29 ;
  wire \u2_Display/lt100_c3 ;
  wire \u2_Display/lt100_c30 ;
  wire \u2_Display/lt100_c31 ;
  wire \u2_Display/lt100_c32 ;
  wire \u2_Display/lt100_c4 ;
  wire \u2_Display/lt100_c5 ;
  wire \u2_Display/lt100_c6 ;
  wire \u2_Display/lt100_c7 ;
  wire \u2_Display/lt100_c8 ;
  wire \u2_Display/lt100_c9 ;
  wire \u2_Display/lt101_c0 ;
  wire \u2_Display/lt101_c1 ;
  wire \u2_Display/lt101_c10 ;
  wire \u2_Display/lt101_c11 ;
  wire \u2_Display/lt101_c12 ;
  wire \u2_Display/lt101_c13 ;
  wire \u2_Display/lt101_c14 ;
  wire \u2_Display/lt101_c15 ;
  wire \u2_Display/lt101_c16 ;
  wire \u2_Display/lt101_c17 ;
  wire \u2_Display/lt101_c18 ;
  wire \u2_Display/lt101_c19 ;
  wire \u2_Display/lt101_c2 ;
  wire \u2_Display/lt101_c20 ;
  wire \u2_Display/lt101_c21 ;
  wire \u2_Display/lt101_c22 ;
  wire \u2_Display/lt101_c23 ;
  wire \u2_Display/lt101_c24 ;
  wire \u2_Display/lt101_c25 ;
  wire \u2_Display/lt101_c26 ;
  wire \u2_Display/lt101_c27 ;
  wire \u2_Display/lt101_c28 ;
  wire \u2_Display/lt101_c29 ;
  wire \u2_Display/lt101_c3 ;
  wire \u2_Display/lt101_c30 ;
  wire \u2_Display/lt101_c31 ;
  wire \u2_Display/lt101_c32 ;
  wire \u2_Display/lt101_c4 ;
  wire \u2_Display/lt101_c5 ;
  wire \u2_Display/lt101_c6 ;
  wire \u2_Display/lt101_c7 ;
  wire \u2_Display/lt101_c8 ;
  wire \u2_Display/lt101_c9 ;
  wire \u2_Display/lt102_c0 ;
  wire \u2_Display/lt102_c1 ;
  wire \u2_Display/lt102_c10 ;
  wire \u2_Display/lt102_c11 ;
  wire \u2_Display/lt102_c12 ;
  wire \u2_Display/lt102_c13 ;
  wire \u2_Display/lt102_c14 ;
  wire \u2_Display/lt102_c15 ;
  wire \u2_Display/lt102_c16 ;
  wire \u2_Display/lt102_c17 ;
  wire \u2_Display/lt102_c18 ;
  wire \u2_Display/lt102_c19 ;
  wire \u2_Display/lt102_c2 ;
  wire \u2_Display/lt102_c20 ;
  wire \u2_Display/lt102_c21 ;
  wire \u2_Display/lt102_c22 ;
  wire \u2_Display/lt102_c23 ;
  wire \u2_Display/lt102_c24 ;
  wire \u2_Display/lt102_c25 ;
  wire \u2_Display/lt102_c26 ;
  wire \u2_Display/lt102_c27 ;
  wire \u2_Display/lt102_c28 ;
  wire \u2_Display/lt102_c29 ;
  wire \u2_Display/lt102_c3 ;
  wire \u2_Display/lt102_c30 ;
  wire \u2_Display/lt102_c31 ;
  wire \u2_Display/lt102_c32 ;
  wire \u2_Display/lt102_c4 ;
  wire \u2_Display/lt102_c5 ;
  wire \u2_Display/lt102_c6 ;
  wire \u2_Display/lt102_c7 ;
  wire \u2_Display/lt102_c8 ;
  wire \u2_Display/lt102_c9 ;
  wire \u2_Display/lt103_c0 ;
  wire \u2_Display/lt103_c1 ;
  wire \u2_Display/lt103_c10 ;
  wire \u2_Display/lt103_c11 ;
  wire \u2_Display/lt103_c12 ;
  wire \u2_Display/lt103_c13 ;
  wire \u2_Display/lt103_c14 ;
  wire \u2_Display/lt103_c15 ;
  wire \u2_Display/lt103_c16 ;
  wire \u2_Display/lt103_c17 ;
  wire \u2_Display/lt103_c18 ;
  wire \u2_Display/lt103_c19 ;
  wire \u2_Display/lt103_c2 ;
  wire \u2_Display/lt103_c20 ;
  wire \u2_Display/lt103_c21 ;
  wire \u2_Display/lt103_c22 ;
  wire \u2_Display/lt103_c23 ;
  wire \u2_Display/lt103_c24 ;
  wire \u2_Display/lt103_c25 ;
  wire \u2_Display/lt103_c26 ;
  wire \u2_Display/lt103_c27 ;
  wire \u2_Display/lt103_c28 ;
  wire \u2_Display/lt103_c29 ;
  wire \u2_Display/lt103_c3 ;
  wire \u2_Display/lt103_c30 ;
  wire \u2_Display/lt103_c31 ;
  wire \u2_Display/lt103_c32 ;
  wire \u2_Display/lt103_c4 ;
  wire \u2_Display/lt103_c5 ;
  wire \u2_Display/lt103_c6 ;
  wire \u2_Display/lt103_c7 ;
  wire \u2_Display/lt103_c8 ;
  wire \u2_Display/lt103_c9 ;
  wire \u2_Display/lt104_c0 ;
  wire \u2_Display/lt104_c1 ;
  wire \u2_Display/lt104_c10 ;
  wire \u2_Display/lt104_c11 ;
  wire \u2_Display/lt104_c12 ;
  wire \u2_Display/lt104_c13 ;
  wire \u2_Display/lt104_c14 ;
  wire \u2_Display/lt104_c15 ;
  wire \u2_Display/lt104_c16 ;
  wire \u2_Display/lt104_c17 ;
  wire \u2_Display/lt104_c18 ;
  wire \u2_Display/lt104_c19 ;
  wire \u2_Display/lt104_c2 ;
  wire \u2_Display/lt104_c20 ;
  wire \u2_Display/lt104_c21 ;
  wire \u2_Display/lt104_c22 ;
  wire \u2_Display/lt104_c23 ;
  wire \u2_Display/lt104_c24 ;
  wire \u2_Display/lt104_c25 ;
  wire \u2_Display/lt104_c26 ;
  wire \u2_Display/lt104_c27 ;
  wire \u2_Display/lt104_c28 ;
  wire \u2_Display/lt104_c29 ;
  wire \u2_Display/lt104_c3 ;
  wire \u2_Display/lt104_c30 ;
  wire \u2_Display/lt104_c31 ;
  wire \u2_Display/lt104_c32 ;
  wire \u2_Display/lt104_c4 ;
  wire \u2_Display/lt104_c5 ;
  wire \u2_Display/lt104_c6 ;
  wire \u2_Display/lt104_c7 ;
  wire \u2_Display/lt104_c8 ;
  wire \u2_Display/lt104_c9 ;
  wire \u2_Display/lt105_c0 ;
  wire \u2_Display/lt105_c1 ;
  wire \u2_Display/lt105_c10 ;
  wire \u2_Display/lt105_c11 ;
  wire \u2_Display/lt105_c12 ;
  wire \u2_Display/lt105_c13 ;
  wire \u2_Display/lt105_c14 ;
  wire \u2_Display/lt105_c15 ;
  wire \u2_Display/lt105_c16 ;
  wire \u2_Display/lt105_c17 ;
  wire \u2_Display/lt105_c18 ;
  wire \u2_Display/lt105_c19 ;
  wire \u2_Display/lt105_c2 ;
  wire \u2_Display/lt105_c20 ;
  wire \u2_Display/lt105_c21 ;
  wire \u2_Display/lt105_c22 ;
  wire \u2_Display/lt105_c23 ;
  wire \u2_Display/lt105_c24 ;
  wire \u2_Display/lt105_c25 ;
  wire \u2_Display/lt105_c26 ;
  wire \u2_Display/lt105_c27 ;
  wire \u2_Display/lt105_c28 ;
  wire \u2_Display/lt105_c29 ;
  wire \u2_Display/lt105_c3 ;
  wire \u2_Display/lt105_c30 ;
  wire \u2_Display/lt105_c31 ;
  wire \u2_Display/lt105_c32 ;
  wire \u2_Display/lt105_c4 ;
  wire \u2_Display/lt105_c5 ;
  wire \u2_Display/lt105_c6 ;
  wire \u2_Display/lt105_c7 ;
  wire \u2_Display/lt105_c8 ;
  wire \u2_Display/lt105_c9 ;
  wire \u2_Display/lt106_c0 ;
  wire \u2_Display/lt106_c1 ;
  wire \u2_Display/lt106_c10 ;
  wire \u2_Display/lt106_c11 ;
  wire \u2_Display/lt106_c12 ;
  wire \u2_Display/lt106_c13 ;
  wire \u2_Display/lt106_c14 ;
  wire \u2_Display/lt106_c15 ;
  wire \u2_Display/lt106_c16 ;
  wire \u2_Display/lt106_c17 ;
  wire \u2_Display/lt106_c18 ;
  wire \u2_Display/lt106_c19 ;
  wire \u2_Display/lt106_c2 ;
  wire \u2_Display/lt106_c20 ;
  wire \u2_Display/lt106_c21 ;
  wire \u2_Display/lt106_c22 ;
  wire \u2_Display/lt106_c23 ;
  wire \u2_Display/lt106_c24 ;
  wire \u2_Display/lt106_c25 ;
  wire \u2_Display/lt106_c26 ;
  wire \u2_Display/lt106_c27 ;
  wire \u2_Display/lt106_c28 ;
  wire \u2_Display/lt106_c29 ;
  wire \u2_Display/lt106_c3 ;
  wire \u2_Display/lt106_c30 ;
  wire \u2_Display/lt106_c31 ;
  wire \u2_Display/lt106_c32 ;
  wire \u2_Display/lt106_c4 ;
  wire \u2_Display/lt106_c5 ;
  wire \u2_Display/lt106_c6 ;
  wire \u2_Display/lt106_c7 ;
  wire \u2_Display/lt106_c8 ;
  wire \u2_Display/lt106_c9 ;
  wire \u2_Display/lt107_c0 ;
  wire \u2_Display/lt107_c1 ;
  wire \u2_Display/lt107_c10 ;
  wire \u2_Display/lt107_c11 ;
  wire \u2_Display/lt107_c12 ;
  wire \u2_Display/lt107_c13 ;
  wire \u2_Display/lt107_c14 ;
  wire \u2_Display/lt107_c15 ;
  wire \u2_Display/lt107_c16 ;
  wire \u2_Display/lt107_c17 ;
  wire \u2_Display/lt107_c18 ;
  wire \u2_Display/lt107_c19 ;
  wire \u2_Display/lt107_c2 ;
  wire \u2_Display/lt107_c20 ;
  wire \u2_Display/lt107_c21 ;
  wire \u2_Display/lt107_c22 ;
  wire \u2_Display/lt107_c23 ;
  wire \u2_Display/lt107_c24 ;
  wire \u2_Display/lt107_c25 ;
  wire \u2_Display/lt107_c26 ;
  wire \u2_Display/lt107_c27 ;
  wire \u2_Display/lt107_c28 ;
  wire \u2_Display/lt107_c29 ;
  wire \u2_Display/lt107_c3 ;
  wire \u2_Display/lt107_c30 ;
  wire \u2_Display/lt107_c31 ;
  wire \u2_Display/lt107_c32 ;
  wire \u2_Display/lt107_c4 ;
  wire \u2_Display/lt107_c5 ;
  wire \u2_Display/lt107_c6 ;
  wire \u2_Display/lt107_c7 ;
  wire \u2_Display/lt107_c8 ;
  wire \u2_Display/lt107_c9 ;
  wire \u2_Display/lt108_c0 ;
  wire \u2_Display/lt108_c1 ;
  wire \u2_Display/lt108_c10 ;
  wire \u2_Display/lt108_c11 ;
  wire \u2_Display/lt108_c12 ;
  wire \u2_Display/lt108_c13 ;
  wire \u2_Display/lt108_c14 ;
  wire \u2_Display/lt108_c15 ;
  wire \u2_Display/lt108_c16 ;
  wire \u2_Display/lt108_c17 ;
  wire \u2_Display/lt108_c18 ;
  wire \u2_Display/lt108_c19 ;
  wire \u2_Display/lt108_c2 ;
  wire \u2_Display/lt108_c20 ;
  wire \u2_Display/lt108_c21 ;
  wire \u2_Display/lt108_c22 ;
  wire \u2_Display/lt108_c23 ;
  wire \u2_Display/lt108_c24 ;
  wire \u2_Display/lt108_c25 ;
  wire \u2_Display/lt108_c26 ;
  wire \u2_Display/lt108_c27 ;
  wire \u2_Display/lt108_c28 ;
  wire \u2_Display/lt108_c29 ;
  wire \u2_Display/lt108_c3 ;
  wire \u2_Display/lt108_c30 ;
  wire \u2_Display/lt108_c31 ;
  wire \u2_Display/lt108_c32 ;
  wire \u2_Display/lt108_c4 ;
  wire \u2_Display/lt108_c5 ;
  wire \u2_Display/lt108_c6 ;
  wire \u2_Display/lt108_c7 ;
  wire \u2_Display/lt108_c8 ;
  wire \u2_Display/lt108_c9 ;
  wire \u2_Display/lt109_c0 ;
  wire \u2_Display/lt109_c1 ;
  wire \u2_Display/lt109_c10 ;
  wire \u2_Display/lt109_c11 ;
  wire \u2_Display/lt109_c12 ;
  wire \u2_Display/lt109_c13 ;
  wire \u2_Display/lt109_c14 ;
  wire \u2_Display/lt109_c15 ;
  wire \u2_Display/lt109_c16 ;
  wire \u2_Display/lt109_c17 ;
  wire \u2_Display/lt109_c18 ;
  wire \u2_Display/lt109_c19 ;
  wire \u2_Display/lt109_c2 ;
  wire \u2_Display/lt109_c20 ;
  wire \u2_Display/lt109_c21 ;
  wire \u2_Display/lt109_c22 ;
  wire \u2_Display/lt109_c23 ;
  wire \u2_Display/lt109_c24 ;
  wire \u2_Display/lt109_c25 ;
  wire \u2_Display/lt109_c26 ;
  wire \u2_Display/lt109_c27 ;
  wire \u2_Display/lt109_c28 ;
  wire \u2_Display/lt109_c29 ;
  wire \u2_Display/lt109_c3 ;
  wire \u2_Display/lt109_c30 ;
  wire \u2_Display/lt109_c31 ;
  wire \u2_Display/lt109_c32 ;
  wire \u2_Display/lt109_c4 ;
  wire \u2_Display/lt109_c5 ;
  wire \u2_Display/lt109_c6 ;
  wire \u2_Display/lt109_c7 ;
  wire \u2_Display/lt109_c8 ;
  wire \u2_Display/lt109_c9 ;
  wire \u2_Display/lt10_2_c0 ;
  wire \u2_Display/lt10_2_c1 ;
  wire \u2_Display/lt10_2_c10 ;
  wire \u2_Display/lt10_2_c11 ;
  wire \u2_Display/lt10_2_c12 ;
  wire \u2_Display/lt10_2_c2 ;
  wire \u2_Display/lt10_2_c3 ;
  wire \u2_Display/lt10_2_c4 ;
  wire \u2_Display/lt10_2_c5 ;
  wire \u2_Display/lt10_2_c6 ;
  wire \u2_Display/lt10_2_c7 ;
  wire \u2_Display/lt10_2_c8 ;
  wire \u2_Display/lt10_2_c9 ;
  wire \u2_Display/lt110_c0 ;
  wire \u2_Display/lt110_c1 ;
  wire \u2_Display/lt110_c10 ;
  wire \u2_Display/lt110_c11 ;
  wire \u2_Display/lt110_c12 ;
  wire \u2_Display/lt110_c13 ;
  wire \u2_Display/lt110_c14 ;
  wire \u2_Display/lt110_c15 ;
  wire \u2_Display/lt110_c16 ;
  wire \u2_Display/lt110_c17 ;
  wire \u2_Display/lt110_c18 ;
  wire \u2_Display/lt110_c19 ;
  wire \u2_Display/lt110_c2 ;
  wire \u2_Display/lt110_c20 ;
  wire \u2_Display/lt110_c21 ;
  wire \u2_Display/lt110_c22 ;
  wire \u2_Display/lt110_c23 ;
  wire \u2_Display/lt110_c24 ;
  wire \u2_Display/lt110_c25 ;
  wire \u2_Display/lt110_c26 ;
  wire \u2_Display/lt110_c27 ;
  wire \u2_Display/lt110_c28 ;
  wire \u2_Display/lt110_c29 ;
  wire \u2_Display/lt110_c3 ;
  wire \u2_Display/lt110_c30 ;
  wire \u2_Display/lt110_c31 ;
  wire \u2_Display/lt110_c32 ;
  wire \u2_Display/lt110_c4 ;
  wire \u2_Display/lt110_c5 ;
  wire \u2_Display/lt110_c6 ;
  wire \u2_Display/lt110_c7 ;
  wire \u2_Display/lt110_c8 ;
  wire \u2_Display/lt110_c9 ;
  wire \u2_Display/lt11_2_c0 ;
  wire \u2_Display/lt11_2_c1 ;
  wire \u2_Display/lt11_2_c10 ;
  wire \u2_Display/lt11_2_c11 ;
  wire \u2_Display/lt11_2_c12 ;
  wire \u2_Display/lt11_2_c13 ;
  wire \u2_Display/lt11_2_c2 ;
  wire \u2_Display/lt11_2_c3 ;
  wire \u2_Display/lt11_2_c4 ;
  wire \u2_Display/lt11_2_c5 ;
  wire \u2_Display/lt11_2_c6 ;
  wire \u2_Display/lt11_2_c7 ;
  wire \u2_Display/lt11_2_c8 ;
  wire \u2_Display/lt11_2_c9 ;
  wire \u2_Display/lt121_c0 ;
  wire \u2_Display/lt121_c1 ;
  wire \u2_Display/lt121_c10 ;
  wire \u2_Display/lt121_c11 ;
  wire \u2_Display/lt121_c12 ;
  wire \u2_Display/lt121_c13 ;
  wire \u2_Display/lt121_c14 ;
  wire \u2_Display/lt121_c15 ;
  wire \u2_Display/lt121_c16 ;
  wire \u2_Display/lt121_c17 ;
  wire \u2_Display/lt121_c18 ;
  wire \u2_Display/lt121_c19 ;
  wire \u2_Display/lt121_c2 ;
  wire \u2_Display/lt121_c20 ;
  wire \u2_Display/lt121_c21 ;
  wire \u2_Display/lt121_c22 ;
  wire \u2_Display/lt121_c23 ;
  wire \u2_Display/lt121_c24 ;
  wire \u2_Display/lt121_c25 ;
  wire \u2_Display/lt121_c26 ;
  wire \u2_Display/lt121_c27 ;
  wire \u2_Display/lt121_c28 ;
  wire \u2_Display/lt121_c29 ;
  wire \u2_Display/lt121_c3 ;
  wire \u2_Display/lt121_c30 ;
  wire \u2_Display/lt121_c31 ;
  wire \u2_Display/lt121_c32 ;
  wire \u2_Display/lt121_c4 ;
  wire \u2_Display/lt121_c5 ;
  wire \u2_Display/lt121_c6 ;
  wire \u2_Display/lt121_c7 ;
  wire \u2_Display/lt121_c8 ;
  wire \u2_Display/lt121_c9 ;
  wire \u2_Display/lt122_c0 ;
  wire \u2_Display/lt122_c1 ;
  wire \u2_Display/lt122_c10 ;
  wire \u2_Display/lt122_c11 ;
  wire \u2_Display/lt122_c12 ;
  wire \u2_Display/lt122_c13 ;
  wire \u2_Display/lt122_c14 ;
  wire \u2_Display/lt122_c15 ;
  wire \u2_Display/lt122_c16 ;
  wire \u2_Display/lt122_c17 ;
  wire \u2_Display/lt122_c18 ;
  wire \u2_Display/lt122_c19 ;
  wire \u2_Display/lt122_c2 ;
  wire \u2_Display/lt122_c20 ;
  wire \u2_Display/lt122_c21 ;
  wire \u2_Display/lt122_c22 ;
  wire \u2_Display/lt122_c23 ;
  wire \u2_Display/lt122_c24 ;
  wire \u2_Display/lt122_c25 ;
  wire \u2_Display/lt122_c26 ;
  wire \u2_Display/lt122_c27 ;
  wire \u2_Display/lt122_c28 ;
  wire \u2_Display/lt122_c29 ;
  wire \u2_Display/lt122_c3 ;
  wire \u2_Display/lt122_c30 ;
  wire \u2_Display/lt122_c31 ;
  wire \u2_Display/lt122_c32 ;
  wire \u2_Display/lt122_c4 ;
  wire \u2_Display/lt122_c5 ;
  wire \u2_Display/lt122_c6 ;
  wire \u2_Display/lt122_c7 ;
  wire \u2_Display/lt122_c8 ;
  wire \u2_Display/lt122_c9 ;
  wire \u2_Display/lt123_c0 ;
  wire \u2_Display/lt123_c1 ;
  wire \u2_Display/lt123_c10 ;
  wire \u2_Display/lt123_c11 ;
  wire \u2_Display/lt123_c12 ;
  wire \u2_Display/lt123_c13 ;
  wire \u2_Display/lt123_c14 ;
  wire \u2_Display/lt123_c15 ;
  wire \u2_Display/lt123_c16 ;
  wire \u2_Display/lt123_c17 ;
  wire \u2_Display/lt123_c18 ;
  wire \u2_Display/lt123_c19 ;
  wire \u2_Display/lt123_c2 ;
  wire \u2_Display/lt123_c20 ;
  wire \u2_Display/lt123_c21 ;
  wire \u2_Display/lt123_c22 ;
  wire \u2_Display/lt123_c23 ;
  wire \u2_Display/lt123_c24 ;
  wire \u2_Display/lt123_c25 ;
  wire \u2_Display/lt123_c26 ;
  wire \u2_Display/lt123_c27 ;
  wire \u2_Display/lt123_c28 ;
  wire \u2_Display/lt123_c29 ;
  wire \u2_Display/lt123_c3 ;
  wire \u2_Display/lt123_c30 ;
  wire \u2_Display/lt123_c31 ;
  wire \u2_Display/lt123_c32 ;
  wire \u2_Display/lt123_c4 ;
  wire \u2_Display/lt123_c5 ;
  wire \u2_Display/lt123_c6 ;
  wire \u2_Display/lt123_c7 ;
  wire \u2_Display/lt123_c8 ;
  wire \u2_Display/lt123_c9 ;
  wire \u2_Display/lt124_c0 ;
  wire \u2_Display/lt124_c1 ;
  wire \u2_Display/lt124_c10 ;
  wire \u2_Display/lt124_c11 ;
  wire \u2_Display/lt124_c12 ;
  wire \u2_Display/lt124_c13 ;
  wire \u2_Display/lt124_c14 ;
  wire \u2_Display/lt124_c15 ;
  wire \u2_Display/lt124_c16 ;
  wire \u2_Display/lt124_c17 ;
  wire \u2_Display/lt124_c18 ;
  wire \u2_Display/lt124_c19 ;
  wire \u2_Display/lt124_c2 ;
  wire \u2_Display/lt124_c20 ;
  wire \u2_Display/lt124_c21 ;
  wire \u2_Display/lt124_c22 ;
  wire \u2_Display/lt124_c23 ;
  wire \u2_Display/lt124_c24 ;
  wire \u2_Display/lt124_c25 ;
  wire \u2_Display/lt124_c26 ;
  wire \u2_Display/lt124_c27 ;
  wire \u2_Display/lt124_c28 ;
  wire \u2_Display/lt124_c29 ;
  wire \u2_Display/lt124_c3 ;
  wire \u2_Display/lt124_c30 ;
  wire \u2_Display/lt124_c31 ;
  wire \u2_Display/lt124_c32 ;
  wire \u2_Display/lt124_c4 ;
  wire \u2_Display/lt124_c5 ;
  wire \u2_Display/lt124_c6 ;
  wire \u2_Display/lt124_c7 ;
  wire \u2_Display/lt124_c8 ;
  wire \u2_Display/lt124_c9 ;
  wire \u2_Display/lt125_c0 ;
  wire \u2_Display/lt125_c1 ;
  wire \u2_Display/lt125_c10 ;
  wire \u2_Display/lt125_c11 ;
  wire \u2_Display/lt125_c12 ;
  wire \u2_Display/lt125_c13 ;
  wire \u2_Display/lt125_c14 ;
  wire \u2_Display/lt125_c15 ;
  wire \u2_Display/lt125_c16 ;
  wire \u2_Display/lt125_c17 ;
  wire \u2_Display/lt125_c18 ;
  wire \u2_Display/lt125_c19 ;
  wire \u2_Display/lt125_c2 ;
  wire \u2_Display/lt125_c20 ;
  wire \u2_Display/lt125_c21 ;
  wire \u2_Display/lt125_c22 ;
  wire \u2_Display/lt125_c23 ;
  wire \u2_Display/lt125_c24 ;
  wire \u2_Display/lt125_c25 ;
  wire \u2_Display/lt125_c26 ;
  wire \u2_Display/lt125_c27 ;
  wire \u2_Display/lt125_c28 ;
  wire \u2_Display/lt125_c29 ;
  wire \u2_Display/lt125_c3 ;
  wire \u2_Display/lt125_c30 ;
  wire \u2_Display/lt125_c31 ;
  wire \u2_Display/lt125_c32 ;
  wire \u2_Display/lt125_c4 ;
  wire \u2_Display/lt125_c5 ;
  wire \u2_Display/lt125_c6 ;
  wire \u2_Display/lt125_c7 ;
  wire \u2_Display/lt125_c8 ;
  wire \u2_Display/lt125_c9 ;
  wire \u2_Display/lt126_c0 ;
  wire \u2_Display/lt126_c1 ;
  wire \u2_Display/lt126_c10 ;
  wire \u2_Display/lt126_c11 ;
  wire \u2_Display/lt126_c12 ;
  wire \u2_Display/lt126_c13 ;
  wire \u2_Display/lt126_c14 ;
  wire \u2_Display/lt126_c15 ;
  wire \u2_Display/lt126_c16 ;
  wire \u2_Display/lt126_c17 ;
  wire \u2_Display/lt126_c18 ;
  wire \u2_Display/lt126_c19 ;
  wire \u2_Display/lt126_c2 ;
  wire \u2_Display/lt126_c20 ;
  wire \u2_Display/lt126_c21 ;
  wire \u2_Display/lt126_c22 ;
  wire \u2_Display/lt126_c23 ;
  wire \u2_Display/lt126_c24 ;
  wire \u2_Display/lt126_c25 ;
  wire \u2_Display/lt126_c26 ;
  wire \u2_Display/lt126_c27 ;
  wire \u2_Display/lt126_c28 ;
  wire \u2_Display/lt126_c29 ;
  wire \u2_Display/lt126_c3 ;
  wire \u2_Display/lt126_c30 ;
  wire \u2_Display/lt126_c31 ;
  wire \u2_Display/lt126_c32 ;
  wire \u2_Display/lt126_c4 ;
  wire \u2_Display/lt126_c5 ;
  wire \u2_Display/lt126_c6 ;
  wire \u2_Display/lt126_c7 ;
  wire \u2_Display/lt126_c8 ;
  wire \u2_Display/lt126_c9 ;
  wire \u2_Display/lt127_c0 ;
  wire \u2_Display/lt127_c1 ;
  wire \u2_Display/lt127_c10 ;
  wire \u2_Display/lt127_c11 ;
  wire \u2_Display/lt127_c12 ;
  wire \u2_Display/lt127_c13 ;
  wire \u2_Display/lt127_c14 ;
  wire \u2_Display/lt127_c15 ;
  wire \u2_Display/lt127_c16 ;
  wire \u2_Display/lt127_c17 ;
  wire \u2_Display/lt127_c18 ;
  wire \u2_Display/lt127_c19 ;
  wire \u2_Display/lt127_c2 ;
  wire \u2_Display/lt127_c20 ;
  wire \u2_Display/lt127_c21 ;
  wire \u2_Display/lt127_c22 ;
  wire \u2_Display/lt127_c23 ;
  wire \u2_Display/lt127_c24 ;
  wire \u2_Display/lt127_c25 ;
  wire \u2_Display/lt127_c26 ;
  wire \u2_Display/lt127_c27 ;
  wire \u2_Display/lt127_c28 ;
  wire \u2_Display/lt127_c29 ;
  wire \u2_Display/lt127_c3 ;
  wire \u2_Display/lt127_c30 ;
  wire \u2_Display/lt127_c31 ;
  wire \u2_Display/lt127_c32 ;
  wire \u2_Display/lt127_c4 ;
  wire \u2_Display/lt127_c5 ;
  wire \u2_Display/lt127_c6 ;
  wire \u2_Display/lt127_c7 ;
  wire \u2_Display/lt127_c8 ;
  wire \u2_Display/lt127_c9 ;
  wire \u2_Display/lt128_c0 ;
  wire \u2_Display/lt128_c1 ;
  wire \u2_Display/lt128_c10 ;
  wire \u2_Display/lt128_c11 ;
  wire \u2_Display/lt128_c12 ;
  wire \u2_Display/lt128_c13 ;
  wire \u2_Display/lt128_c14 ;
  wire \u2_Display/lt128_c15 ;
  wire \u2_Display/lt128_c16 ;
  wire \u2_Display/lt128_c17 ;
  wire \u2_Display/lt128_c18 ;
  wire \u2_Display/lt128_c19 ;
  wire \u2_Display/lt128_c2 ;
  wire \u2_Display/lt128_c20 ;
  wire \u2_Display/lt128_c21 ;
  wire \u2_Display/lt128_c22 ;
  wire \u2_Display/lt128_c23 ;
  wire \u2_Display/lt128_c24 ;
  wire \u2_Display/lt128_c25 ;
  wire \u2_Display/lt128_c26 ;
  wire \u2_Display/lt128_c27 ;
  wire \u2_Display/lt128_c28 ;
  wire \u2_Display/lt128_c29 ;
  wire \u2_Display/lt128_c3 ;
  wire \u2_Display/lt128_c30 ;
  wire \u2_Display/lt128_c31 ;
  wire \u2_Display/lt128_c32 ;
  wire \u2_Display/lt128_c4 ;
  wire \u2_Display/lt128_c5 ;
  wire \u2_Display/lt128_c6 ;
  wire \u2_Display/lt128_c7 ;
  wire \u2_Display/lt128_c8 ;
  wire \u2_Display/lt128_c9 ;
  wire \u2_Display/lt129_c0 ;
  wire \u2_Display/lt129_c1 ;
  wire \u2_Display/lt129_c10 ;
  wire \u2_Display/lt129_c11 ;
  wire \u2_Display/lt129_c12 ;
  wire \u2_Display/lt129_c13 ;
  wire \u2_Display/lt129_c14 ;
  wire \u2_Display/lt129_c15 ;
  wire \u2_Display/lt129_c16 ;
  wire \u2_Display/lt129_c17 ;
  wire \u2_Display/lt129_c18 ;
  wire \u2_Display/lt129_c19 ;
  wire \u2_Display/lt129_c2 ;
  wire \u2_Display/lt129_c20 ;
  wire \u2_Display/lt129_c21 ;
  wire \u2_Display/lt129_c22 ;
  wire \u2_Display/lt129_c23 ;
  wire \u2_Display/lt129_c24 ;
  wire \u2_Display/lt129_c25 ;
  wire \u2_Display/lt129_c26 ;
  wire \u2_Display/lt129_c27 ;
  wire \u2_Display/lt129_c28 ;
  wire \u2_Display/lt129_c29 ;
  wire \u2_Display/lt129_c3 ;
  wire \u2_Display/lt129_c30 ;
  wire \u2_Display/lt129_c31 ;
  wire \u2_Display/lt129_c32 ;
  wire \u2_Display/lt129_c4 ;
  wire \u2_Display/lt129_c5 ;
  wire \u2_Display/lt129_c6 ;
  wire \u2_Display/lt129_c7 ;
  wire \u2_Display/lt129_c8 ;
  wire \u2_Display/lt129_c9 ;
  wire \u2_Display/lt130_c0 ;
  wire \u2_Display/lt130_c1 ;
  wire \u2_Display/lt130_c10 ;
  wire \u2_Display/lt130_c11 ;
  wire \u2_Display/lt130_c12 ;
  wire \u2_Display/lt130_c13 ;
  wire \u2_Display/lt130_c14 ;
  wire \u2_Display/lt130_c15 ;
  wire \u2_Display/lt130_c16 ;
  wire \u2_Display/lt130_c17 ;
  wire \u2_Display/lt130_c18 ;
  wire \u2_Display/lt130_c19 ;
  wire \u2_Display/lt130_c2 ;
  wire \u2_Display/lt130_c20 ;
  wire \u2_Display/lt130_c21 ;
  wire \u2_Display/lt130_c22 ;
  wire \u2_Display/lt130_c23 ;
  wire \u2_Display/lt130_c24 ;
  wire \u2_Display/lt130_c25 ;
  wire \u2_Display/lt130_c26 ;
  wire \u2_Display/lt130_c27 ;
  wire \u2_Display/lt130_c28 ;
  wire \u2_Display/lt130_c29 ;
  wire \u2_Display/lt130_c3 ;
  wire \u2_Display/lt130_c30 ;
  wire \u2_Display/lt130_c31 ;
  wire \u2_Display/lt130_c32 ;
  wire \u2_Display/lt130_c4 ;
  wire \u2_Display/lt130_c5 ;
  wire \u2_Display/lt130_c6 ;
  wire \u2_Display/lt130_c7 ;
  wire \u2_Display/lt130_c8 ;
  wire \u2_Display/lt130_c9 ;
  wire \u2_Display/lt131_c0 ;
  wire \u2_Display/lt131_c1 ;
  wire \u2_Display/lt131_c10 ;
  wire \u2_Display/lt131_c11 ;
  wire \u2_Display/lt131_c12 ;
  wire \u2_Display/lt131_c13 ;
  wire \u2_Display/lt131_c14 ;
  wire \u2_Display/lt131_c15 ;
  wire \u2_Display/lt131_c16 ;
  wire \u2_Display/lt131_c17 ;
  wire \u2_Display/lt131_c18 ;
  wire \u2_Display/lt131_c19 ;
  wire \u2_Display/lt131_c2 ;
  wire \u2_Display/lt131_c20 ;
  wire \u2_Display/lt131_c21 ;
  wire \u2_Display/lt131_c22 ;
  wire \u2_Display/lt131_c23 ;
  wire \u2_Display/lt131_c24 ;
  wire \u2_Display/lt131_c25 ;
  wire \u2_Display/lt131_c26 ;
  wire \u2_Display/lt131_c27 ;
  wire \u2_Display/lt131_c28 ;
  wire \u2_Display/lt131_c29 ;
  wire \u2_Display/lt131_c3 ;
  wire \u2_Display/lt131_c30 ;
  wire \u2_Display/lt131_c31 ;
  wire \u2_Display/lt131_c32 ;
  wire \u2_Display/lt131_c4 ;
  wire \u2_Display/lt131_c5 ;
  wire \u2_Display/lt131_c6 ;
  wire \u2_Display/lt131_c7 ;
  wire \u2_Display/lt131_c8 ;
  wire \u2_Display/lt131_c9 ;
  wire \u2_Display/lt132_c0 ;
  wire \u2_Display/lt132_c1 ;
  wire \u2_Display/lt132_c10 ;
  wire \u2_Display/lt132_c11 ;
  wire \u2_Display/lt132_c12 ;
  wire \u2_Display/lt132_c13 ;
  wire \u2_Display/lt132_c14 ;
  wire \u2_Display/lt132_c15 ;
  wire \u2_Display/lt132_c16 ;
  wire \u2_Display/lt132_c17 ;
  wire \u2_Display/lt132_c18 ;
  wire \u2_Display/lt132_c19 ;
  wire \u2_Display/lt132_c2 ;
  wire \u2_Display/lt132_c20 ;
  wire \u2_Display/lt132_c21 ;
  wire \u2_Display/lt132_c22 ;
  wire \u2_Display/lt132_c23 ;
  wire \u2_Display/lt132_c24 ;
  wire \u2_Display/lt132_c25 ;
  wire \u2_Display/lt132_c26 ;
  wire \u2_Display/lt132_c27 ;
  wire \u2_Display/lt132_c28 ;
  wire \u2_Display/lt132_c29 ;
  wire \u2_Display/lt132_c3 ;
  wire \u2_Display/lt132_c30 ;
  wire \u2_Display/lt132_c31 ;
  wire \u2_Display/lt132_c32 ;
  wire \u2_Display/lt132_c4 ;
  wire \u2_Display/lt132_c5 ;
  wire \u2_Display/lt132_c6 ;
  wire \u2_Display/lt132_c7 ;
  wire \u2_Display/lt132_c8 ;
  wire \u2_Display/lt132_c9 ;
  wire \u2_Display/lt133_c0 ;
  wire \u2_Display/lt133_c1 ;
  wire \u2_Display/lt133_c10 ;
  wire \u2_Display/lt133_c11 ;
  wire \u2_Display/lt133_c12 ;
  wire \u2_Display/lt133_c13 ;
  wire \u2_Display/lt133_c14 ;
  wire \u2_Display/lt133_c15 ;
  wire \u2_Display/lt133_c16 ;
  wire \u2_Display/lt133_c17 ;
  wire \u2_Display/lt133_c18 ;
  wire \u2_Display/lt133_c19 ;
  wire \u2_Display/lt133_c2 ;
  wire \u2_Display/lt133_c20 ;
  wire \u2_Display/lt133_c21 ;
  wire \u2_Display/lt133_c22 ;
  wire \u2_Display/lt133_c23 ;
  wire \u2_Display/lt133_c24 ;
  wire \u2_Display/lt133_c25 ;
  wire \u2_Display/lt133_c26 ;
  wire \u2_Display/lt133_c27 ;
  wire \u2_Display/lt133_c28 ;
  wire \u2_Display/lt133_c29 ;
  wire \u2_Display/lt133_c3 ;
  wire \u2_Display/lt133_c30 ;
  wire \u2_Display/lt133_c31 ;
  wire \u2_Display/lt133_c32 ;
  wire \u2_Display/lt133_c4 ;
  wire \u2_Display/lt133_c5 ;
  wire \u2_Display/lt133_c6 ;
  wire \u2_Display/lt133_c7 ;
  wire \u2_Display/lt133_c8 ;
  wire \u2_Display/lt133_c9 ;
  wire \u2_Display/lt134_c0 ;
  wire \u2_Display/lt134_c1 ;
  wire \u2_Display/lt134_c10 ;
  wire \u2_Display/lt134_c11 ;
  wire \u2_Display/lt134_c12 ;
  wire \u2_Display/lt134_c13 ;
  wire \u2_Display/lt134_c14 ;
  wire \u2_Display/lt134_c15 ;
  wire \u2_Display/lt134_c16 ;
  wire \u2_Display/lt134_c17 ;
  wire \u2_Display/lt134_c18 ;
  wire \u2_Display/lt134_c19 ;
  wire \u2_Display/lt134_c2 ;
  wire \u2_Display/lt134_c20 ;
  wire \u2_Display/lt134_c21 ;
  wire \u2_Display/lt134_c22 ;
  wire \u2_Display/lt134_c23 ;
  wire \u2_Display/lt134_c24 ;
  wire \u2_Display/lt134_c25 ;
  wire \u2_Display/lt134_c26 ;
  wire \u2_Display/lt134_c27 ;
  wire \u2_Display/lt134_c28 ;
  wire \u2_Display/lt134_c29 ;
  wire \u2_Display/lt134_c3 ;
  wire \u2_Display/lt134_c30 ;
  wire \u2_Display/lt134_c31 ;
  wire \u2_Display/lt134_c32 ;
  wire \u2_Display/lt134_c4 ;
  wire \u2_Display/lt134_c5 ;
  wire \u2_Display/lt134_c6 ;
  wire \u2_Display/lt134_c7 ;
  wire \u2_Display/lt134_c8 ;
  wire \u2_Display/lt134_c9 ;
  wire \u2_Display/lt135_c0 ;
  wire \u2_Display/lt135_c1 ;
  wire \u2_Display/lt135_c10 ;
  wire \u2_Display/lt135_c11 ;
  wire \u2_Display/lt135_c12 ;
  wire \u2_Display/lt135_c13 ;
  wire \u2_Display/lt135_c14 ;
  wire \u2_Display/lt135_c15 ;
  wire \u2_Display/lt135_c16 ;
  wire \u2_Display/lt135_c17 ;
  wire \u2_Display/lt135_c18 ;
  wire \u2_Display/lt135_c19 ;
  wire \u2_Display/lt135_c2 ;
  wire \u2_Display/lt135_c20 ;
  wire \u2_Display/lt135_c21 ;
  wire \u2_Display/lt135_c22 ;
  wire \u2_Display/lt135_c23 ;
  wire \u2_Display/lt135_c24 ;
  wire \u2_Display/lt135_c25 ;
  wire \u2_Display/lt135_c26 ;
  wire \u2_Display/lt135_c27 ;
  wire \u2_Display/lt135_c28 ;
  wire \u2_Display/lt135_c29 ;
  wire \u2_Display/lt135_c3 ;
  wire \u2_Display/lt135_c30 ;
  wire \u2_Display/lt135_c31 ;
  wire \u2_Display/lt135_c32 ;
  wire \u2_Display/lt135_c4 ;
  wire \u2_Display/lt135_c5 ;
  wire \u2_Display/lt135_c6 ;
  wire \u2_Display/lt135_c7 ;
  wire \u2_Display/lt135_c8 ;
  wire \u2_Display/lt135_c9 ;
  wire \u2_Display/lt136_c0 ;
  wire \u2_Display/lt136_c1 ;
  wire \u2_Display/lt136_c10 ;
  wire \u2_Display/lt136_c11 ;
  wire \u2_Display/lt136_c12 ;
  wire \u2_Display/lt136_c13 ;
  wire \u2_Display/lt136_c14 ;
  wire \u2_Display/lt136_c15 ;
  wire \u2_Display/lt136_c16 ;
  wire \u2_Display/lt136_c17 ;
  wire \u2_Display/lt136_c18 ;
  wire \u2_Display/lt136_c19 ;
  wire \u2_Display/lt136_c2 ;
  wire \u2_Display/lt136_c20 ;
  wire \u2_Display/lt136_c21 ;
  wire \u2_Display/lt136_c22 ;
  wire \u2_Display/lt136_c23 ;
  wire \u2_Display/lt136_c24 ;
  wire \u2_Display/lt136_c25 ;
  wire \u2_Display/lt136_c26 ;
  wire \u2_Display/lt136_c27 ;
  wire \u2_Display/lt136_c28 ;
  wire \u2_Display/lt136_c29 ;
  wire \u2_Display/lt136_c3 ;
  wire \u2_Display/lt136_c30 ;
  wire \u2_Display/lt136_c31 ;
  wire \u2_Display/lt136_c32 ;
  wire \u2_Display/lt136_c4 ;
  wire \u2_Display/lt136_c5 ;
  wire \u2_Display/lt136_c6 ;
  wire \u2_Display/lt136_c7 ;
  wire \u2_Display/lt136_c8 ;
  wire \u2_Display/lt136_c9 ;
  wire \u2_Display/lt137_c0 ;
  wire \u2_Display/lt137_c1 ;
  wire \u2_Display/lt137_c10 ;
  wire \u2_Display/lt137_c11 ;
  wire \u2_Display/lt137_c12 ;
  wire \u2_Display/lt137_c13 ;
  wire \u2_Display/lt137_c14 ;
  wire \u2_Display/lt137_c15 ;
  wire \u2_Display/lt137_c16 ;
  wire \u2_Display/lt137_c17 ;
  wire \u2_Display/lt137_c18 ;
  wire \u2_Display/lt137_c19 ;
  wire \u2_Display/lt137_c2 ;
  wire \u2_Display/lt137_c20 ;
  wire \u2_Display/lt137_c21 ;
  wire \u2_Display/lt137_c22 ;
  wire \u2_Display/lt137_c23 ;
  wire \u2_Display/lt137_c24 ;
  wire \u2_Display/lt137_c25 ;
  wire \u2_Display/lt137_c26 ;
  wire \u2_Display/lt137_c27 ;
  wire \u2_Display/lt137_c28 ;
  wire \u2_Display/lt137_c29 ;
  wire \u2_Display/lt137_c3 ;
  wire \u2_Display/lt137_c30 ;
  wire \u2_Display/lt137_c31 ;
  wire \u2_Display/lt137_c32 ;
  wire \u2_Display/lt137_c4 ;
  wire \u2_Display/lt137_c5 ;
  wire \u2_Display/lt137_c6 ;
  wire \u2_Display/lt137_c7 ;
  wire \u2_Display/lt137_c8 ;
  wire \u2_Display/lt137_c9 ;
  wire \u2_Display/lt138_c0 ;
  wire \u2_Display/lt138_c1 ;
  wire \u2_Display/lt138_c10 ;
  wire \u2_Display/lt138_c11 ;
  wire \u2_Display/lt138_c12 ;
  wire \u2_Display/lt138_c13 ;
  wire \u2_Display/lt138_c14 ;
  wire \u2_Display/lt138_c15 ;
  wire \u2_Display/lt138_c16 ;
  wire \u2_Display/lt138_c17 ;
  wire \u2_Display/lt138_c18 ;
  wire \u2_Display/lt138_c19 ;
  wire \u2_Display/lt138_c2 ;
  wire \u2_Display/lt138_c20 ;
  wire \u2_Display/lt138_c21 ;
  wire \u2_Display/lt138_c22 ;
  wire \u2_Display/lt138_c23 ;
  wire \u2_Display/lt138_c24 ;
  wire \u2_Display/lt138_c25 ;
  wire \u2_Display/lt138_c26 ;
  wire \u2_Display/lt138_c27 ;
  wire \u2_Display/lt138_c28 ;
  wire \u2_Display/lt138_c29 ;
  wire \u2_Display/lt138_c3 ;
  wire \u2_Display/lt138_c30 ;
  wire \u2_Display/lt138_c31 ;
  wire \u2_Display/lt138_c32 ;
  wire \u2_Display/lt138_c4 ;
  wire \u2_Display/lt138_c5 ;
  wire \u2_Display/lt138_c6 ;
  wire \u2_Display/lt138_c7 ;
  wire \u2_Display/lt138_c8 ;
  wire \u2_Display/lt138_c9 ;
  wire \u2_Display/lt139_c0 ;
  wire \u2_Display/lt139_c1 ;
  wire \u2_Display/lt139_c10 ;
  wire \u2_Display/lt139_c11 ;
  wire \u2_Display/lt139_c12 ;
  wire \u2_Display/lt139_c13 ;
  wire \u2_Display/lt139_c14 ;
  wire \u2_Display/lt139_c15 ;
  wire \u2_Display/lt139_c16 ;
  wire \u2_Display/lt139_c17 ;
  wire \u2_Display/lt139_c18 ;
  wire \u2_Display/lt139_c19 ;
  wire \u2_Display/lt139_c2 ;
  wire \u2_Display/lt139_c20 ;
  wire \u2_Display/lt139_c21 ;
  wire \u2_Display/lt139_c22 ;
  wire \u2_Display/lt139_c23 ;
  wire \u2_Display/lt139_c24 ;
  wire \u2_Display/lt139_c25 ;
  wire \u2_Display/lt139_c26 ;
  wire \u2_Display/lt139_c27 ;
  wire \u2_Display/lt139_c28 ;
  wire \u2_Display/lt139_c29 ;
  wire \u2_Display/lt139_c3 ;
  wire \u2_Display/lt139_c30 ;
  wire \u2_Display/lt139_c31 ;
  wire \u2_Display/lt139_c32 ;
  wire \u2_Display/lt139_c4 ;
  wire \u2_Display/lt139_c5 ;
  wire \u2_Display/lt139_c6 ;
  wire \u2_Display/lt139_c7 ;
  wire \u2_Display/lt139_c8 ;
  wire \u2_Display/lt139_c9 ;
  wire \u2_Display/lt140_c0 ;
  wire \u2_Display/lt140_c1 ;
  wire \u2_Display/lt140_c10 ;
  wire \u2_Display/lt140_c11 ;
  wire \u2_Display/lt140_c12 ;
  wire \u2_Display/lt140_c13 ;
  wire \u2_Display/lt140_c14 ;
  wire \u2_Display/lt140_c15 ;
  wire \u2_Display/lt140_c16 ;
  wire \u2_Display/lt140_c17 ;
  wire \u2_Display/lt140_c18 ;
  wire \u2_Display/lt140_c19 ;
  wire \u2_Display/lt140_c2 ;
  wire \u2_Display/lt140_c20 ;
  wire \u2_Display/lt140_c21 ;
  wire \u2_Display/lt140_c22 ;
  wire \u2_Display/lt140_c23 ;
  wire \u2_Display/lt140_c24 ;
  wire \u2_Display/lt140_c25 ;
  wire \u2_Display/lt140_c26 ;
  wire \u2_Display/lt140_c27 ;
  wire \u2_Display/lt140_c28 ;
  wire \u2_Display/lt140_c29 ;
  wire \u2_Display/lt140_c3 ;
  wire \u2_Display/lt140_c30 ;
  wire \u2_Display/lt140_c31 ;
  wire \u2_Display/lt140_c32 ;
  wire \u2_Display/lt140_c4 ;
  wire \u2_Display/lt140_c5 ;
  wire \u2_Display/lt140_c6 ;
  wire \u2_Display/lt140_c7 ;
  wire \u2_Display/lt140_c8 ;
  wire \u2_Display/lt140_c9 ;
  wire \u2_Display/lt141_c0 ;
  wire \u2_Display/lt141_c1 ;
  wire \u2_Display/lt141_c10 ;
  wire \u2_Display/lt141_c11 ;
  wire \u2_Display/lt141_c12 ;
  wire \u2_Display/lt141_c13 ;
  wire \u2_Display/lt141_c14 ;
  wire \u2_Display/lt141_c15 ;
  wire \u2_Display/lt141_c16 ;
  wire \u2_Display/lt141_c17 ;
  wire \u2_Display/lt141_c18 ;
  wire \u2_Display/lt141_c19 ;
  wire \u2_Display/lt141_c2 ;
  wire \u2_Display/lt141_c20 ;
  wire \u2_Display/lt141_c21 ;
  wire \u2_Display/lt141_c22 ;
  wire \u2_Display/lt141_c23 ;
  wire \u2_Display/lt141_c24 ;
  wire \u2_Display/lt141_c25 ;
  wire \u2_Display/lt141_c26 ;
  wire \u2_Display/lt141_c27 ;
  wire \u2_Display/lt141_c28 ;
  wire \u2_Display/lt141_c29 ;
  wire \u2_Display/lt141_c3 ;
  wire \u2_Display/lt141_c30 ;
  wire \u2_Display/lt141_c31 ;
  wire \u2_Display/lt141_c32 ;
  wire \u2_Display/lt141_c4 ;
  wire \u2_Display/lt141_c5 ;
  wire \u2_Display/lt141_c6 ;
  wire \u2_Display/lt141_c7 ;
  wire \u2_Display/lt141_c8 ;
  wire \u2_Display/lt141_c9 ;
  wire \u2_Display/lt142_c0 ;
  wire \u2_Display/lt142_c1 ;
  wire \u2_Display/lt142_c10 ;
  wire \u2_Display/lt142_c11 ;
  wire \u2_Display/lt142_c12 ;
  wire \u2_Display/lt142_c13 ;
  wire \u2_Display/lt142_c14 ;
  wire \u2_Display/lt142_c15 ;
  wire \u2_Display/lt142_c16 ;
  wire \u2_Display/lt142_c17 ;
  wire \u2_Display/lt142_c18 ;
  wire \u2_Display/lt142_c19 ;
  wire \u2_Display/lt142_c2 ;
  wire \u2_Display/lt142_c20 ;
  wire \u2_Display/lt142_c21 ;
  wire \u2_Display/lt142_c22 ;
  wire \u2_Display/lt142_c23 ;
  wire \u2_Display/lt142_c24 ;
  wire \u2_Display/lt142_c25 ;
  wire \u2_Display/lt142_c26 ;
  wire \u2_Display/lt142_c27 ;
  wire \u2_Display/lt142_c28 ;
  wire \u2_Display/lt142_c29 ;
  wire \u2_Display/lt142_c3 ;
  wire \u2_Display/lt142_c30 ;
  wire \u2_Display/lt142_c31 ;
  wire \u2_Display/lt142_c32 ;
  wire \u2_Display/lt142_c4 ;
  wire \u2_Display/lt142_c5 ;
  wire \u2_Display/lt142_c6 ;
  wire \u2_Display/lt142_c7 ;
  wire \u2_Display/lt142_c8 ;
  wire \u2_Display/lt142_c9 ;
  wire \u2_Display/lt143_c0 ;
  wire \u2_Display/lt143_c1 ;
  wire \u2_Display/lt143_c10 ;
  wire \u2_Display/lt143_c11 ;
  wire \u2_Display/lt143_c12 ;
  wire \u2_Display/lt143_c13 ;
  wire \u2_Display/lt143_c14 ;
  wire \u2_Display/lt143_c15 ;
  wire \u2_Display/lt143_c16 ;
  wire \u2_Display/lt143_c17 ;
  wire \u2_Display/lt143_c18 ;
  wire \u2_Display/lt143_c19 ;
  wire \u2_Display/lt143_c2 ;
  wire \u2_Display/lt143_c20 ;
  wire \u2_Display/lt143_c21 ;
  wire \u2_Display/lt143_c22 ;
  wire \u2_Display/lt143_c23 ;
  wire \u2_Display/lt143_c24 ;
  wire \u2_Display/lt143_c25 ;
  wire \u2_Display/lt143_c26 ;
  wire \u2_Display/lt143_c27 ;
  wire \u2_Display/lt143_c28 ;
  wire \u2_Display/lt143_c29 ;
  wire \u2_Display/lt143_c3 ;
  wire \u2_Display/lt143_c30 ;
  wire \u2_Display/lt143_c31 ;
  wire \u2_Display/lt143_c32 ;
  wire \u2_Display/lt143_c4 ;
  wire \u2_Display/lt143_c5 ;
  wire \u2_Display/lt143_c6 ;
  wire \u2_Display/lt143_c7 ;
  wire \u2_Display/lt143_c8 ;
  wire \u2_Display/lt143_c9 ;
  wire \u2_Display/lt154_c0 ;
  wire \u2_Display/lt154_c1 ;
  wire \u2_Display/lt154_c10 ;
  wire \u2_Display/lt154_c11 ;
  wire \u2_Display/lt154_c12 ;
  wire \u2_Display/lt154_c13 ;
  wire \u2_Display/lt154_c14 ;
  wire \u2_Display/lt154_c15 ;
  wire \u2_Display/lt154_c16 ;
  wire \u2_Display/lt154_c17 ;
  wire \u2_Display/lt154_c18 ;
  wire \u2_Display/lt154_c19 ;
  wire \u2_Display/lt154_c2 ;
  wire \u2_Display/lt154_c20 ;
  wire \u2_Display/lt154_c21 ;
  wire \u2_Display/lt154_c22 ;
  wire \u2_Display/lt154_c23 ;
  wire \u2_Display/lt154_c24 ;
  wire \u2_Display/lt154_c25 ;
  wire \u2_Display/lt154_c26 ;
  wire \u2_Display/lt154_c27 ;
  wire \u2_Display/lt154_c28 ;
  wire \u2_Display/lt154_c29 ;
  wire \u2_Display/lt154_c3 ;
  wire \u2_Display/lt154_c30 ;
  wire \u2_Display/lt154_c31 ;
  wire \u2_Display/lt154_c32 ;
  wire \u2_Display/lt154_c4 ;
  wire \u2_Display/lt154_c5 ;
  wire \u2_Display/lt154_c6 ;
  wire \u2_Display/lt154_c7 ;
  wire \u2_Display/lt154_c8 ;
  wire \u2_Display/lt154_c9 ;
  wire \u2_Display/lt155_c0 ;
  wire \u2_Display/lt155_c1 ;
  wire \u2_Display/lt155_c10 ;
  wire \u2_Display/lt155_c11 ;
  wire \u2_Display/lt155_c12 ;
  wire \u2_Display/lt155_c13 ;
  wire \u2_Display/lt155_c14 ;
  wire \u2_Display/lt155_c15 ;
  wire \u2_Display/lt155_c16 ;
  wire \u2_Display/lt155_c17 ;
  wire \u2_Display/lt155_c18 ;
  wire \u2_Display/lt155_c19 ;
  wire \u2_Display/lt155_c2 ;
  wire \u2_Display/lt155_c20 ;
  wire \u2_Display/lt155_c21 ;
  wire \u2_Display/lt155_c22 ;
  wire \u2_Display/lt155_c23 ;
  wire \u2_Display/lt155_c24 ;
  wire \u2_Display/lt155_c25 ;
  wire \u2_Display/lt155_c26 ;
  wire \u2_Display/lt155_c27 ;
  wire \u2_Display/lt155_c28 ;
  wire \u2_Display/lt155_c29 ;
  wire \u2_Display/lt155_c3 ;
  wire \u2_Display/lt155_c30 ;
  wire \u2_Display/lt155_c31 ;
  wire \u2_Display/lt155_c32 ;
  wire \u2_Display/lt155_c4 ;
  wire \u2_Display/lt155_c5 ;
  wire \u2_Display/lt155_c6 ;
  wire \u2_Display/lt155_c7 ;
  wire \u2_Display/lt155_c8 ;
  wire \u2_Display/lt155_c9 ;
  wire \u2_Display/lt156_c0 ;
  wire \u2_Display/lt156_c1 ;
  wire \u2_Display/lt156_c10 ;
  wire \u2_Display/lt156_c11 ;
  wire \u2_Display/lt156_c12 ;
  wire \u2_Display/lt156_c13 ;
  wire \u2_Display/lt156_c14 ;
  wire \u2_Display/lt156_c15 ;
  wire \u2_Display/lt156_c16 ;
  wire \u2_Display/lt156_c17 ;
  wire \u2_Display/lt156_c18 ;
  wire \u2_Display/lt156_c19 ;
  wire \u2_Display/lt156_c2 ;
  wire \u2_Display/lt156_c20 ;
  wire \u2_Display/lt156_c21 ;
  wire \u2_Display/lt156_c22 ;
  wire \u2_Display/lt156_c23 ;
  wire \u2_Display/lt156_c24 ;
  wire \u2_Display/lt156_c25 ;
  wire \u2_Display/lt156_c26 ;
  wire \u2_Display/lt156_c27 ;
  wire \u2_Display/lt156_c28 ;
  wire \u2_Display/lt156_c29 ;
  wire \u2_Display/lt156_c3 ;
  wire \u2_Display/lt156_c30 ;
  wire \u2_Display/lt156_c31 ;
  wire \u2_Display/lt156_c32 ;
  wire \u2_Display/lt156_c4 ;
  wire \u2_Display/lt156_c5 ;
  wire \u2_Display/lt156_c6 ;
  wire \u2_Display/lt156_c7 ;
  wire \u2_Display/lt156_c8 ;
  wire \u2_Display/lt156_c9 ;
  wire \u2_Display/lt157_c0 ;
  wire \u2_Display/lt157_c1 ;
  wire \u2_Display/lt157_c10 ;
  wire \u2_Display/lt157_c11 ;
  wire \u2_Display/lt157_c12 ;
  wire \u2_Display/lt157_c13 ;
  wire \u2_Display/lt157_c14 ;
  wire \u2_Display/lt157_c15 ;
  wire \u2_Display/lt157_c16 ;
  wire \u2_Display/lt157_c17 ;
  wire \u2_Display/lt157_c18 ;
  wire \u2_Display/lt157_c19 ;
  wire \u2_Display/lt157_c2 ;
  wire \u2_Display/lt157_c20 ;
  wire \u2_Display/lt157_c21 ;
  wire \u2_Display/lt157_c22 ;
  wire \u2_Display/lt157_c23 ;
  wire \u2_Display/lt157_c24 ;
  wire \u2_Display/lt157_c25 ;
  wire \u2_Display/lt157_c26 ;
  wire \u2_Display/lt157_c27 ;
  wire \u2_Display/lt157_c28 ;
  wire \u2_Display/lt157_c29 ;
  wire \u2_Display/lt157_c3 ;
  wire \u2_Display/lt157_c30 ;
  wire \u2_Display/lt157_c31 ;
  wire \u2_Display/lt157_c32 ;
  wire \u2_Display/lt157_c4 ;
  wire \u2_Display/lt157_c5 ;
  wire \u2_Display/lt157_c6 ;
  wire \u2_Display/lt157_c7 ;
  wire \u2_Display/lt157_c8 ;
  wire \u2_Display/lt157_c9 ;
  wire \u2_Display/lt158_c0 ;
  wire \u2_Display/lt158_c1 ;
  wire \u2_Display/lt158_c10 ;
  wire \u2_Display/lt158_c11 ;
  wire \u2_Display/lt158_c12 ;
  wire \u2_Display/lt158_c13 ;
  wire \u2_Display/lt158_c14 ;
  wire \u2_Display/lt158_c15 ;
  wire \u2_Display/lt158_c16 ;
  wire \u2_Display/lt158_c17 ;
  wire \u2_Display/lt158_c18 ;
  wire \u2_Display/lt158_c19 ;
  wire \u2_Display/lt158_c2 ;
  wire \u2_Display/lt158_c20 ;
  wire \u2_Display/lt158_c21 ;
  wire \u2_Display/lt158_c22 ;
  wire \u2_Display/lt158_c23 ;
  wire \u2_Display/lt158_c24 ;
  wire \u2_Display/lt158_c25 ;
  wire \u2_Display/lt158_c26 ;
  wire \u2_Display/lt158_c27 ;
  wire \u2_Display/lt158_c28 ;
  wire \u2_Display/lt158_c29 ;
  wire \u2_Display/lt158_c3 ;
  wire \u2_Display/lt158_c30 ;
  wire \u2_Display/lt158_c31 ;
  wire \u2_Display/lt158_c32 ;
  wire \u2_Display/lt158_c4 ;
  wire \u2_Display/lt158_c5 ;
  wire \u2_Display/lt158_c6 ;
  wire \u2_Display/lt158_c7 ;
  wire \u2_Display/lt158_c8 ;
  wire \u2_Display/lt158_c9 ;
  wire \u2_Display/lt159_c0 ;
  wire \u2_Display/lt159_c1 ;
  wire \u2_Display/lt159_c10 ;
  wire \u2_Display/lt159_c11 ;
  wire \u2_Display/lt159_c12 ;
  wire \u2_Display/lt159_c13 ;
  wire \u2_Display/lt159_c14 ;
  wire \u2_Display/lt159_c15 ;
  wire \u2_Display/lt159_c16 ;
  wire \u2_Display/lt159_c17 ;
  wire \u2_Display/lt159_c18 ;
  wire \u2_Display/lt159_c19 ;
  wire \u2_Display/lt159_c2 ;
  wire \u2_Display/lt159_c20 ;
  wire \u2_Display/lt159_c21 ;
  wire \u2_Display/lt159_c22 ;
  wire \u2_Display/lt159_c23 ;
  wire \u2_Display/lt159_c24 ;
  wire \u2_Display/lt159_c25 ;
  wire \u2_Display/lt159_c26 ;
  wire \u2_Display/lt159_c27 ;
  wire \u2_Display/lt159_c28 ;
  wire \u2_Display/lt159_c29 ;
  wire \u2_Display/lt159_c3 ;
  wire \u2_Display/lt159_c30 ;
  wire \u2_Display/lt159_c31 ;
  wire \u2_Display/lt159_c32 ;
  wire \u2_Display/lt159_c4 ;
  wire \u2_Display/lt159_c5 ;
  wire \u2_Display/lt159_c6 ;
  wire \u2_Display/lt159_c7 ;
  wire \u2_Display/lt159_c8 ;
  wire \u2_Display/lt159_c9 ;
  wire \u2_Display/lt160_c0 ;
  wire \u2_Display/lt160_c1 ;
  wire \u2_Display/lt160_c10 ;
  wire \u2_Display/lt160_c11 ;
  wire \u2_Display/lt160_c12 ;
  wire \u2_Display/lt160_c13 ;
  wire \u2_Display/lt160_c14 ;
  wire \u2_Display/lt160_c15 ;
  wire \u2_Display/lt160_c16 ;
  wire \u2_Display/lt160_c17 ;
  wire \u2_Display/lt160_c18 ;
  wire \u2_Display/lt160_c19 ;
  wire \u2_Display/lt160_c2 ;
  wire \u2_Display/lt160_c20 ;
  wire \u2_Display/lt160_c21 ;
  wire \u2_Display/lt160_c22 ;
  wire \u2_Display/lt160_c23 ;
  wire \u2_Display/lt160_c24 ;
  wire \u2_Display/lt160_c25 ;
  wire \u2_Display/lt160_c26 ;
  wire \u2_Display/lt160_c27 ;
  wire \u2_Display/lt160_c28 ;
  wire \u2_Display/lt160_c29 ;
  wire \u2_Display/lt160_c3 ;
  wire \u2_Display/lt160_c30 ;
  wire \u2_Display/lt160_c31 ;
  wire \u2_Display/lt160_c32 ;
  wire \u2_Display/lt160_c4 ;
  wire \u2_Display/lt160_c5 ;
  wire \u2_Display/lt160_c6 ;
  wire \u2_Display/lt160_c7 ;
  wire \u2_Display/lt160_c8 ;
  wire \u2_Display/lt160_c9 ;
  wire \u2_Display/lt161_c0 ;
  wire \u2_Display/lt161_c1 ;
  wire \u2_Display/lt161_c10 ;
  wire \u2_Display/lt161_c11 ;
  wire \u2_Display/lt161_c12 ;
  wire \u2_Display/lt161_c13 ;
  wire \u2_Display/lt161_c14 ;
  wire \u2_Display/lt161_c15 ;
  wire \u2_Display/lt161_c16 ;
  wire \u2_Display/lt161_c17 ;
  wire \u2_Display/lt161_c18 ;
  wire \u2_Display/lt161_c19 ;
  wire \u2_Display/lt161_c2 ;
  wire \u2_Display/lt161_c20 ;
  wire \u2_Display/lt161_c21 ;
  wire \u2_Display/lt161_c22 ;
  wire \u2_Display/lt161_c23 ;
  wire \u2_Display/lt161_c24 ;
  wire \u2_Display/lt161_c25 ;
  wire \u2_Display/lt161_c26 ;
  wire \u2_Display/lt161_c27 ;
  wire \u2_Display/lt161_c28 ;
  wire \u2_Display/lt161_c29 ;
  wire \u2_Display/lt161_c3 ;
  wire \u2_Display/lt161_c30 ;
  wire \u2_Display/lt161_c31 ;
  wire \u2_Display/lt161_c32 ;
  wire \u2_Display/lt161_c4 ;
  wire \u2_Display/lt161_c5 ;
  wire \u2_Display/lt161_c6 ;
  wire \u2_Display/lt161_c7 ;
  wire \u2_Display/lt161_c8 ;
  wire \u2_Display/lt161_c9 ;
  wire \u2_Display/lt162_c0 ;
  wire \u2_Display/lt162_c1 ;
  wire \u2_Display/lt162_c10 ;
  wire \u2_Display/lt162_c11 ;
  wire \u2_Display/lt162_c12 ;
  wire \u2_Display/lt162_c13 ;
  wire \u2_Display/lt162_c14 ;
  wire \u2_Display/lt162_c15 ;
  wire \u2_Display/lt162_c16 ;
  wire \u2_Display/lt162_c17 ;
  wire \u2_Display/lt162_c18 ;
  wire \u2_Display/lt162_c19 ;
  wire \u2_Display/lt162_c2 ;
  wire \u2_Display/lt162_c20 ;
  wire \u2_Display/lt162_c21 ;
  wire \u2_Display/lt162_c22 ;
  wire \u2_Display/lt162_c23 ;
  wire \u2_Display/lt162_c24 ;
  wire \u2_Display/lt162_c25 ;
  wire \u2_Display/lt162_c26 ;
  wire \u2_Display/lt162_c27 ;
  wire \u2_Display/lt162_c28 ;
  wire \u2_Display/lt162_c29 ;
  wire \u2_Display/lt162_c3 ;
  wire \u2_Display/lt162_c30 ;
  wire \u2_Display/lt162_c31 ;
  wire \u2_Display/lt162_c32 ;
  wire \u2_Display/lt162_c4 ;
  wire \u2_Display/lt162_c5 ;
  wire \u2_Display/lt162_c6 ;
  wire \u2_Display/lt162_c7 ;
  wire \u2_Display/lt162_c8 ;
  wire \u2_Display/lt162_c9 ;
  wire \u2_Display/lt163_c0 ;
  wire \u2_Display/lt163_c1 ;
  wire \u2_Display/lt163_c10 ;
  wire \u2_Display/lt163_c11 ;
  wire \u2_Display/lt163_c12 ;
  wire \u2_Display/lt163_c13 ;
  wire \u2_Display/lt163_c14 ;
  wire \u2_Display/lt163_c15 ;
  wire \u2_Display/lt163_c16 ;
  wire \u2_Display/lt163_c17 ;
  wire \u2_Display/lt163_c18 ;
  wire \u2_Display/lt163_c19 ;
  wire \u2_Display/lt163_c2 ;
  wire \u2_Display/lt163_c20 ;
  wire \u2_Display/lt163_c21 ;
  wire \u2_Display/lt163_c22 ;
  wire \u2_Display/lt163_c23 ;
  wire \u2_Display/lt163_c24 ;
  wire \u2_Display/lt163_c25 ;
  wire \u2_Display/lt163_c26 ;
  wire \u2_Display/lt163_c27 ;
  wire \u2_Display/lt163_c28 ;
  wire \u2_Display/lt163_c29 ;
  wire \u2_Display/lt163_c3 ;
  wire \u2_Display/lt163_c30 ;
  wire \u2_Display/lt163_c31 ;
  wire \u2_Display/lt163_c32 ;
  wire \u2_Display/lt163_c4 ;
  wire \u2_Display/lt163_c5 ;
  wire \u2_Display/lt163_c6 ;
  wire \u2_Display/lt163_c7 ;
  wire \u2_Display/lt163_c8 ;
  wire \u2_Display/lt163_c9 ;
  wire \u2_Display/lt164_c0 ;
  wire \u2_Display/lt164_c1 ;
  wire \u2_Display/lt164_c10 ;
  wire \u2_Display/lt164_c11 ;
  wire \u2_Display/lt164_c12 ;
  wire \u2_Display/lt164_c13 ;
  wire \u2_Display/lt164_c14 ;
  wire \u2_Display/lt164_c15 ;
  wire \u2_Display/lt164_c16 ;
  wire \u2_Display/lt164_c17 ;
  wire \u2_Display/lt164_c18 ;
  wire \u2_Display/lt164_c19 ;
  wire \u2_Display/lt164_c2 ;
  wire \u2_Display/lt164_c20 ;
  wire \u2_Display/lt164_c21 ;
  wire \u2_Display/lt164_c22 ;
  wire \u2_Display/lt164_c23 ;
  wire \u2_Display/lt164_c24 ;
  wire \u2_Display/lt164_c25 ;
  wire \u2_Display/lt164_c26 ;
  wire \u2_Display/lt164_c27 ;
  wire \u2_Display/lt164_c28 ;
  wire \u2_Display/lt164_c29 ;
  wire \u2_Display/lt164_c3 ;
  wire \u2_Display/lt164_c30 ;
  wire \u2_Display/lt164_c31 ;
  wire \u2_Display/lt164_c32 ;
  wire \u2_Display/lt164_c4 ;
  wire \u2_Display/lt164_c5 ;
  wire \u2_Display/lt164_c6 ;
  wire \u2_Display/lt164_c7 ;
  wire \u2_Display/lt164_c8 ;
  wire \u2_Display/lt164_c9 ;
  wire \u2_Display/lt165_c0 ;
  wire \u2_Display/lt165_c1 ;
  wire \u2_Display/lt165_c10 ;
  wire \u2_Display/lt165_c11 ;
  wire \u2_Display/lt165_c12 ;
  wire \u2_Display/lt165_c13 ;
  wire \u2_Display/lt165_c14 ;
  wire \u2_Display/lt165_c15 ;
  wire \u2_Display/lt165_c16 ;
  wire \u2_Display/lt165_c17 ;
  wire \u2_Display/lt165_c18 ;
  wire \u2_Display/lt165_c19 ;
  wire \u2_Display/lt165_c2 ;
  wire \u2_Display/lt165_c20 ;
  wire \u2_Display/lt165_c21 ;
  wire \u2_Display/lt165_c22 ;
  wire \u2_Display/lt165_c23 ;
  wire \u2_Display/lt165_c24 ;
  wire \u2_Display/lt165_c25 ;
  wire \u2_Display/lt165_c26 ;
  wire \u2_Display/lt165_c27 ;
  wire \u2_Display/lt165_c28 ;
  wire \u2_Display/lt165_c29 ;
  wire \u2_Display/lt165_c3 ;
  wire \u2_Display/lt165_c30 ;
  wire \u2_Display/lt165_c31 ;
  wire \u2_Display/lt165_c32 ;
  wire \u2_Display/lt165_c4 ;
  wire \u2_Display/lt165_c5 ;
  wire \u2_Display/lt165_c6 ;
  wire \u2_Display/lt165_c7 ;
  wire \u2_Display/lt165_c8 ;
  wire \u2_Display/lt165_c9 ;
  wire \u2_Display/lt166_c0 ;
  wire \u2_Display/lt166_c1 ;
  wire \u2_Display/lt166_c10 ;
  wire \u2_Display/lt166_c11 ;
  wire \u2_Display/lt166_c12 ;
  wire \u2_Display/lt166_c13 ;
  wire \u2_Display/lt166_c14 ;
  wire \u2_Display/lt166_c15 ;
  wire \u2_Display/lt166_c16 ;
  wire \u2_Display/lt166_c17 ;
  wire \u2_Display/lt166_c18 ;
  wire \u2_Display/lt166_c19 ;
  wire \u2_Display/lt166_c2 ;
  wire \u2_Display/lt166_c20 ;
  wire \u2_Display/lt166_c21 ;
  wire \u2_Display/lt166_c22 ;
  wire \u2_Display/lt166_c23 ;
  wire \u2_Display/lt166_c24 ;
  wire \u2_Display/lt166_c25 ;
  wire \u2_Display/lt166_c26 ;
  wire \u2_Display/lt166_c27 ;
  wire \u2_Display/lt166_c28 ;
  wire \u2_Display/lt166_c29 ;
  wire \u2_Display/lt166_c3 ;
  wire \u2_Display/lt166_c30 ;
  wire \u2_Display/lt166_c31 ;
  wire \u2_Display/lt166_c32 ;
  wire \u2_Display/lt166_c4 ;
  wire \u2_Display/lt166_c5 ;
  wire \u2_Display/lt166_c6 ;
  wire \u2_Display/lt166_c7 ;
  wire \u2_Display/lt166_c8 ;
  wire \u2_Display/lt166_c9 ;
  wire \u2_Display/lt167_c0 ;
  wire \u2_Display/lt167_c1 ;
  wire \u2_Display/lt167_c10 ;
  wire \u2_Display/lt167_c11 ;
  wire \u2_Display/lt167_c12 ;
  wire \u2_Display/lt167_c13 ;
  wire \u2_Display/lt167_c14 ;
  wire \u2_Display/lt167_c15 ;
  wire \u2_Display/lt167_c16 ;
  wire \u2_Display/lt167_c17 ;
  wire \u2_Display/lt167_c18 ;
  wire \u2_Display/lt167_c19 ;
  wire \u2_Display/lt167_c2 ;
  wire \u2_Display/lt167_c20 ;
  wire \u2_Display/lt167_c21 ;
  wire \u2_Display/lt167_c22 ;
  wire \u2_Display/lt167_c23 ;
  wire \u2_Display/lt167_c24 ;
  wire \u2_Display/lt167_c25 ;
  wire \u2_Display/lt167_c26 ;
  wire \u2_Display/lt167_c27 ;
  wire \u2_Display/lt167_c28 ;
  wire \u2_Display/lt167_c29 ;
  wire \u2_Display/lt167_c3 ;
  wire \u2_Display/lt167_c30 ;
  wire \u2_Display/lt167_c31 ;
  wire \u2_Display/lt167_c32 ;
  wire \u2_Display/lt167_c4 ;
  wire \u2_Display/lt167_c5 ;
  wire \u2_Display/lt167_c6 ;
  wire \u2_Display/lt167_c7 ;
  wire \u2_Display/lt167_c8 ;
  wire \u2_Display/lt167_c9 ;
  wire \u2_Display/lt168_c0 ;
  wire \u2_Display/lt168_c1 ;
  wire \u2_Display/lt168_c10 ;
  wire \u2_Display/lt168_c11 ;
  wire \u2_Display/lt168_c12 ;
  wire \u2_Display/lt168_c13 ;
  wire \u2_Display/lt168_c14 ;
  wire \u2_Display/lt168_c15 ;
  wire \u2_Display/lt168_c16 ;
  wire \u2_Display/lt168_c17 ;
  wire \u2_Display/lt168_c18 ;
  wire \u2_Display/lt168_c19 ;
  wire \u2_Display/lt168_c2 ;
  wire \u2_Display/lt168_c20 ;
  wire \u2_Display/lt168_c21 ;
  wire \u2_Display/lt168_c22 ;
  wire \u2_Display/lt168_c23 ;
  wire \u2_Display/lt168_c24 ;
  wire \u2_Display/lt168_c25 ;
  wire \u2_Display/lt168_c26 ;
  wire \u2_Display/lt168_c27 ;
  wire \u2_Display/lt168_c28 ;
  wire \u2_Display/lt168_c29 ;
  wire \u2_Display/lt168_c3 ;
  wire \u2_Display/lt168_c30 ;
  wire \u2_Display/lt168_c31 ;
  wire \u2_Display/lt168_c32 ;
  wire \u2_Display/lt168_c4 ;
  wire \u2_Display/lt168_c5 ;
  wire \u2_Display/lt168_c6 ;
  wire \u2_Display/lt168_c7 ;
  wire \u2_Display/lt168_c8 ;
  wire \u2_Display/lt168_c9 ;
  wire \u2_Display/lt169_c0 ;
  wire \u2_Display/lt169_c1 ;
  wire \u2_Display/lt169_c10 ;
  wire \u2_Display/lt169_c11 ;
  wire \u2_Display/lt169_c12 ;
  wire \u2_Display/lt169_c13 ;
  wire \u2_Display/lt169_c14 ;
  wire \u2_Display/lt169_c15 ;
  wire \u2_Display/lt169_c16 ;
  wire \u2_Display/lt169_c17 ;
  wire \u2_Display/lt169_c18 ;
  wire \u2_Display/lt169_c19 ;
  wire \u2_Display/lt169_c2 ;
  wire \u2_Display/lt169_c20 ;
  wire \u2_Display/lt169_c21 ;
  wire \u2_Display/lt169_c22 ;
  wire \u2_Display/lt169_c23 ;
  wire \u2_Display/lt169_c24 ;
  wire \u2_Display/lt169_c25 ;
  wire \u2_Display/lt169_c26 ;
  wire \u2_Display/lt169_c27 ;
  wire \u2_Display/lt169_c28 ;
  wire \u2_Display/lt169_c29 ;
  wire \u2_Display/lt169_c3 ;
  wire \u2_Display/lt169_c30 ;
  wire \u2_Display/lt169_c31 ;
  wire \u2_Display/lt169_c32 ;
  wire \u2_Display/lt169_c4 ;
  wire \u2_Display/lt169_c5 ;
  wire \u2_Display/lt169_c6 ;
  wire \u2_Display/lt169_c7 ;
  wire \u2_Display/lt169_c8 ;
  wire \u2_Display/lt169_c9 ;
  wire \u2_Display/lt170_c0 ;
  wire \u2_Display/lt170_c1 ;
  wire \u2_Display/lt170_c10 ;
  wire \u2_Display/lt170_c11 ;
  wire \u2_Display/lt170_c12 ;
  wire \u2_Display/lt170_c13 ;
  wire \u2_Display/lt170_c14 ;
  wire \u2_Display/lt170_c15 ;
  wire \u2_Display/lt170_c16 ;
  wire \u2_Display/lt170_c17 ;
  wire \u2_Display/lt170_c18 ;
  wire \u2_Display/lt170_c19 ;
  wire \u2_Display/lt170_c2 ;
  wire \u2_Display/lt170_c20 ;
  wire \u2_Display/lt170_c21 ;
  wire \u2_Display/lt170_c22 ;
  wire \u2_Display/lt170_c23 ;
  wire \u2_Display/lt170_c24 ;
  wire \u2_Display/lt170_c25 ;
  wire \u2_Display/lt170_c26 ;
  wire \u2_Display/lt170_c27 ;
  wire \u2_Display/lt170_c28 ;
  wire \u2_Display/lt170_c29 ;
  wire \u2_Display/lt170_c3 ;
  wire \u2_Display/lt170_c30 ;
  wire \u2_Display/lt170_c31 ;
  wire \u2_Display/lt170_c32 ;
  wire \u2_Display/lt170_c4 ;
  wire \u2_Display/lt170_c5 ;
  wire \u2_Display/lt170_c6 ;
  wire \u2_Display/lt170_c7 ;
  wire \u2_Display/lt170_c8 ;
  wire \u2_Display/lt170_c9 ;
  wire \u2_Display/lt171_c0 ;
  wire \u2_Display/lt171_c1 ;
  wire \u2_Display/lt171_c10 ;
  wire \u2_Display/lt171_c11 ;
  wire \u2_Display/lt171_c12 ;
  wire \u2_Display/lt171_c13 ;
  wire \u2_Display/lt171_c14 ;
  wire \u2_Display/lt171_c15 ;
  wire \u2_Display/lt171_c16 ;
  wire \u2_Display/lt171_c17 ;
  wire \u2_Display/lt171_c18 ;
  wire \u2_Display/lt171_c19 ;
  wire \u2_Display/lt171_c2 ;
  wire \u2_Display/lt171_c20 ;
  wire \u2_Display/lt171_c21 ;
  wire \u2_Display/lt171_c22 ;
  wire \u2_Display/lt171_c23 ;
  wire \u2_Display/lt171_c24 ;
  wire \u2_Display/lt171_c25 ;
  wire \u2_Display/lt171_c26 ;
  wire \u2_Display/lt171_c27 ;
  wire \u2_Display/lt171_c28 ;
  wire \u2_Display/lt171_c29 ;
  wire \u2_Display/lt171_c3 ;
  wire \u2_Display/lt171_c30 ;
  wire \u2_Display/lt171_c31 ;
  wire \u2_Display/lt171_c32 ;
  wire \u2_Display/lt171_c4 ;
  wire \u2_Display/lt171_c5 ;
  wire \u2_Display/lt171_c6 ;
  wire \u2_Display/lt171_c7 ;
  wire \u2_Display/lt171_c8 ;
  wire \u2_Display/lt171_c9 ;
  wire \u2_Display/lt172_c0 ;
  wire \u2_Display/lt172_c1 ;
  wire \u2_Display/lt172_c10 ;
  wire \u2_Display/lt172_c11 ;
  wire \u2_Display/lt172_c12 ;
  wire \u2_Display/lt172_c13 ;
  wire \u2_Display/lt172_c14 ;
  wire \u2_Display/lt172_c15 ;
  wire \u2_Display/lt172_c16 ;
  wire \u2_Display/lt172_c17 ;
  wire \u2_Display/lt172_c18 ;
  wire \u2_Display/lt172_c19 ;
  wire \u2_Display/lt172_c2 ;
  wire \u2_Display/lt172_c20 ;
  wire \u2_Display/lt172_c21 ;
  wire \u2_Display/lt172_c22 ;
  wire \u2_Display/lt172_c23 ;
  wire \u2_Display/lt172_c24 ;
  wire \u2_Display/lt172_c25 ;
  wire \u2_Display/lt172_c26 ;
  wire \u2_Display/lt172_c27 ;
  wire \u2_Display/lt172_c28 ;
  wire \u2_Display/lt172_c29 ;
  wire \u2_Display/lt172_c3 ;
  wire \u2_Display/lt172_c30 ;
  wire \u2_Display/lt172_c31 ;
  wire \u2_Display/lt172_c32 ;
  wire \u2_Display/lt172_c4 ;
  wire \u2_Display/lt172_c5 ;
  wire \u2_Display/lt172_c6 ;
  wire \u2_Display/lt172_c7 ;
  wire \u2_Display/lt172_c8 ;
  wire \u2_Display/lt172_c9 ;
  wire \u2_Display/lt173_c0 ;
  wire \u2_Display/lt173_c1 ;
  wire \u2_Display/lt173_c10 ;
  wire \u2_Display/lt173_c11 ;
  wire \u2_Display/lt173_c12 ;
  wire \u2_Display/lt173_c13 ;
  wire \u2_Display/lt173_c14 ;
  wire \u2_Display/lt173_c15 ;
  wire \u2_Display/lt173_c16 ;
  wire \u2_Display/lt173_c17 ;
  wire \u2_Display/lt173_c18 ;
  wire \u2_Display/lt173_c19 ;
  wire \u2_Display/lt173_c2 ;
  wire \u2_Display/lt173_c20 ;
  wire \u2_Display/lt173_c21 ;
  wire \u2_Display/lt173_c22 ;
  wire \u2_Display/lt173_c23 ;
  wire \u2_Display/lt173_c24 ;
  wire \u2_Display/lt173_c25 ;
  wire \u2_Display/lt173_c26 ;
  wire \u2_Display/lt173_c27 ;
  wire \u2_Display/lt173_c28 ;
  wire \u2_Display/lt173_c29 ;
  wire \u2_Display/lt173_c3 ;
  wire \u2_Display/lt173_c30 ;
  wire \u2_Display/lt173_c31 ;
  wire \u2_Display/lt173_c32 ;
  wire \u2_Display/lt173_c4 ;
  wire \u2_Display/lt173_c5 ;
  wire \u2_Display/lt173_c6 ;
  wire \u2_Display/lt173_c7 ;
  wire \u2_Display/lt173_c8 ;
  wire \u2_Display/lt173_c9 ;
  wire \u2_Display/lt174_c0 ;
  wire \u2_Display/lt174_c1 ;
  wire \u2_Display/lt174_c10 ;
  wire \u2_Display/lt174_c11 ;
  wire \u2_Display/lt174_c12 ;
  wire \u2_Display/lt174_c13 ;
  wire \u2_Display/lt174_c14 ;
  wire \u2_Display/lt174_c15 ;
  wire \u2_Display/lt174_c16 ;
  wire \u2_Display/lt174_c17 ;
  wire \u2_Display/lt174_c18 ;
  wire \u2_Display/lt174_c19 ;
  wire \u2_Display/lt174_c2 ;
  wire \u2_Display/lt174_c20 ;
  wire \u2_Display/lt174_c21 ;
  wire \u2_Display/lt174_c22 ;
  wire \u2_Display/lt174_c23 ;
  wire \u2_Display/lt174_c24 ;
  wire \u2_Display/lt174_c25 ;
  wire \u2_Display/lt174_c26 ;
  wire \u2_Display/lt174_c27 ;
  wire \u2_Display/lt174_c28 ;
  wire \u2_Display/lt174_c29 ;
  wire \u2_Display/lt174_c3 ;
  wire \u2_Display/lt174_c30 ;
  wire \u2_Display/lt174_c31 ;
  wire \u2_Display/lt174_c32 ;
  wire \u2_Display/lt174_c4 ;
  wire \u2_Display/lt174_c5 ;
  wire \u2_Display/lt174_c6 ;
  wire \u2_Display/lt174_c7 ;
  wire \u2_Display/lt174_c8 ;
  wire \u2_Display/lt174_c9 ;
  wire \u2_Display/lt175_c0 ;
  wire \u2_Display/lt175_c1 ;
  wire \u2_Display/lt175_c10 ;
  wire \u2_Display/lt175_c11 ;
  wire \u2_Display/lt175_c12 ;
  wire \u2_Display/lt175_c13 ;
  wire \u2_Display/lt175_c14 ;
  wire \u2_Display/lt175_c15 ;
  wire \u2_Display/lt175_c16 ;
  wire \u2_Display/lt175_c17 ;
  wire \u2_Display/lt175_c18 ;
  wire \u2_Display/lt175_c19 ;
  wire \u2_Display/lt175_c2 ;
  wire \u2_Display/lt175_c20 ;
  wire \u2_Display/lt175_c21 ;
  wire \u2_Display/lt175_c22 ;
  wire \u2_Display/lt175_c23 ;
  wire \u2_Display/lt175_c24 ;
  wire \u2_Display/lt175_c25 ;
  wire \u2_Display/lt175_c26 ;
  wire \u2_Display/lt175_c27 ;
  wire \u2_Display/lt175_c28 ;
  wire \u2_Display/lt175_c29 ;
  wire \u2_Display/lt175_c3 ;
  wire \u2_Display/lt175_c30 ;
  wire \u2_Display/lt175_c31 ;
  wire \u2_Display/lt175_c32 ;
  wire \u2_Display/lt175_c4 ;
  wire \u2_Display/lt175_c5 ;
  wire \u2_Display/lt175_c6 ;
  wire \u2_Display/lt175_c7 ;
  wire \u2_Display/lt175_c8 ;
  wire \u2_Display/lt175_c9 ;
  wire \u2_Display/lt176_c0 ;
  wire \u2_Display/lt176_c1 ;
  wire \u2_Display/lt176_c10 ;
  wire \u2_Display/lt176_c11 ;
  wire \u2_Display/lt176_c12 ;
  wire \u2_Display/lt176_c13 ;
  wire \u2_Display/lt176_c14 ;
  wire \u2_Display/lt176_c15 ;
  wire \u2_Display/lt176_c16 ;
  wire \u2_Display/lt176_c17 ;
  wire \u2_Display/lt176_c18 ;
  wire \u2_Display/lt176_c19 ;
  wire \u2_Display/lt176_c2 ;
  wire \u2_Display/lt176_c20 ;
  wire \u2_Display/lt176_c21 ;
  wire \u2_Display/lt176_c22 ;
  wire \u2_Display/lt176_c23 ;
  wire \u2_Display/lt176_c24 ;
  wire \u2_Display/lt176_c25 ;
  wire \u2_Display/lt176_c26 ;
  wire \u2_Display/lt176_c27 ;
  wire \u2_Display/lt176_c28 ;
  wire \u2_Display/lt176_c29 ;
  wire \u2_Display/lt176_c3 ;
  wire \u2_Display/lt176_c30 ;
  wire \u2_Display/lt176_c31 ;
  wire \u2_Display/lt176_c32 ;
  wire \u2_Display/lt176_c4 ;
  wire \u2_Display/lt176_c5 ;
  wire \u2_Display/lt176_c6 ;
  wire \u2_Display/lt176_c7 ;
  wire \u2_Display/lt176_c8 ;
  wire \u2_Display/lt176_c9 ;
  wire \u2_Display/lt1_c0 ;
  wire \u2_Display/lt1_c1 ;
  wire \u2_Display/lt1_c10 ;
  wire \u2_Display/lt1_c11 ;
  wire \u2_Display/lt1_c12 ;
  wire \u2_Display/lt1_c2 ;
  wire \u2_Display/lt1_c3 ;
  wire \u2_Display/lt1_c4 ;
  wire \u2_Display/lt1_c5 ;
  wire \u2_Display/lt1_c6 ;
  wire \u2_Display/lt1_c7 ;
  wire \u2_Display/lt1_c8 ;
  wire \u2_Display/lt1_c9 ;
  wire \u2_Display/lt22_c0 ;
  wire \u2_Display/lt22_c1 ;
  wire \u2_Display/lt22_c10 ;
  wire \u2_Display/lt22_c11 ;
  wire \u2_Display/lt22_c12 ;
  wire \u2_Display/lt22_c13 ;
  wire \u2_Display/lt22_c14 ;
  wire \u2_Display/lt22_c15 ;
  wire \u2_Display/lt22_c16 ;
  wire \u2_Display/lt22_c17 ;
  wire \u2_Display/lt22_c18 ;
  wire \u2_Display/lt22_c19 ;
  wire \u2_Display/lt22_c2 ;
  wire \u2_Display/lt22_c20 ;
  wire \u2_Display/lt22_c21 ;
  wire \u2_Display/lt22_c22 ;
  wire \u2_Display/lt22_c23 ;
  wire \u2_Display/lt22_c24 ;
  wire \u2_Display/lt22_c25 ;
  wire \u2_Display/lt22_c26 ;
  wire \u2_Display/lt22_c27 ;
  wire \u2_Display/lt22_c28 ;
  wire \u2_Display/lt22_c29 ;
  wire \u2_Display/lt22_c3 ;
  wire \u2_Display/lt22_c30 ;
  wire \u2_Display/lt22_c31 ;
  wire \u2_Display/lt22_c32 ;
  wire \u2_Display/lt22_c4 ;
  wire \u2_Display/lt22_c5 ;
  wire \u2_Display/lt22_c6 ;
  wire \u2_Display/lt22_c7 ;
  wire \u2_Display/lt22_c8 ;
  wire \u2_Display/lt22_c9 ;
  wire \u2_Display/lt23_c0 ;
  wire \u2_Display/lt23_c1 ;
  wire \u2_Display/lt23_c10 ;
  wire \u2_Display/lt23_c11 ;
  wire \u2_Display/lt23_c12 ;
  wire \u2_Display/lt23_c13 ;
  wire \u2_Display/lt23_c14 ;
  wire \u2_Display/lt23_c15 ;
  wire \u2_Display/lt23_c16 ;
  wire \u2_Display/lt23_c17 ;
  wire \u2_Display/lt23_c18 ;
  wire \u2_Display/lt23_c19 ;
  wire \u2_Display/lt23_c2 ;
  wire \u2_Display/lt23_c20 ;
  wire \u2_Display/lt23_c21 ;
  wire \u2_Display/lt23_c22 ;
  wire \u2_Display/lt23_c23 ;
  wire \u2_Display/lt23_c24 ;
  wire \u2_Display/lt23_c25 ;
  wire \u2_Display/lt23_c26 ;
  wire \u2_Display/lt23_c27 ;
  wire \u2_Display/lt23_c28 ;
  wire \u2_Display/lt23_c29 ;
  wire \u2_Display/lt23_c3 ;
  wire \u2_Display/lt23_c30 ;
  wire \u2_Display/lt23_c31 ;
  wire \u2_Display/lt23_c32 ;
  wire \u2_Display/lt23_c4 ;
  wire \u2_Display/lt23_c5 ;
  wire \u2_Display/lt23_c6 ;
  wire \u2_Display/lt23_c7 ;
  wire \u2_Display/lt23_c8 ;
  wire \u2_Display/lt23_c9 ;
  wire \u2_Display/lt24_c0 ;
  wire \u2_Display/lt24_c1 ;
  wire \u2_Display/lt24_c10 ;
  wire \u2_Display/lt24_c11 ;
  wire \u2_Display/lt24_c12 ;
  wire \u2_Display/lt24_c13 ;
  wire \u2_Display/lt24_c14 ;
  wire \u2_Display/lt24_c15 ;
  wire \u2_Display/lt24_c16 ;
  wire \u2_Display/lt24_c17 ;
  wire \u2_Display/lt24_c18 ;
  wire \u2_Display/lt24_c19 ;
  wire \u2_Display/lt24_c2 ;
  wire \u2_Display/lt24_c20 ;
  wire \u2_Display/lt24_c21 ;
  wire \u2_Display/lt24_c22 ;
  wire \u2_Display/lt24_c23 ;
  wire \u2_Display/lt24_c24 ;
  wire \u2_Display/lt24_c25 ;
  wire \u2_Display/lt24_c26 ;
  wire \u2_Display/lt24_c27 ;
  wire \u2_Display/lt24_c28 ;
  wire \u2_Display/lt24_c29 ;
  wire \u2_Display/lt24_c3 ;
  wire \u2_Display/lt24_c30 ;
  wire \u2_Display/lt24_c31 ;
  wire \u2_Display/lt24_c32 ;
  wire \u2_Display/lt24_c4 ;
  wire \u2_Display/lt24_c5 ;
  wire \u2_Display/lt24_c6 ;
  wire \u2_Display/lt24_c7 ;
  wire \u2_Display/lt24_c8 ;
  wire \u2_Display/lt24_c9 ;
  wire \u2_Display/lt25_c0 ;
  wire \u2_Display/lt25_c1 ;
  wire \u2_Display/lt25_c10 ;
  wire \u2_Display/lt25_c11 ;
  wire \u2_Display/lt25_c12 ;
  wire \u2_Display/lt25_c13 ;
  wire \u2_Display/lt25_c14 ;
  wire \u2_Display/lt25_c15 ;
  wire \u2_Display/lt25_c16 ;
  wire \u2_Display/lt25_c17 ;
  wire \u2_Display/lt25_c18 ;
  wire \u2_Display/lt25_c19 ;
  wire \u2_Display/lt25_c2 ;
  wire \u2_Display/lt25_c20 ;
  wire \u2_Display/lt25_c21 ;
  wire \u2_Display/lt25_c22 ;
  wire \u2_Display/lt25_c23 ;
  wire \u2_Display/lt25_c24 ;
  wire \u2_Display/lt25_c25 ;
  wire \u2_Display/lt25_c26 ;
  wire \u2_Display/lt25_c27 ;
  wire \u2_Display/lt25_c28 ;
  wire \u2_Display/lt25_c29 ;
  wire \u2_Display/lt25_c3 ;
  wire \u2_Display/lt25_c30 ;
  wire \u2_Display/lt25_c31 ;
  wire \u2_Display/lt25_c32 ;
  wire \u2_Display/lt25_c4 ;
  wire \u2_Display/lt25_c5 ;
  wire \u2_Display/lt25_c6 ;
  wire \u2_Display/lt25_c7 ;
  wire \u2_Display/lt25_c8 ;
  wire \u2_Display/lt25_c9 ;
  wire \u2_Display/lt26_c0 ;
  wire \u2_Display/lt26_c1 ;
  wire \u2_Display/lt26_c10 ;
  wire \u2_Display/lt26_c11 ;
  wire \u2_Display/lt26_c12 ;
  wire \u2_Display/lt26_c13 ;
  wire \u2_Display/lt26_c14 ;
  wire \u2_Display/lt26_c15 ;
  wire \u2_Display/lt26_c16 ;
  wire \u2_Display/lt26_c17 ;
  wire \u2_Display/lt26_c18 ;
  wire \u2_Display/lt26_c19 ;
  wire \u2_Display/lt26_c2 ;
  wire \u2_Display/lt26_c20 ;
  wire \u2_Display/lt26_c21 ;
  wire \u2_Display/lt26_c22 ;
  wire \u2_Display/lt26_c23 ;
  wire \u2_Display/lt26_c24 ;
  wire \u2_Display/lt26_c25 ;
  wire \u2_Display/lt26_c26 ;
  wire \u2_Display/lt26_c27 ;
  wire \u2_Display/lt26_c28 ;
  wire \u2_Display/lt26_c29 ;
  wire \u2_Display/lt26_c3 ;
  wire \u2_Display/lt26_c30 ;
  wire \u2_Display/lt26_c31 ;
  wire \u2_Display/lt26_c32 ;
  wire \u2_Display/lt26_c4 ;
  wire \u2_Display/lt26_c5 ;
  wire \u2_Display/lt26_c6 ;
  wire \u2_Display/lt26_c7 ;
  wire \u2_Display/lt26_c8 ;
  wire \u2_Display/lt26_c9 ;
  wire \u2_Display/lt27_c0 ;
  wire \u2_Display/lt27_c1 ;
  wire \u2_Display/lt27_c10 ;
  wire \u2_Display/lt27_c11 ;
  wire \u2_Display/lt27_c12 ;
  wire \u2_Display/lt27_c13 ;
  wire \u2_Display/lt27_c14 ;
  wire \u2_Display/lt27_c15 ;
  wire \u2_Display/lt27_c16 ;
  wire \u2_Display/lt27_c17 ;
  wire \u2_Display/lt27_c18 ;
  wire \u2_Display/lt27_c19 ;
  wire \u2_Display/lt27_c2 ;
  wire \u2_Display/lt27_c20 ;
  wire \u2_Display/lt27_c21 ;
  wire \u2_Display/lt27_c22 ;
  wire \u2_Display/lt27_c23 ;
  wire \u2_Display/lt27_c24 ;
  wire \u2_Display/lt27_c25 ;
  wire \u2_Display/lt27_c26 ;
  wire \u2_Display/lt27_c27 ;
  wire \u2_Display/lt27_c28 ;
  wire \u2_Display/lt27_c29 ;
  wire \u2_Display/lt27_c3 ;
  wire \u2_Display/lt27_c30 ;
  wire \u2_Display/lt27_c31 ;
  wire \u2_Display/lt27_c32 ;
  wire \u2_Display/lt27_c4 ;
  wire \u2_Display/lt27_c5 ;
  wire \u2_Display/lt27_c6 ;
  wire \u2_Display/lt27_c7 ;
  wire \u2_Display/lt27_c8 ;
  wire \u2_Display/lt27_c9 ;
  wire \u2_Display/lt28_c0 ;
  wire \u2_Display/lt28_c1 ;
  wire \u2_Display/lt28_c10 ;
  wire \u2_Display/lt28_c11 ;
  wire \u2_Display/lt28_c12 ;
  wire \u2_Display/lt28_c13 ;
  wire \u2_Display/lt28_c14 ;
  wire \u2_Display/lt28_c15 ;
  wire \u2_Display/lt28_c16 ;
  wire \u2_Display/lt28_c17 ;
  wire \u2_Display/lt28_c18 ;
  wire \u2_Display/lt28_c19 ;
  wire \u2_Display/lt28_c2 ;
  wire \u2_Display/lt28_c20 ;
  wire \u2_Display/lt28_c21 ;
  wire \u2_Display/lt28_c22 ;
  wire \u2_Display/lt28_c23 ;
  wire \u2_Display/lt28_c24 ;
  wire \u2_Display/lt28_c25 ;
  wire \u2_Display/lt28_c26 ;
  wire \u2_Display/lt28_c27 ;
  wire \u2_Display/lt28_c28 ;
  wire \u2_Display/lt28_c29 ;
  wire \u2_Display/lt28_c3 ;
  wire \u2_Display/lt28_c30 ;
  wire \u2_Display/lt28_c31 ;
  wire \u2_Display/lt28_c32 ;
  wire \u2_Display/lt28_c4 ;
  wire \u2_Display/lt28_c5 ;
  wire \u2_Display/lt28_c6 ;
  wire \u2_Display/lt28_c7 ;
  wire \u2_Display/lt28_c8 ;
  wire \u2_Display/lt28_c9 ;
  wire \u2_Display/lt29_c0 ;
  wire \u2_Display/lt29_c1 ;
  wire \u2_Display/lt29_c10 ;
  wire \u2_Display/lt29_c11 ;
  wire \u2_Display/lt29_c12 ;
  wire \u2_Display/lt29_c13 ;
  wire \u2_Display/lt29_c14 ;
  wire \u2_Display/lt29_c15 ;
  wire \u2_Display/lt29_c16 ;
  wire \u2_Display/lt29_c17 ;
  wire \u2_Display/lt29_c18 ;
  wire \u2_Display/lt29_c19 ;
  wire \u2_Display/lt29_c2 ;
  wire \u2_Display/lt29_c20 ;
  wire \u2_Display/lt29_c21 ;
  wire \u2_Display/lt29_c22 ;
  wire \u2_Display/lt29_c23 ;
  wire \u2_Display/lt29_c24 ;
  wire \u2_Display/lt29_c25 ;
  wire \u2_Display/lt29_c26 ;
  wire \u2_Display/lt29_c27 ;
  wire \u2_Display/lt29_c28 ;
  wire \u2_Display/lt29_c29 ;
  wire \u2_Display/lt29_c3 ;
  wire \u2_Display/lt29_c30 ;
  wire \u2_Display/lt29_c31 ;
  wire \u2_Display/lt29_c32 ;
  wire \u2_Display/lt29_c4 ;
  wire \u2_Display/lt29_c5 ;
  wire \u2_Display/lt29_c6 ;
  wire \u2_Display/lt29_c7 ;
  wire \u2_Display/lt29_c8 ;
  wire \u2_Display/lt29_c9 ;
  wire \u2_Display/lt2_2_c0 ;
  wire \u2_Display/lt2_2_c1 ;
  wire \u2_Display/lt2_2_c10 ;
  wire \u2_Display/lt2_2_c11 ;
  wire \u2_Display/lt2_2_c12 ;
  wire \u2_Display/lt2_2_c2 ;
  wire \u2_Display/lt2_2_c3 ;
  wire \u2_Display/lt2_2_c4 ;
  wire \u2_Display/lt2_2_c5 ;
  wire \u2_Display/lt2_2_c6 ;
  wire \u2_Display/lt2_2_c7 ;
  wire \u2_Display/lt2_2_c8 ;
  wire \u2_Display/lt2_2_c9 ;
  wire \u2_Display/lt30_c0 ;
  wire \u2_Display/lt30_c1 ;
  wire \u2_Display/lt30_c10 ;
  wire \u2_Display/lt30_c11 ;
  wire \u2_Display/lt30_c12 ;
  wire \u2_Display/lt30_c13 ;
  wire \u2_Display/lt30_c14 ;
  wire \u2_Display/lt30_c15 ;
  wire \u2_Display/lt30_c16 ;
  wire \u2_Display/lt30_c17 ;
  wire \u2_Display/lt30_c18 ;
  wire \u2_Display/lt30_c19 ;
  wire \u2_Display/lt30_c2 ;
  wire \u2_Display/lt30_c20 ;
  wire \u2_Display/lt30_c21 ;
  wire \u2_Display/lt30_c22 ;
  wire \u2_Display/lt30_c23 ;
  wire \u2_Display/lt30_c24 ;
  wire \u2_Display/lt30_c25 ;
  wire \u2_Display/lt30_c26 ;
  wire \u2_Display/lt30_c27 ;
  wire \u2_Display/lt30_c28 ;
  wire \u2_Display/lt30_c29 ;
  wire \u2_Display/lt30_c3 ;
  wire \u2_Display/lt30_c30 ;
  wire \u2_Display/lt30_c31 ;
  wire \u2_Display/lt30_c32 ;
  wire \u2_Display/lt30_c4 ;
  wire \u2_Display/lt30_c5 ;
  wire \u2_Display/lt30_c6 ;
  wire \u2_Display/lt30_c7 ;
  wire \u2_Display/lt30_c8 ;
  wire \u2_Display/lt30_c9 ;
  wire \u2_Display/lt31_c0 ;
  wire \u2_Display/lt31_c1 ;
  wire \u2_Display/lt31_c10 ;
  wire \u2_Display/lt31_c11 ;
  wire \u2_Display/lt31_c12 ;
  wire \u2_Display/lt31_c13 ;
  wire \u2_Display/lt31_c14 ;
  wire \u2_Display/lt31_c15 ;
  wire \u2_Display/lt31_c16 ;
  wire \u2_Display/lt31_c17 ;
  wire \u2_Display/lt31_c18 ;
  wire \u2_Display/lt31_c19 ;
  wire \u2_Display/lt31_c2 ;
  wire \u2_Display/lt31_c20 ;
  wire \u2_Display/lt31_c21 ;
  wire \u2_Display/lt31_c22 ;
  wire \u2_Display/lt31_c23 ;
  wire \u2_Display/lt31_c24 ;
  wire \u2_Display/lt31_c25 ;
  wire \u2_Display/lt31_c26 ;
  wire \u2_Display/lt31_c27 ;
  wire \u2_Display/lt31_c28 ;
  wire \u2_Display/lt31_c29 ;
  wire \u2_Display/lt31_c3 ;
  wire \u2_Display/lt31_c30 ;
  wire \u2_Display/lt31_c31 ;
  wire \u2_Display/lt31_c32 ;
  wire \u2_Display/lt31_c4 ;
  wire \u2_Display/lt31_c5 ;
  wire \u2_Display/lt31_c6 ;
  wire \u2_Display/lt31_c7 ;
  wire \u2_Display/lt31_c8 ;
  wire \u2_Display/lt31_c9 ;
  wire \u2_Display/lt32_c0 ;
  wire \u2_Display/lt32_c1 ;
  wire \u2_Display/lt32_c10 ;
  wire \u2_Display/lt32_c11 ;
  wire \u2_Display/lt32_c12 ;
  wire \u2_Display/lt32_c13 ;
  wire \u2_Display/lt32_c14 ;
  wire \u2_Display/lt32_c15 ;
  wire \u2_Display/lt32_c16 ;
  wire \u2_Display/lt32_c17 ;
  wire \u2_Display/lt32_c18 ;
  wire \u2_Display/lt32_c19 ;
  wire \u2_Display/lt32_c2 ;
  wire \u2_Display/lt32_c20 ;
  wire \u2_Display/lt32_c21 ;
  wire \u2_Display/lt32_c22 ;
  wire \u2_Display/lt32_c23 ;
  wire \u2_Display/lt32_c24 ;
  wire \u2_Display/lt32_c25 ;
  wire \u2_Display/lt32_c26 ;
  wire \u2_Display/lt32_c27 ;
  wire \u2_Display/lt32_c28 ;
  wire \u2_Display/lt32_c29 ;
  wire \u2_Display/lt32_c3 ;
  wire \u2_Display/lt32_c30 ;
  wire \u2_Display/lt32_c31 ;
  wire \u2_Display/lt32_c32 ;
  wire \u2_Display/lt32_c4 ;
  wire \u2_Display/lt32_c5 ;
  wire \u2_Display/lt32_c6 ;
  wire \u2_Display/lt32_c7 ;
  wire \u2_Display/lt32_c8 ;
  wire \u2_Display/lt32_c9 ;
  wire \u2_Display/lt33_c0 ;
  wire \u2_Display/lt33_c1 ;
  wire \u2_Display/lt33_c10 ;
  wire \u2_Display/lt33_c11 ;
  wire \u2_Display/lt33_c12 ;
  wire \u2_Display/lt33_c13 ;
  wire \u2_Display/lt33_c14 ;
  wire \u2_Display/lt33_c15 ;
  wire \u2_Display/lt33_c16 ;
  wire \u2_Display/lt33_c17 ;
  wire \u2_Display/lt33_c18 ;
  wire \u2_Display/lt33_c19 ;
  wire \u2_Display/lt33_c2 ;
  wire \u2_Display/lt33_c20 ;
  wire \u2_Display/lt33_c21 ;
  wire \u2_Display/lt33_c22 ;
  wire \u2_Display/lt33_c23 ;
  wire \u2_Display/lt33_c24 ;
  wire \u2_Display/lt33_c25 ;
  wire \u2_Display/lt33_c26 ;
  wire \u2_Display/lt33_c27 ;
  wire \u2_Display/lt33_c28 ;
  wire \u2_Display/lt33_c29 ;
  wire \u2_Display/lt33_c3 ;
  wire \u2_Display/lt33_c30 ;
  wire \u2_Display/lt33_c31 ;
  wire \u2_Display/lt33_c32 ;
  wire \u2_Display/lt33_c4 ;
  wire \u2_Display/lt33_c5 ;
  wire \u2_Display/lt33_c6 ;
  wire \u2_Display/lt33_c7 ;
  wire \u2_Display/lt33_c8 ;
  wire \u2_Display/lt33_c9 ;
  wire \u2_Display/lt34_c0 ;
  wire \u2_Display/lt34_c1 ;
  wire \u2_Display/lt34_c10 ;
  wire \u2_Display/lt34_c11 ;
  wire \u2_Display/lt34_c12 ;
  wire \u2_Display/lt34_c13 ;
  wire \u2_Display/lt34_c14 ;
  wire \u2_Display/lt34_c15 ;
  wire \u2_Display/lt34_c16 ;
  wire \u2_Display/lt34_c17 ;
  wire \u2_Display/lt34_c18 ;
  wire \u2_Display/lt34_c19 ;
  wire \u2_Display/lt34_c2 ;
  wire \u2_Display/lt34_c20 ;
  wire \u2_Display/lt34_c21 ;
  wire \u2_Display/lt34_c22 ;
  wire \u2_Display/lt34_c23 ;
  wire \u2_Display/lt34_c24 ;
  wire \u2_Display/lt34_c25 ;
  wire \u2_Display/lt34_c26 ;
  wire \u2_Display/lt34_c27 ;
  wire \u2_Display/lt34_c28 ;
  wire \u2_Display/lt34_c29 ;
  wire \u2_Display/lt34_c3 ;
  wire \u2_Display/lt34_c30 ;
  wire \u2_Display/lt34_c31 ;
  wire \u2_Display/lt34_c32 ;
  wire \u2_Display/lt34_c4 ;
  wire \u2_Display/lt34_c5 ;
  wire \u2_Display/lt34_c6 ;
  wire \u2_Display/lt34_c7 ;
  wire \u2_Display/lt34_c8 ;
  wire \u2_Display/lt34_c9 ;
  wire \u2_Display/lt35_c0 ;
  wire \u2_Display/lt35_c1 ;
  wire \u2_Display/lt35_c10 ;
  wire \u2_Display/lt35_c11 ;
  wire \u2_Display/lt35_c12 ;
  wire \u2_Display/lt35_c13 ;
  wire \u2_Display/lt35_c14 ;
  wire \u2_Display/lt35_c15 ;
  wire \u2_Display/lt35_c16 ;
  wire \u2_Display/lt35_c17 ;
  wire \u2_Display/lt35_c18 ;
  wire \u2_Display/lt35_c19 ;
  wire \u2_Display/lt35_c2 ;
  wire \u2_Display/lt35_c20 ;
  wire \u2_Display/lt35_c21 ;
  wire \u2_Display/lt35_c22 ;
  wire \u2_Display/lt35_c23 ;
  wire \u2_Display/lt35_c24 ;
  wire \u2_Display/lt35_c25 ;
  wire \u2_Display/lt35_c26 ;
  wire \u2_Display/lt35_c27 ;
  wire \u2_Display/lt35_c28 ;
  wire \u2_Display/lt35_c29 ;
  wire \u2_Display/lt35_c3 ;
  wire \u2_Display/lt35_c30 ;
  wire \u2_Display/lt35_c31 ;
  wire \u2_Display/lt35_c32 ;
  wire \u2_Display/lt35_c4 ;
  wire \u2_Display/lt35_c5 ;
  wire \u2_Display/lt35_c6 ;
  wire \u2_Display/lt35_c7 ;
  wire \u2_Display/lt35_c8 ;
  wire \u2_Display/lt35_c9 ;
  wire \u2_Display/lt36_c0 ;
  wire \u2_Display/lt36_c1 ;
  wire \u2_Display/lt36_c10 ;
  wire \u2_Display/lt36_c11 ;
  wire \u2_Display/lt36_c12 ;
  wire \u2_Display/lt36_c13 ;
  wire \u2_Display/lt36_c14 ;
  wire \u2_Display/lt36_c15 ;
  wire \u2_Display/lt36_c16 ;
  wire \u2_Display/lt36_c17 ;
  wire \u2_Display/lt36_c18 ;
  wire \u2_Display/lt36_c19 ;
  wire \u2_Display/lt36_c2 ;
  wire \u2_Display/lt36_c20 ;
  wire \u2_Display/lt36_c21 ;
  wire \u2_Display/lt36_c22 ;
  wire \u2_Display/lt36_c23 ;
  wire \u2_Display/lt36_c24 ;
  wire \u2_Display/lt36_c25 ;
  wire \u2_Display/lt36_c26 ;
  wire \u2_Display/lt36_c27 ;
  wire \u2_Display/lt36_c28 ;
  wire \u2_Display/lt36_c29 ;
  wire \u2_Display/lt36_c3 ;
  wire \u2_Display/lt36_c30 ;
  wire \u2_Display/lt36_c31 ;
  wire \u2_Display/lt36_c32 ;
  wire \u2_Display/lt36_c4 ;
  wire \u2_Display/lt36_c5 ;
  wire \u2_Display/lt36_c6 ;
  wire \u2_Display/lt36_c7 ;
  wire \u2_Display/lt36_c8 ;
  wire \u2_Display/lt36_c9 ;
  wire \u2_Display/lt37_c0 ;
  wire \u2_Display/lt37_c1 ;
  wire \u2_Display/lt37_c10 ;
  wire \u2_Display/lt37_c11 ;
  wire \u2_Display/lt37_c12 ;
  wire \u2_Display/lt37_c13 ;
  wire \u2_Display/lt37_c14 ;
  wire \u2_Display/lt37_c15 ;
  wire \u2_Display/lt37_c16 ;
  wire \u2_Display/lt37_c17 ;
  wire \u2_Display/lt37_c18 ;
  wire \u2_Display/lt37_c19 ;
  wire \u2_Display/lt37_c2 ;
  wire \u2_Display/lt37_c20 ;
  wire \u2_Display/lt37_c21 ;
  wire \u2_Display/lt37_c22 ;
  wire \u2_Display/lt37_c23 ;
  wire \u2_Display/lt37_c24 ;
  wire \u2_Display/lt37_c25 ;
  wire \u2_Display/lt37_c26 ;
  wire \u2_Display/lt37_c27 ;
  wire \u2_Display/lt37_c28 ;
  wire \u2_Display/lt37_c29 ;
  wire \u2_Display/lt37_c3 ;
  wire \u2_Display/lt37_c30 ;
  wire \u2_Display/lt37_c31 ;
  wire \u2_Display/lt37_c32 ;
  wire \u2_Display/lt37_c4 ;
  wire \u2_Display/lt37_c5 ;
  wire \u2_Display/lt37_c6 ;
  wire \u2_Display/lt37_c7 ;
  wire \u2_Display/lt37_c8 ;
  wire \u2_Display/lt37_c9 ;
  wire \u2_Display/lt38_c0 ;
  wire \u2_Display/lt38_c1 ;
  wire \u2_Display/lt38_c10 ;
  wire \u2_Display/lt38_c11 ;
  wire \u2_Display/lt38_c12 ;
  wire \u2_Display/lt38_c13 ;
  wire \u2_Display/lt38_c14 ;
  wire \u2_Display/lt38_c15 ;
  wire \u2_Display/lt38_c16 ;
  wire \u2_Display/lt38_c17 ;
  wire \u2_Display/lt38_c18 ;
  wire \u2_Display/lt38_c19 ;
  wire \u2_Display/lt38_c2 ;
  wire \u2_Display/lt38_c20 ;
  wire \u2_Display/lt38_c21 ;
  wire \u2_Display/lt38_c22 ;
  wire \u2_Display/lt38_c23 ;
  wire \u2_Display/lt38_c24 ;
  wire \u2_Display/lt38_c25 ;
  wire \u2_Display/lt38_c26 ;
  wire \u2_Display/lt38_c27 ;
  wire \u2_Display/lt38_c28 ;
  wire \u2_Display/lt38_c29 ;
  wire \u2_Display/lt38_c3 ;
  wire \u2_Display/lt38_c30 ;
  wire \u2_Display/lt38_c31 ;
  wire \u2_Display/lt38_c32 ;
  wire \u2_Display/lt38_c4 ;
  wire \u2_Display/lt38_c5 ;
  wire \u2_Display/lt38_c6 ;
  wire \u2_Display/lt38_c7 ;
  wire \u2_Display/lt38_c8 ;
  wire \u2_Display/lt38_c9 ;
  wire \u2_Display/lt39_c0 ;
  wire \u2_Display/lt39_c1 ;
  wire \u2_Display/lt39_c10 ;
  wire \u2_Display/lt39_c11 ;
  wire \u2_Display/lt39_c12 ;
  wire \u2_Display/lt39_c13 ;
  wire \u2_Display/lt39_c14 ;
  wire \u2_Display/lt39_c15 ;
  wire \u2_Display/lt39_c16 ;
  wire \u2_Display/lt39_c17 ;
  wire \u2_Display/lt39_c18 ;
  wire \u2_Display/lt39_c19 ;
  wire \u2_Display/lt39_c2 ;
  wire \u2_Display/lt39_c20 ;
  wire \u2_Display/lt39_c21 ;
  wire \u2_Display/lt39_c22 ;
  wire \u2_Display/lt39_c23 ;
  wire \u2_Display/lt39_c24 ;
  wire \u2_Display/lt39_c25 ;
  wire \u2_Display/lt39_c26 ;
  wire \u2_Display/lt39_c27 ;
  wire \u2_Display/lt39_c28 ;
  wire \u2_Display/lt39_c29 ;
  wire \u2_Display/lt39_c3 ;
  wire \u2_Display/lt39_c30 ;
  wire \u2_Display/lt39_c31 ;
  wire \u2_Display/lt39_c32 ;
  wire \u2_Display/lt39_c4 ;
  wire \u2_Display/lt39_c5 ;
  wire \u2_Display/lt39_c6 ;
  wire \u2_Display/lt39_c7 ;
  wire \u2_Display/lt39_c8 ;
  wire \u2_Display/lt39_c9 ;
  wire \u2_Display/lt3_c0 ;
  wire \u2_Display/lt3_c1 ;
  wire \u2_Display/lt3_c10 ;
  wire \u2_Display/lt3_c11 ;
  wire \u2_Display/lt3_c12 ;
  wire \u2_Display/lt3_c2 ;
  wire \u2_Display/lt3_c3 ;
  wire \u2_Display/lt3_c4 ;
  wire \u2_Display/lt3_c5 ;
  wire \u2_Display/lt3_c6 ;
  wire \u2_Display/lt3_c7 ;
  wire \u2_Display/lt3_c8 ;
  wire \u2_Display/lt3_c9 ;
  wire \u2_Display/lt40_c0 ;
  wire \u2_Display/lt40_c1 ;
  wire \u2_Display/lt40_c10 ;
  wire \u2_Display/lt40_c11 ;
  wire \u2_Display/lt40_c12 ;
  wire \u2_Display/lt40_c13 ;
  wire \u2_Display/lt40_c14 ;
  wire \u2_Display/lt40_c15 ;
  wire \u2_Display/lt40_c16 ;
  wire \u2_Display/lt40_c17 ;
  wire \u2_Display/lt40_c18 ;
  wire \u2_Display/lt40_c19 ;
  wire \u2_Display/lt40_c2 ;
  wire \u2_Display/lt40_c20 ;
  wire \u2_Display/lt40_c21 ;
  wire \u2_Display/lt40_c22 ;
  wire \u2_Display/lt40_c23 ;
  wire \u2_Display/lt40_c24 ;
  wire \u2_Display/lt40_c25 ;
  wire \u2_Display/lt40_c26 ;
  wire \u2_Display/lt40_c27 ;
  wire \u2_Display/lt40_c28 ;
  wire \u2_Display/lt40_c29 ;
  wire \u2_Display/lt40_c3 ;
  wire \u2_Display/lt40_c30 ;
  wire \u2_Display/lt40_c31 ;
  wire \u2_Display/lt40_c32 ;
  wire \u2_Display/lt40_c4 ;
  wire \u2_Display/lt40_c5 ;
  wire \u2_Display/lt40_c6 ;
  wire \u2_Display/lt40_c7 ;
  wire \u2_Display/lt40_c8 ;
  wire \u2_Display/lt40_c9 ;
  wire \u2_Display/lt41_c0 ;
  wire \u2_Display/lt41_c1 ;
  wire \u2_Display/lt41_c10 ;
  wire \u2_Display/lt41_c11 ;
  wire \u2_Display/lt41_c12 ;
  wire \u2_Display/lt41_c13 ;
  wire \u2_Display/lt41_c14 ;
  wire \u2_Display/lt41_c15 ;
  wire \u2_Display/lt41_c16 ;
  wire \u2_Display/lt41_c17 ;
  wire \u2_Display/lt41_c18 ;
  wire \u2_Display/lt41_c19 ;
  wire \u2_Display/lt41_c2 ;
  wire \u2_Display/lt41_c20 ;
  wire \u2_Display/lt41_c21 ;
  wire \u2_Display/lt41_c22 ;
  wire \u2_Display/lt41_c23 ;
  wire \u2_Display/lt41_c24 ;
  wire \u2_Display/lt41_c25 ;
  wire \u2_Display/lt41_c26 ;
  wire \u2_Display/lt41_c27 ;
  wire \u2_Display/lt41_c28 ;
  wire \u2_Display/lt41_c29 ;
  wire \u2_Display/lt41_c3 ;
  wire \u2_Display/lt41_c30 ;
  wire \u2_Display/lt41_c31 ;
  wire \u2_Display/lt41_c32 ;
  wire \u2_Display/lt41_c4 ;
  wire \u2_Display/lt41_c5 ;
  wire \u2_Display/lt41_c6 ;
  wire \u2_Display/lt41_c7 ;
  wire \u2_Display/lt41_c8 ;
  wire \u2_Display/lt41_c9 ;
  wire \u2_Display/lt42_c0 ;
  wire \u2_Display/lt42_c1 ;
  wire \u2_Display/lt42_c10 ;
  wire \u2_Display/lt42_c11 ;
  wire \u2_Display/lt42_c12 ;
  wire \u2_Display/lt42_c13 ;
  wire \u2_Display/lt42_c14 ;
  wire \u2_Display/lt42_c15 ;
  wire \u2_Display/lt42_c16 ;
  wire \u2_Display/lt42_c17 ;
  wire \u2_Display/lt42_c18 ;
  wire \u2_Display/lt42_c19 ;
  wire \u2_Display/lt42_c2 ;
  wire \u2_Display/lt42_c20 ;
  wire \u2_Display/lt42_c21 ;
  wire \u2_Display/lt42_c22 ;
  wire \u2_Display/lt42_c23 ;
  wire \u2_Display/lt42_c24 ;
  wire \u2_Display/lt42_c25 ;
  wire \u2_Display/lt42_c26 ;
  wire \u2_Display/lt42_c27 ;
  wire \u2_Display/lt42_c28 ;
  wire \u2_Display/lt42_c29 ;
  wire \u2_Display/lt42_c3 ;
  wire \u2_Display/lt42_c30 ;
  wire \u2_Display/lt42_c31 ;
  wire \u2_Display/lt42_c32 ;
  wire \u2_Display/lt42_c4 ;
  wire \u2_Display/lt42_c5 ;
  wire \u2_Display/lt42_c6 ;
  wire \u2_Display/lt42_c7 ;
  wire \u2_Display/lt42_c8 ;
  wire \u2_Display/lt42_c9 ;
  wire \u2_Display/lt43_c0 ;
  wire \u2_Display/lt43_c1 ;
  wire \u2_Display/lt43_c10 ;
  wire \u2_Display/lt43_c11 ;
  wire \u2_Display/lt43_c12 ;
  wire \u2_Display/lt43_c13 ;
  wire \u2_Display/lt43_c14 ;
  wire \u2_Display/lt43_c15 ;
  wire \u2_Display/lt43_c16 ;
  wire \u2_Display/lt43_c17 ;
  wire \u2_Display/lt43_c18 ;
  wire \u2_Display/lt43_c19 ;
  wire \u2_Display/lt43_c2 ;
  wire \u2_Display/lt43_c20 ;
  wire \u2_Display/lt43_c21 ;
  wire \u2_Display/lt43_c22 ;
  wire \u2_Display/lt43_c23 ;
  wire \u2_Display/lt43_c24 ;
  wire \u2_Display/lt43_c25 ;
  wire \u2_Display/lt43_c26 ;
  wire \u2_Display/lt43_c27 ;
  wire \u2_Display/lt43_c28 ;
  wire \u2_Display/lt43_c29 ;
  wire \u2_Display/lt43_c3 ;
  wire \u2_Display/lt43_c30 ;
  wire \u2_Display/lt43_c31 ;
  wire \u2_Display/lt43_c32 ;
  wire \u2_Display/lt43_c4 ;
  wire \u2_Display/lt43_c5 ;
  wire \u2_Display/lt43_c6 ;
  wire \u2_Display/lt43_c7 ;
  wire \u2_Display/lt43_c8 ;
  wire \u2_Display/lt43_c9 ;
  wire \u2_Display/lt44_c0 ;
  wire \u2_Display/lt44_c1 ;
  wire \u2_Display/lt44_c10 ;
  wire \u2_Display/lt44_c11 ;
  wire \u2_Display/lt44_c12 ;
  wire \u2_Display/lt44_c13 ;
  wire \u2_Display/lt44_c14 ;
  wire \u2_Display/lt44_c15 ;
  wire \u2_Display/lt44_c16 ;
  wire \u2_Display/lt44_c17 ;
  wire \u2_Display/lt44_c18 ;
  wire \u2_Display/lt44_c19 ;
  wire \u2_Display/lt44_c2 ;
  wire \u2_Display/lt44_c20 ;
  wire \u2_Display/lt44_c21 ;
  wire \u2_Display/lt44_c22 ;
  wire \u2_Display/lt44_c23 ;
  wire \u2_Display/lt44_c24 ;
  wire \u2_Display/lt44_c25 ;
  wire \u2_Display/lt44_c26 ;
  wire \u2_Display/lt44_c27 ;
  wire \u2_Display/lt44_c28 ;
  wire \u2_Display/lt44_c29 ;
  wire \u2_Display/lt44_c3 ;
  wire \u2_Display/lt44_c30 ;
  wire \u2_Display/lt44_c31 ;
  wire \u2_Display/lt44_c32 ;
  wire \u2_Display/lt44_c4 ;
  wire \u2_Display/lt44_c5 ;
  wire \u2_Display/lt44_c6 ;
  wire \u2_Display/lt44_c7 ;
  wire \u2_Display/lt44_c8 ;
  wire \u2_Display/lt44_c9 ;
  wire \u2_Display/lt4_2_c0 ;
  wire \u2_Display/lt4_2_c1 ;
  wire \u2_Display/lt4_2_c10 ;
  wire \u2_Display/lt4_2_c11 ;
  wire \u2_Display/lt4_2_c12 ;
  wire \u2_Display/lt4_2_c2 ;
  wire \u2_Display/lt4_2_c3 ;
  wire \u2_Display/lt4_2_c4 ;
  wire \u2_Display/lt4_2_c5 ;
  wire \u2_Display/lt4_2_c6 ;
  wire \u2_Display/lt4_2_c7 ;
  wire \u2_Display/lt4_2_c8 ;
  wire \u2_Display/lt4_2_c9 ;
  wire \u2_Display/lt55_c0 ;
  wire \u2_Display/lt55_c1 ;
  wire \u2_Display/lt55_c10 ;
  wire \u2_Display/lt55_c11 ;
  wire \u2_Display/lt55_c12 ;
  wire \u2_Display/lt55_c13 ;
  wire \u2_Display/lt55_c14 ;
  wire \u2_Display/lt55_c15 ;
  wire \u2_Display/lt55_c16 ;
  wire \u2_Display/lt55_c17 ;
  wire \u2_Display/lt55_c18 ;
  wire \u2_Display/lt55_c19 ;
  wire \u2_Display/lt55_c2 ;
  wire \u2_Display/lt55_c20 ;
  wire \u2_Display/lt55_c21 ;
  wire \u2_Display/lt55_c22 ;
  wire \u2_Display/lt55_c23 ;
  wire \u2_Display/lt55_c24 ;
  wire \u2_Display/lt55_c25 ;
  wire \u2_Display/lt55_c26 ;
  wire \u2_Display/lt55_c27 ;
  wire \u2_Display/lt55_c28 ;
  wire \u2_Display/lt55_c29 ;
  wire \u2_Display/lt55_c3 ;
  wire \u2_Display/lt55_c30 ;
  wire \u2_Display/lt55_c31 ;
  wire \u2_Display/lt55_c32 ;
  wire \u2_Display/lt55_c4 ;
  wire \u2_Display/lt55_c5 ;
  wire \u2_Display/lt55_c6 ;
  wire \u2_Display/lt55_c7 ;
  wire \u2_Display/lt55_c8 ;
  wire \u2_Display/lt55_c9 ;
  wire \u2_Display/lt56_c0 ;
  wire \u2_Display/lt56_c1 ;
  wire \u2_Display/lt56_c10 ;
  wire \u2_Display/lt56_c11 ;
  wire \u2_Display/lt56_c12 ;
  wire \u2_Display/lt56_c13 ;
  wire \u2_Display/lt56_c14 ;
  wire \u2_Display/lt56_c15 ;
  wire \u2_Display/lt56_c16 ;
  wire \u2_Display/lt56_c17 ;
  wire \u2_Display/lt56_c18 ;
  wire \u2_Display/lt56_c19 ;
  wire \u2_Display/lt56_c2 ;
  wire \u2_Display/lt56_c20 ;
  wire \u2_Display/lt56_c21 ;
  wire \u2_Display/lt56_c22 ;
  wire \u2_Display/lt56_c23 ;
  wire \u2_Display/lt56_c24 ;
  wire \u2_Display/lt56_c25 ;
  wire \u2_Display/lt56_c26 ;
  wire \u2_Display/lt56_c27 ;
  wire \u2_Display/lt56_c28 ;
  wire \u2_Display/lt56_c29 ;
  wire \u2_Display/lt56_c3 ;
  wire \u2_Display/lt56_c30 ;
  wire \u2_Display/lt56_c31 ;
  wire \u2_Display/lt56_c32 ;
  wire \u2_Display/lt56_c4 ;
  wire \u2_Display/lt56_c5 ;
  wire \u2_Display/lt56_c6 ;
  wire \u2_Display/lt56_c7 ;
  wire \u2_Display/lt56_c8 ;
  wire \u2_Display/lt56_c9 ;
  wire \u2_Display/lt57_c0 ;
  wire \u2_Display/lt57_c1 ;
  wire \u2_Display/lt57_c10 ;
  wire \u2_Display/lt57_c11 ;
  wire \u2_Display/lt57_c12 ;
  wire \u2_Display/lt57_c13 ;
  wire \u2_Display/lt57_c14 ;
  wire \u2_Display/lt57_c15 ;
  wire \u2_Display/lt57_c16 ;
  wire \u2_Display/lt57_c17 ;
  wire \u2_Display/lt57_c18 ;
  wire \u2_Display/lt57_c19 ;
  wire \u2_Display/lt57_c2 ;
  wire \u2_Display/lt57_c20 ;
  wire \u2_Display/lt57_c21 ;
  wire \u2_Display/lt57_c22 ;
  wire \u2_Display/lt57_c23 ;
  wire \u2_Display/lt57_c24 ;
  wire \u2_Display/lt57_c25 ;
  wire \u2_Display/lt57_c26 ;
  wire \u2_Display/lt57_c27 ;
  wire \u2_Display/lt57_c28 ;
  wire \u2_Display/lt57_c29 ;
  wire \u2_Display/lt57_c3 ;
  wire \u2_Display/lt57_c30 ;
  wire \u2_Display/lt57_c31 ;
  wire \u2_Display/lt57_c32 ;
  wire \u2_Display/lt57_c4 ;
  wire \u2_Display/lt57_c5 ;
  wire \u2_Display/lt57_c6 ;
  wire \u2_Display/lt57_c7 ;
  wire \u2_Display/lt57_c8 ;
  wire \u2_Display/lt57_c9 ;
  wire \u2_Display/lt58_c0 ;
  wire \u2_Display/lt58_c1 ;
  wire \u2_Display/lt58_c10 ;
  wire \u2_Display/lt58_c11 ;
  wire \u2_Display/lt58_c12 ;
  wire \u2_Display/lt58_c13 ;
  wire \u2_Display/lt58_c14 ;
  wire \u2_Display/lt58_c15 ;
  wire \u2_Display/lt58_c16 ;
  wire \u2_Display/lt58_c17 ;
  wire \u2_Display/lt58_c18 ;
  wire \u2_Display/lt58_c19 ;
  wire \u2_Display/lt58_c2 ;
  wire \u2_Display/lt58_c20 ;
  wire \u2_Display/lt58_c21 ;
  wire \u2_Display/lt58_c22 ;
  wire \u2_Display/lt58_c23 ;
  wire \u2_Display/lt58_c24 ;
  wire \u2_Display/lt58_c25 ;
  wire \u2_Display/lt58_c26 ;
  wire \u2_Display/lt58_c27 ;
  wire \u2_Display/lt58_c28 ;
  wire \u2_Display/lt58_c29 ;
  wire \u2_Display/lt58_c3 ;
  wire \u2_Display/lt58_c30 ;
  wire \u2_Display/lt58_c31 ;
  wire \u2_Display/lt58_c32 ;
  wire \u2_Display/lt58_c4 ;
  wire \u2_Display/lt58_c5 ;
  wire \u2_Display/lt58_c6 ;
  wire \u2_Display/lt58_c7 ;
  wire \u2_Display/lt58_c8 ;
  wire \u2_Display/lt58_c9 ;
  wire \u2_Display/lt59_c0 ;
  wire \u2_Display/lt59_c1 ;
  wire \u2_Display/lt59_c10 ;
  wire \u2_Display/lt59_c11 ;
  wire \u2_Display/lt59_c12 ;
  wire \u2_Display/lt59_c13 ;
  wire \u2_Display/lt59_c14 ;
  wire \u2_Display/lt59_c15 ;
  wire \u2_Display/lt59_c16 ;
  wire \u2_Display/lt59_c17 ;
  wire \u2_Display/lt59_c18 ;
  wire \u2_Display/lt59_c19 ;
  wire \u2_Display/lt59_c2 ;
  wire \u2_Display/lt59_c20 ;
  wire \u2_Display/lt59_c21 ;
  wire \u2_Display/lt59_c22 ;
  wire \u2_Display/lt59_c23 ;
  wire \u2_Display/lt59_c24 ;
  wire \u2_Display/lt59_c25 ;
  wire \u2_Display/lt59_c26 ;
  wire \u2_Display/lt59_c27 ;
  wire \u2_Display/lt59_c28 ;
  wire \u2_Display/lt59_c29 ;
  wire \u2_Display/lt59_c3 ;
  wire \u2_Display/lt59_c30 ;
  wire \u2_Display/lt59_c31 ;
  wire \u2_Display/lt59_c32 ;
  wire \u2_Display/lt59_c4 ;
  wire \u2_Display/lt59_c5 ;
  wire \u2_Display/lt59_c6 ;
  wire \u2_Display/lt59_c7 ;
  wire \u2_Display/lt59_c8 ;
  wire \u2_Display/lt59_c9 ;
  wire \u2_Display/lt5_2_c0 ;
  wire \u2_Display/lt5_2_c1 ;
  wire \u2_Display/lt5_2_c10 ;
  wire \u2_Display/lt5_2_c11 ;
  wire \u2_Display/lt5_2_c12 ;
  wire \u2_Display/lt5_2_c13 ;
  wire \u2_Display/lt5_2_c2 ;
  wire \u2_Display/lt5_2_c3 ;
  wire \u2_Display/lt5_2_c4 ;
  wire \u2_Display/lt5_2_c5 ;
  wire \u2_Display/lt5_2_c6 ;
  wire \u2_Display/lt5_2_c7 ;
  wire \u2_Display/lt5_2_c8 ;
  wire \u2_Display/lt5_2_c9 ;
  wire \u2_Display/lt60_c0 ;
  wire \u2_Display/lt60_c1 ;
  wire \u2_Display/lt60_c10 ;
  wire \u2_Display/lt60_c11 ;
  wire \u2_Display/lt60_c12 ;
  wire \u2_Display/lt60_c13 ;
  wire \u2_Display/lt60_c14 ;
  wire \u2_Display/lt60_c15 ;
  wire \u2_Display/lt60_c16 ;
  wire \u2_Display/lt60_c17 ;
  wire \u2_Display/lt60_c18 ;
  wire \u2_Display/lt60_c19 ;
  wire \u2_Display/lt60_c2 ;
  wire \u2_Display/lt60_c20 ;
  wire \u2_Display/lt60_c21 ;
  wire \u2_Display/lt60_c22 ;
  wire \u2_Display/lt60_c23 ;
  wire \u2_Display/lt60_c24 ;
  wire \u2_Display/lt60_c25 ;
  wire \u2_Display/lt60_c26 ;
  wire \u2_Display/lt60_c27 ;
  wire \u2_Display/lt60_c28 ;
  wire \u2_Display/lt60_c29 ;
  wire \u2_Display/lt60_c3 ;
  wire \u2_Display/lt60_c30 ;
  wire \u2_Display/lt60_c31 ;
  wire \u2_Display/lt60_c32 ;
  wire \u2_Display/lt60_c4 ;
  wire \u2_Display/lt60_c5 ;
  wire \u2_Display/lt60_c6 ;
  wire \u2_Display/lt60_c7 ;
  wire \u2_Display/lt60_c8 ;
  wire \u2_Display/lt60_c9 ;
  wire \u2_Display/lt61_c0 ;
  wire \u2_Display/lt61_c1 ;
  wire \u2_Display/lt61_c10 ;
  wire \u2_Display/lt61_c11 ;
  wire \u2_Display/lt61_c12 ;
  wire \u2_Display/lt61_c13 ;
  wire \u2_Display/lt61_c14 ;
  wire \u2_Display/lt61_c15 ;
  wire \u2_Display/lt61_c16 ;
  wire \u2_Display/lt61_c17 ;
  wire \u2_Display/lt61_c18 ;
  wire \u2_Display/lt61_c19 ;
  wire \u2_Display/lt61_c2 ;
  wire \u2_Display/lt61_c20 ;
  wire \u2_Display/lt61_c21 ;
  wire \u2_Display/lt61_c22 ;
  wire \u2_Display/lt61_c23 ;
  wire \u2_Display/lt61_c24 ;
  wire \u2_Display/lt61_c25 ;
  wire \u2_Display/lt61_c26 ;
  wire \u2_Display/lt61_c27 ;
  wire \u2_Display/lt61_c28 ;
  wire \u2_Display/lt61_c29 ;
  wire \u2_Display/lt61_c3 ;
  wire \u2_Display/lt61_c30 ;
  wire \u2_Display/lt61_c31 ;
  wire \u2_Display/lt61_c32 ;
  wire \u2_Display/lt61_c4 ;
  wire \u2_Display/lt61_c5 ;
  wire \u2_Display/lt61_c6 ;
  wire \u2_Display/lt61_c7 ;
  wire \u2_Display/lt61_c8 ;
  wire \u2_Display/lt61_c9 ;
  wire \u2_Display/lt62_c0 ;
  wire \u2_Display/lt62_c1 ;
  wire \u2_Display/lt62_c10 ;
  wire \u2_Display/lt62_c11 ;
  wire \u2_Display/lt62_c12 ;
  wire \u2_Display/lt62_c13 ;
  wire \u2_Display/lt62_c14 ;
  wire \u2_Display/lt62_c15 ;
  wire \u2_Display/lt62_c16 ;
  wire \u2_Display/lt62_c17 ;
  wire \u2_Display/lt62_c18 ;
  wire \u2_Display/lt62_c19 ;
  wire \u2_Display/lt62_c2 ;
  wire \u2_Display/lt62_c20 ;
  wire \u2_Display/lt62_c21 ;
  wire \u2_Display/lt62_c22 ;
  wire \u2_Display/lt62_c23 ;
  wire \u2_Display/lt62_c24 ;
  wire \u2_Display/lt62_c25 ;
  wire \u2_Display/lt62_c26 ;
  wire \u2_Display/lt62_c27 ;
  wire \u2_Display/lt62_c28 ;
  wire \u2_Display/lt62_c29 ;
  wire \u2_Display/lt62_c3 ;
  wire \u2_Display/lt62_c30 ;
  wire \u2_Display/lt62_c31 ;
  wire \u2_Display/lt62_c32 ;
  wire \u2_Display/lt62_c4 ;
  wire \u2_Display/lt62_c5 ;
  wire \u2_Display/lt62_c6 ;
  wire \u2_Display/lt62_c7 ;
  wire \u2_Display/lt62_c8 ;
  wire \u2_Display/lt62_c9 ;
  wire \u2_Display/lt63_c0 ;
  wire \u2_Display/lt63_c1 ;
  wire \u2_Display/lt63_c10 ;
  wire \u2_Display/lt63_c11 ;
  wire \u2_Display/lt63_c12 ;
  wire \u2_Display/lt63_c13 ;
  wire \u2_Display/lt63_c14 ;
  wire \u2_Display/lt63_c15 ;
  wire \u2_Display/lt63_c16 ;
  wire \u2_Display/lt63_c17 ;
  wire \u2_Display/lt63_c18 ;
  wire \u2_Display/lt63_c19 ;
  wire \u2_Display/lt63_c2 ;
  wire \u2_Display/lt63_c20 ;
  wire \u2_Display/lt63_c21 ;
  wire \u2_Display/lt63_c22 ;
  wire \u2_Display/lt63_c23 ;
  wire \u2_Display/lt63_c24 ;
  wire \u2_Display/lt63_c25 ;
  wire \u2_Display/lt63_c26 ;
  wire \u2_Display/lt63_c27 ;
  wire \u2_Display/lt63_c28 ;
  wire \u2_Display/lt63_c29 ;
  wire \u2_Display/lt63_c3 ;
  wire \u2_Display/lt63_c30 ;
  wire \u2_Display/lt63_c31 ;
  wire \u2_Display/lt63_c32 ;
  wire \u2_Display/lt63_c4 ;
  wire \u2_Display/lt63_c5 ;
  wire \u2_Display/lt63_c6 ;
  wire \u2_Display/lt63_c7 ;
  wire \u2_Display/lt63_c8 ;
  wire \u2_Display/lt63_c9 ;
  wire \u2_Display/lt64_c0 ;
  wire \u2_Display/lt64_c1 ;
  wire \u2_Display/lt64_c10 ;
  wire \u2_Display/lt64_c11 ;
  wire \u2_Display/lt64_c12 ;
  wire \u2_Display/lt64_c13 ;
  wire \u2_Display/lt64_c14 ;
  wire \u2_Display/lt64_c15 ;
  wire \u2_Display/lt64_c16 ;
  wire \u2_Display/lt64_c17 ;
  wire \u2_Display/lt64_c18 ;
  wire \u2_Display/lt64_c19 ;
  wire \u2_Display/lt64_c2 ;
  wire \u2_Display/lt64_c20 ;
  wire \u2_Display/lt64_c21 ;
  wire \u2_Display/lt64_c22 ;
  wire \u2_Display/lt64_c23 ;
  wire \u2_Display/lt64_c24 ;
  wire \u2_Display/lt64_c25 ;
  wire \u2_Display/lt64_c26 ;
  wire \u2_Display/lt64_c27 ;
  wire \u2_Display/lt64_c28 ;
  wire \u2_Display/lt64_c29 ;
  wire \u2_Display/lt64_c3 ;
  wire \u2_Display/lt64_c30 ;
  wire \u2_Display/lt64_c31 ;
  wire \u2_Display/lt64_c32 ;
  wire \u2_Display/lt64_c4 ;
  wire \u2_Display/lt64_c5 ;
  wire \u2_Display/lt64_c6 ;
  wire \u2_Display/lt64_c7 ;
  wire \u2_Display/lt64_c8 ;
  wire \u2_Display/lt64_c9 ;
  wire \u2_Display/lt65_c0 ;
  wire \u2_Display/lt65_c1 ;
  wire \u2_Display/lt65_c10 ;
  wire \u2_Display/lt65_c11 ;
  wire \u2_Display/lt65_c12 ;
  wire \u2_Display/lt65_c13 ;
  wire \u2_Display/lt65_c14 ;
  wire \u2_Display/lt65_c15 ;
  wire \u2_Display/lt65_c16 ;
  wire \u2_Display/lt65_c17 ;
  wire \u2_Display/lt65_c18 ;
  wire \u2_Display/lt65_c19 ;
  wire \u2_Display/lt65_c2 ;
  wire \u2_Display/lt65_c20 ;
  wire \u2_Display/lt65_c21 ;
  wire \u2_Display/lt65_c22 ;
  wire \u2_Display/lt65_c23 ;
  wire \u2_Display/lt65_c24 ;
  wire \u2_Display/lt65_c25 ;
  wire \u2_Display/lt65_c26 ;
  wire \u2_Display/lt65_c27 ;
  wire \u2_Display/lt65_c28 ;
  wire \u2_Display/lt65_c29 ;
  wire \u2_Display/lt65_c3 ;
  wire \u2_Display/lt65_c30 ;
  wire \u2_Display/lt65_c31 ;
  wire \u2_Display/lt65_c32 ;
  wire \u2_Display/lt65_c4 ;
  wire \u2_Display/lt65_c5 ;
  wire \u2_Display/lt65_c6 ;
  wire \u2_Display/lt65_c7 ;
  wire \u2_Display/lt65_c8 ;
  wire \u2_Display/lt65_c9 ;
  wire \u2_Display/lt66_c0 ;
  wire \u2_Display/lt66_c1 ;
  wire \u2_Display/lt66_c10 ;
  wire \u2_Display/lt66_c11 ;
  wire \u2_Display/lt66_c12 ;
  wire \u2_Display/lt66_c13 ;
  wire \u2_Display/lt66_c14 ;
  wire \u2_Display/lt66_c15 ;
  wire \u2_Display/lt66_c16 ;
  wire \u2_Display/lt66_c17 ;
  wire \u2_Display/lt66_c18 ;
  wire \u2_Display/lt66_c19 ;
  wire \u2_Display/lt66_c2 ;
  wire \u2_Display/lt66_c20 ;
  wire \u2_Display/lt66_c21 ;
  wire \u2_Display/lt66_c22 ;
  wire \u2_Display/lt66_c23 ;
  wire \u2_Display/lt66_c24 ;
  wire \u2_Display/lt66_c25 ;
  wire \u2_Display/lt66_c26 ;
  wire \u2_Display/lt66_c27 ;
  wire \u2_Display/lt66_c28 ;
  wire \u2_Display/lt66_c29 ;
  wire \u2_Display/lt66_c3 ;
  wire \u2_Display/lt66_c30 ;
  wire \u2_Display/lt66_c31 ;
  wire \u2_Display/lt66_c32 ;
  wire \u2_Display/lt66_c4 ;
  wire \u2_Display/lt66_c5 ;
  wire \u2_Display/lt66_c6 ;
  wire \u2_Display/lt66_c7 ;
  wire \u2_Display/lt66_c8 ;
  wire \u2_Display/lt66_c9 ;
  wire \u2_Display/lt67_c0 ;
  wire \u2_Display/lt67_c1 ;
  wire \u2_Display/lt67_c10 ;
  wire \u2_Display/lt67_c11 ;
  wire \u2_Display/lt67_c12 ;
  wire \u2_Display/lt67_c13 ;
  wire \u2_Display/lt67_c14 ;
  wire \u2_Display/lt67_c15 ;
  wire \u2_Display/lt67_c16 ;
  wire \u2_Display/lt67_c17 ;
  wire \u2_Display/lt67_c18 ;
  wire \u2_Display/lt67_c19 ;
  wire \u2_Display/lt67_c2 ;
  wire \u2_Display/lt67_c20 ;
  wire \u2_Display/lt67_c21 ;
  wire \u2_Display/lt67_c22 ;
  wire \u2_Display/lt67_c23 ;
  wire \u2_Display/lt67_c24 ;
  wire \u2_Display/lt67_c25 ;
  wire \u2_Display/lt67_c26 ;
  wire \u2_Display/lt67_c27 ;
  wire \u2_Display/lt67_c28 ;
  wire \u2_Display/lt67_c29 ;
  wire \u2_Display/lt67_c3 ;
  wire \u2_Display/lt67_c30 ;
  wire \u2_Display/lt67_c31 ;
  wire \u2_Display/lt67_c32 ;
  wire \u2_Display/lt67_c4 ;
  wire \u2_Display/lt67_c5 ;
  wire \u2_Display/lt67_c6 ;
  wire \u2_Display/lt67_c7 ;
  wire \u2_Display/lt67_c8 ;
  wire \u2_Display/lt67_c9 ;
  wire \u2_Display/lt68_c0 ;
  wire \u2_Display/lt68_c1 ;
  wire \u2_Display/lt68_c10 ;
  wire \u2_Display/lt68_c11 ;
  wire \u2_Display/lt68_c12 ;
  wire \u2_Display/lt68_c13 ;
  wire \u2_Display/lt68_c14 ;
  wire \u2_Display/lt68_c15 ;
  wire \u2_Display/lt68_c16 ;
  wire \u2_Display/lt68_c17 ;
  wire \u2_Display/lt68_c18 ;
  wire \u2_Display/lt68_c19 ;
  wire \u2_Display/lt68_c2 ;
  wire \u2_Display/lt68_c20 ;
  wire \u2_Display/lt68_c21 ;
  wire \u2_Display/lt68_c22 ;
  wire \u2_Display/lt68_c23 ;
  wire \u2_Display/lt68_c24 ;
  wire \u2_Display/lt68_c25 ;
  wire \u2_Display/lt68_c26 ;
  wire \u2_Display/lt68_c27 ;
  wire \u2_Display/lt68_c28 ;
  wire \u2_Display/lt68_c29 ;
  wire \u2_Display/lt68_c3 ;
  wire \u2_Display/lt68_c30 ;
  wire \u2_Display/lt68_c31 ;
  wire \u2_Display/lt68_c32 ;
  wire \u2_Display/lt68_c4 ;
  wire \u2_Display/lt68_c5 ;
  wire \u2_Display/lt68_c6 ;
  wire \u2_Display/lt68_c7 ;
  wire \u2_Display/lt68_c8 ;
  wire \u2_Display/lt68_c9 ;
  wire \u2_Display/lt69_c0 ;
  wire \u2_Display/lt69_c1 ;
  wire \u2_Display/lt69_c10 ;
  wire \u2_Display/lt69_c11 ;
  wire \u2_Display/lt69_c12 ;
  wire \u2_Display/lt69_c13 ;
  wire \u2_Display/lt69_c14 ;
  wire \u2_Display/lt69_c15 ;
  wire \u2_Display/lt69_c16 ;
  wire \u2_Display/lt69_c17 ;
  wire \u2_Display/lt69_c18 ;
  wire \u2_Display/lt69_c19 ;
  wire \u2_Display/lt69_c2 ;
  wire \u2_Display/lt69_c20 ;
  wire \u2_Display/lt69_c21 ;
  wire \u2_Display/lt69_c22 ;
  wire \u2_Display/lt69_c23 ;
  wire \u2_Display/lt69_c24 ;
  wire \u2_Display/lt69_c25 ;
  wire \u2_Display/lt69_c26 ;
  wire \u2_Display/lt69_c27 ;
  wire \u2_Display/lt69_c28 ;
  wire \u2_Display/lt69_c29 ;
  wire \u2_Display/lt69_c3 ;
  wire \u2_Display/lt69_c30 ;
  wire \u2_Display/lt69_c31 ;
  wire \u2_Display/lt69_c32 ;
  wire \u2_Display/lt69_c4 ;
  wire \u2_Display/lt69_c5 ;
  wire \u2_Display/lt69_c6 ;
  wire \u2_Display/lt69_c7 ;
  wire \u2_Display/lt69_c8 ;
  wire \u2_Display/lt69_c9 ;
  wire \u2_Display/lt6_2_c0 ;
  wire \u2_Display/lt6_2_c1 ;
  wire \u2_Display/lt6_2_c10 ;
  wire \u2_Display/lt6_2_c11 ;
  wire \u2_Display/lt6_2_c12 ;
  wire \u2_Display/lt6_2_c2 ;
  wire \u2_Display/lt6_2_c3 ;
  wire \u2_Display/lt6_2_c4 ;
  wire \u2_Display/lt6_2_c5 ;
  wire \u2_Display/lt6_2_c6 ;
  wire \u2_Display/lt6_2_c7 ;
  wire \u2_Display/lt6_2_c8 ;
  wire \u2_Display/lt6_2_c9 ;
  wire \u2_Display/lt70_c0 ;
  wire \u2_Display/lt70_c1 ;
  wire \u2_Display/lt70_c10 ;
  wire \u2_Display/lt70_c11 ;
  wire \u2_Display/lt70_c12 ;
  wire \u2_Display/lt70_c13 ;
  wire \u2_Display/lt70_c14 ;
  wire \u2_Display/lt70_c15 ;
  wire \u2_Display/lt70_c16 ;
  wire \u2_Display/lt70_c17 ;
  wire \u2_Display/lt70_c18 ;
  wire \u2_Display/lt70_c19 ;
  wire \u2_Display/lt70_c2 ;
  wire \u2_Display/lt70_c20 ;
  wire \u2_Display/lt70_c21 ;
  wire \u2_Display/lt70_c22 ;
  wire \u2_Display/lt70_c23 ;
  wire \u2_Display/lt70_c24 ;
  wire \u2_Display/lt70_c25 ;
  wire \u2_Display/lt70_c26 ;
  wire \u2_Display/lt70_c27 ;
  wire \u2_Display/lt70_c28 ;
  wire \u2_Display/lt70_c29 ;
  wire \u2_Display/lt70_c3 ;
  wire \u2_Display/lt70_c30 ;
  wire \u2_Display/lt70_c31 ;
  wire \u2_Display/lt70_c32 ;
  wire \u2_Display/lt70_c4 ;
  wire \u2_Display/lt70_c5 ;
  wire \u2_Display/lt70_c6 ;
  wire \u2_Display/lt70_c7 ;
  wire \u2_Display/lt70_c8 ;
  wire \u2_Display/lt70_c9 ;
  wire \u2_Display/lt71_c0 ;
  wire \u2_Display/lt71_c1 ;
  wire \u2_Display/lt71_c10 ;
  wire \u2_Display/lt71_c11 ;
  wire \u2_Display/lt71_c12 ;
  wire \u2_Display/lt71_c13 ;
  wire \u2_Display/lt71_c14 ;
  wire \u2_Display/lt71_c15 ;
  wire \u2_Display/lt71_c16 ;
  wire \u2_Display/lt71_c17 ;
  wire \u2_Display/lt71_c18 ;
  wire \u2_Display/lt71_c19 ;
  wire \u2_Display/lt71_c2 ;
  wire \u2_Display/lt71_c20 ;
  wire \u2_Display/lt71_c21 ;
  wire \u2_Display/lt71_c22 ;
  wire \u2_Display/lt71_c23 ;
  wire \u2_Display/lt71_c24 ;
  wire \u2_Display/lt71_c25 ;
  wire \u2_Display/lt71_c26 ;
  wire \u2_Display/lt71_c27 ;
  wire \u2_Display/lt71_c28 ;
  wire \u2_Display/lt71_c29 ;
  wire \u2_Display/lt71_c3 ;
  wire \u2_Display/lt71_c30 ;
  wire \u2_Display/lt71_c31 ;
  wire \u2_Display/lt71_c32 ;
  wire \u2_Display/lt71_c4 ;
  wire \u2_Display/lt71_c5 ;
  wire \u2_Display/lt71_c6 ;
  wire \u2_Display/lt71_c7 ;
  wire \u2_Display/lt71_c8 ;
  wire \u2_Display/lt71_c9 ;
  wire \u2_Display/lt72_c0 ;
  wire \u2_Display/lt72_c1 ;
  wire \u2_Display/lt72_c10 ;
  wire \u2_Display/lt72_c11 ;
  wire \u2_Display/lt72_c12 ;
  wire \u2_Display/lt72_c13 ;
  wire \u2_Display/lt72_c14 ;
  wire \u2_Display/lt72_c15 ;
  wire \u2_Display/lt72_c16 ;
  wire \u2_Display/lt72_c17 ;
  wire \u2_Display/lt72_c18 ;
  wire \u2_Display/lt72_c19 ;
  wire \u2_Display/lt72_c2 ;
  wire \u2_Display/lt72_c20 ;
  wire \u2_Display/lt72_c21 ;
  wire \u2_Display/lt72_c22 ;
  wire \u2_Display/lt72_c23 ;
  wire \u2_Display/lt72_c24 ;
  wire \u2_Display/lt72_c25 ;
  wire \u2_Display/lt72_c26 ;
  wire \u2_Display/lt72_c27 ;
  wire \u2_Display/lt72_c28 ;
  wire \u2_Display/lt72_c29 ;
  wire \u2_Display/lt72_c3 ;
  wire \u2_Display/lt72_c30 ;
  wire \u2_Display/lt72_c31 ;
  wire \u2_Display/lt72_c32 ;
  wire \u2_Display/lt72_c4 ;
  wire \u2_Display/lt72_c5 ;
  wire \u2_Display/lt72_c6 ;
  wire \u2_Display/lt72_c7 ;
  wire \u2_Display/lt72_c8 ;
  wire \u2_Display/lt72_c9 ;
  wire \u2_Display/lt73_c0 ;
  wire \u2_Display/lt73_c1 ;
  wire \u2_Display/lt73_c10 ;
  wire \u2_Display/lt73_c11 ;
  wire \u2_Display/lt73_c12 ;
  wire \u2_Display/lt73_c13 ;
  wire \u2_Display/lt73_c14 ;
  wire \u2_Display/lt73_c15 ;
  wire \u2_Display/lt73_c16 ;
  wire \u2_Display/lt73_c17 ;
  wire \u2_Display/lt73_c18 ;
  wire \u2_Display/lt73_c19 ;
  wire \u2_Display/lt73_c2 ;
  wire \u2_Display/lt73_c20 ;
  wire \u2_Display/lt73_c21 ;
  wire \u2_Display/lt73_c22 ;
  wire \u2_Display/lt73_c23 ;
  wire \u2_Display/lt73_c24 ;
  wire \u2_Display/lt73_c25 ;
  wire \u2_Display/lt73_c26 ;
  wire \u2_Display/lt73_c27 ;
  wire \u2_Display/lt73_c28 ;
  wire \u2_Display/lt73_c29 ;
  wire \u2_Display/lt73_c3 ;
  wire \u2_Display/lt73_c30 ;
  wire \u2_Display/lt73_c31 ;
  wire \u2_Display/lt73_c32 ;
  wire \u2_Display/lt73_c4 ;
  wire \u2_Display/lt73_c5 ;
  wire \u2_Display/lt73_c6 ;
  wire \u2_Display/lt73_c7 ;
  wire \u2_Display/lt73_c8 ;
  wire \u2_Display/lt73_c9 ;
  wire \u2_Display/lt74_c0 ;
  wire \u2_Display/lt74_c1 ;
  wire \u2_Display/lt74_c10 ;
  wire \u2_Display/lt74_c11 ;
  wire \u2_Display/lt74_c12 ;
  wire \u2_Display/lt74_c13 ;
  wire \u2_Display/lt74_c14 ;
  wire \u2_Display/lt74_c15 ;
  wire \u2_Display/lt74_c16 ;
  wire \u2_Display/lt74_c17 ;
  wire \u2_Display/lt74_c18 ;
  wire \u2_Display/lt74_c19 ;
  wire \u2_Display/lt74_c2 ;
  wire \u2_Display/lt74_c20 ;
  wire \u2_Display/lt74_c21 ;
  wire \u2_Display/lt74_c22 ;
  wire \u2_Display/lt74_c23 ;
  wire \u2_Display/lt74_c24 ;
  wire \u2_Display/lt74_c25 ;
  wire \u2_Display/lt74_c26 ;
  wire \u2_Display/lt74_c27 ;
  wire \u2_Display/lt74_c28 ;
  wire \u2_Display/lt74_c29 ;
  wire \u2_Display/lt74_c3 ;
  wire \u2_Display/lt74_c30 ;
  wire \u2_Display/lt74_c31 ;
  wire \u2_Display/lt74_c32 ;
  wire \u2_Display/lt74_c4 ;
  wire \u2_Display/lt74_c5 ;
  wire \u2_Display/lt74_c6 ;
  wire \u2_Display/lt74_c7 ;
  wire \u2_Display/lt74_c8 ;
  wire \u2_Display/lt74_c9 ;
  wire \u2_Display/lt75_c0 ;
  wire \u2_Display/lt75_c1 ;
  wire \u2_Display/lt75_c10 ;
  wire \u2_Display/lt75_c11 ;
  wire \u2_Display/lt75_c12 ;
  wire \u2_Display/lt75_c13 ;
  wire \u2_Display/lt75_c14 ;
  wire \u2_Display/lt75_c15 ;
  wire \u2_Display/lt75_c16 ;
  wire \u2_Display/lt75_c17 ;
  wire \u2_Display/lt75_c18 ;
  wire \u2_Display/lt75_c19 ;
  wire \u2_Display/lt75_c2 ;
  wire \u2_Display/lt75_c20 ;
  wire \u2_Display/lt75_c21 ;
  wire \u2_Display/lt75_c22 ;
  wire \u2_Display/lt75_c23 ;
  wire \u2_Display/lt75_c24 ;
  wire \u2_Display/lt75_c25 ;
  wire \u2_Display/lt75_c26 ;
  wire \u2_Display/lt75_c27 ;
  wire \u2_Display/lt75_c28 ;
  wire \u2_Display/lt75_c29 ;
  wire \u2_Display/lt75_c3 ;
  wire \u2_Display/lt75_c30 ;
  wire \u2_Display/lt75_c31 ;
  wire \u2_Display/lt75_c32 ;
  wire \u2_Display/lt75_c4 ;
  wire \u2_Display/lt75_c5 ;
  wire \u2_Display/lt75_c6 ;
  wire \u2_Display/lt75_c7 ;
  wire \u2_Display/lt75_c8 ;
  wire \u2_Display/lt75_c9 ;
  wire \u2_Display/lt76_c0 ;
  wire \u2_Display/lt76_c1 ;
  wire \u2_Display/lt76_c10 ;
  wire \u2_Display/lt76_c11 ;
  wire \u2_Display/lt76_c12 ;
  wire \u2_Display/lt76_c13 ;
  wire \u2_Display/lt76_c14 ;
  wire \u2_Display/lt76_c15 ;
  wire \u2_Display/lt76_c16 ;
  wire \u2_Display/lt76_c17 ;
  wire \u2_Display/lt76_c18 ;
  wire \u2_Display/lt76_c19 ;
  wire \u2_Display/lt76_c2 ;
  wire \u2_Display/lt76_c20 ;
  wire \u2_Display/lt76_c21 ;
  wire \u2_Display/lt76_c22 ;
  wire \u2_Display/lt76_c23 ;
  wire \u2_Display/lt76_c24 ;
  wire \u2_Display/lt76_c25 ;
  wire \u2_Display/lt76_c26 ;
  wire \u2_Display/lt76_c27 ;
  wire \u2_Display/lt76_c28 ;
  wire \u2_Display/lt76_c29 ;
  wire \u2_Display/lt76_c3 ;
  wire \u2_Display/lt76_c30 ;
  wire \u2_Display/lt76_c31 ;
  wire \u2_Display/lt76_c32 ;
  wire \u2_Display/lt76_c4 ;
  wire \u2_Display/lt76_c5 ;
  wire \u2_Display/lt76_c6 ;
  wire \u2_Display/lt76_c7 ;
  wire \u2_Display/lt76_c8 ;
  wire \u2_Display/lt76_c9 ;
  wire \u2_Display/lt77_c0 ;
  wire \u2_Display/lt77_c1 ;
  wire \u2_Display/lt77_c10 ;
  wire \u2_Display/lt77_c11 ;
  wire \u2_Display/lt77_c12 ;
  wire \u2_Display/lt77_c13 ;
  wire \u2_Display/lt77_c14 ;
  wire \u2_Display/lt77_c15 ;
  wire \u2_Display/lt77_c16 ;
  wire \u2_Display/lt77_c17 ;
  wire \u2_Display/lt77_c18 ;
  wire \u2_Display/lt77_c19 ;
  wire \u2_Display/lt77_c2 ;
  wire \u2_Display/lt77_c20 ;
  wire \u2_Display/lt77_c21 ;
  wire \u2_Display/lt77_c22 ;
  wire \u2_Display/lt77_c23 ;
  wire \u2_Display/lt77_c24 ;
  wire \u2_Display/lt77_c25 ;
  wire \u2_Display/lt77_c26 ;
  wire \u2_Display/lt77_c27 ;
  wire \u2_Display/lt77_c28 ;
  wire \u2_Display/lt77_c29 ;
  wire \u2_Display/lt77_c3 ;
  wire \u2_Display/lt77_c30 ;
  wire \u2_Display/lt77_c31 ;
  wire \u2_Display/lt77_c32 ;
  wire \u2_Display/lt77_c4 ;
  wire \u2_Display/lt77_c5 ;
  wire \u2_Display/lt77_c6 ;
  wire \u2_Display/lt77_c7 ;
  wire \u2_Display/lt77_c8 ;
  wire \u2_Display/lt77_c9 ;
  wire \u2_Display/lt7_2_c0 ;
  wire \u2_Display/lt7_2_c1 ;
  wire \u2_Display/lt7_2_c10 ;
  wire \u2_Display/lt7_2_c11 ;
  wire \u2_Display/lt7_2_c12 ;
  wire \u2_Display/lt7_2_c13 ;
  wire \u2_Display/lt7_2_c2 ;
  wire \u2_Display/lt7_2_c3 ;
  wire \u2_Display/lt7_2_c4 ;
  wire \u2_Display/lt7_2_c5 ;
  wire \u2_Display/lt7_2_c6 ;
  wire \u2_Display/lt7_2_c7 ;
  wire \u2_Display/lt7_2_c8 ;
  wire \u2_Display/lt7_2_c9 ;
  wire \u2_Display/lt88_c0 ;
  wire \u2_Display/lt88_c1 ;
  wire \u2_Display/lt88_c10 ;
  wire \u2_Display/lt88_c11 ;
  wire \u2_Display/lt88_c12 ;
  wire \u2_Display/lt88_c13 ;
  wire \u2_Display/lt88_c14 ;
  wire \u2_Display/lt88_c15 ;
  wire \u2_Display/lt88_c16 ;
  wire \u2_Display/lt88_c17 ;
  wire \u2_Display/lt88_c18 ;
  wire \u2_Display/lt88_c19 ;
  wire \u2_Display/lt88_c2 ;
  wire \u2_Display/lt88_c20 ;
  wire \u2_Display/lt88_c21 ;
  wire \u2_Display/lt88_c22 ;
  wire \u2_Display/lt88_c23 ;
  wire \u2_Display/lt88_c24 ;
  wire \u2_Display/lt88_c25 ;
  wire \u2_Display/lt88_c26 ;
  wire \u2_Display/lt88_c27 ;
  wire \u2_Display/lt88_c28 ;
  wire \u2_Display/lt88_c29 ;
  wire \u2_Display/lt88_c3 ;
  wire \u2_Display/lt88_c30 ;
  wire \u2_Display/lt88_c31 ;
  wire \u2_Display/lt88_c32 ;
  wire \u2_Display/lt88_c4 ;
  wire \u2_Display/lt88_c5 ;
  wire \u2_Display/lt88_c6 ;
  wire \u2_Display/lt88_c7 ;
  wire \u2_Display/lt88_c8 ;
  wire \u2_Display/lt88_c9 ;
  wire \u2_Display/lt89_c0 ;
  wire \u2_Display/lt89_c1 ;
  wire \u2_Display/lt89_c10 ;
  wire \u2_Display/lt89_c11 ;
  wire \u2_Display/lt89_c12 ;
  wire \u2_Display/lt89_c13 ;
  wire \u2_Display/lt89_c14 ;
  wire \u2_Display/lt89_c15 ;
  wire \u2_Display/lt89_c16 ;
  wire \u2_Display/lt89_c17 ;
  wire \u2_Display/lt89_c18 ;
  wire \u2_Display/lt89_c19 ;
  wire \u2_Display/lt89_c2 ;
  wire \u2_Display/lt89_c20 ;
  wire \u2_Display/lt89_c21 ;
  wire \u2_Display/lt89_c22 ;
  wire \u2_Display/lt89_c23 ;
  wire \u2_Display/lt89_c24 ;
  wire \u2_Display/lt89_c25 ;
  wire \u2_Display/lt89_c26 ;
  wire \u2_Display/lt89_c27 ;
  wire \u2_Display/lt89_c28 ;
  wire \u2_Display/lt89_c29 ;
  wire \u2_Display/lt89_c3 ;
  wire \u2_Display/lt89_c30 ;
  wire \u2_Display/lt89_c31 ;
  wire \u2_Display/lt89_c32 ;
  wire \u2_Display/lt89_c4 ;
  wire \u2_Display/lt89_c5 ;
  wire \u2_Display/lt89_c6 ;
  wire \u2_Display/lt89_c7 ;
  wire \u2_Display/lt89_c8 ;
  wire \u2_Display/lt89_c9 ;
  wire \u2_Display/lt8_2_c0 ;
  wire \u2_Display/lt8_2_c1 ;
  wire \u2_Display/lt8_2_c10 ;
  wire \u2_Display/lt8_2_c11 ;
  wire \u2_Display/lt8_2_c12 ;
  wire \u2_Display/lt8_2_c2 ;
  wire \u2_Display/lt8_2_c3 ;
  wire \u2_Display/lt8_2_c4 ;
  wire \u2_Display/lt8_2_c5 ;
  wire \u2_Display/lt8_2_c6 ;
  wire \u2_Display/lt8_2_c7 ;
  wire \u2_Display/lt8_2_c8 ;
  wire \u2_Display/lt8_2_c9 ;
  wire \u2_Display/lt90_c0 ;
  wire \u2_Display/lt90_c1 ;
  wire \u2_Display/lt90_c10 ;
  wire \u2_Display/lt90_c11 ;
  wire \u2_Display/lt90_c12 ;
  wire \u2_Display/lt90_c13 ;
  wire \u2_Display/lt90_c14 ;
  wire \u2_Display/lt90_c15 ;
  wire \u2_Display/lt90_c16 ;
  wire \u2_Display/lt90_c17 ;
  wire \u2_Display/lt90_c18 ;
  wire \u2_Display/lt90_c19 ;
  wire \u2_Display/lt90_c2 ;
  wire \u2_Display/lt90_c20 ;
  wire \u2_Display/lt90_c21 ;
  wire \u2_Display/lt90_c22 ;
  wire \u2_Display/lt90_c23 ;
  wire \u2_Display/lt90_c24 ;
  wire \u2_Display/lt90_c25 ;
  wire \u2_Display/lt90_c26 ;
  wire \u2_Display/lt90_c27 ;
  wire \u2_Display/lt90_c28 ;
  wire \u2_Display/lt90_c29 ;
  wire \u2_Display/lt90_c3 ;
  wire \u2_Display/lt90_c30 ;
  wire \u2_Display/lt90_c31 ;
  wire \u2_Display/lt90_c32 ;
  wire \u2_Display/lt90_c4 ;
  wire \u2_Display/lt90_c5 ;
  wire \u2_Display/lt90_c6 ;
  wire \u2_Display/lt90_c7 ;
  wire \u2_Display/lt90_c8 ;
  wire \u2_Display/lt90_c9 ;
  wire \u2_Display/lt91_c0 ;
  wire \u2_Display/lt91_c1 ;
  wire \u2_Display/lt91_c10 ;
  wire \u2_Display/lt91_c11 ;
  wire \u2_Display/lt91_c12 ;
  wire \u2_Display/lt91_c13 ;
  wire \u2_Display/lt91_c14 ;
  wire \u2_Display/lt91_c15 ;
  wire \u2_Display/lt91_c16 ;
  wire \u2_Display/lt91_c17 ;
  wire \u2_Display/lt91_c18 ;
  wire \u2_Display/lt91_c19 ;
  wire \u2_Display/lt91_c2 ;
  wire \u2_Display/lt91_c20 ;
  wire \u2_Display/lt91_c21 ;
  wire \u2_Display/lt91_c22 ;
  wire \u2_Display/lt91_c23 ;
  wire \u2_Display/lt91_c24 ;
  wire \u2_Display/lt91_c25 ;
  wire \u2_Display/lt91_c26 ;
  wire \u2_Display/lt91_c27 ;
  wire \u2_Display/lt91_c28 ;
  wire \u2_Display/lt91_c29 ;
  wire \u2_Display/lt91_c3 ;
  wire \u2_Display/lt91_c30 ;
  wire \u2_Display/lt91_c31 ;
  wire \u2_Display/lt91_c32 ;
  wire \u2_Display/lt91_c4 ;
  wire \u2_Display/lt91_c5 ;
  wire \u2_Display/lt91_c6 ;
  wire \u2_Display/lt91_c7 ;
  wire \u2_Display/lt91_c8 ;
  wire \u2_Display/lt91_c9 ;
  wire \u2_Display/lt92_c0 ;
  wire \u2_Display/lt92_c1 ;
  wire \u2_Display/lt92_c10 ;
  wire \u2_Display/lt92_c11 ;
  wire \u2_Display/lt92_c12 ;
  wire \u2_Display/lt92_c13 ;
  wire \u2_Display/lt92_c14 ;
  wire \u2_Display/lt92_c15 ;
  wire \u2_Display/lt92_c16 ;
  wire \u2_Display/lt92_c17 ;
  wire \u2_Display/lt92_c18 ;
  wire \u2_Display/lt92_c19 ;
  wire \u2_Display/lt92_c2 ;
  wire \u2_Display/lt92_c20 ;
  wire \u2_Display/lt92_c21 ;
  wire \u2_Display/lt92_c22 ;
  wire \u2_Display/lt92_c23 ;
  wire \u2_Display/lt92_c24 ;
  wire \u2_Display/lt92_c25 ;
  wire \u2_Display/lt92_c26 ;
  wire \u2_Display/lt92_c27 ;
  wire \u2_Display/lt92_c28 ;
  wire \u2_Display/lt92_c29 ;
  wire \u2_Display/lt92_c3 ;
  wire \u2_Display/lt92_c30 ;
  wire \u2_Display/lt92_c31 ;
  wire \u2_Display/lt92_c32 ;
  wire \u2_Display/lt92_c4 ;
  wire \u2_Display/lt92_c5 ;
  wire \u2_Display/lt92_c6 ;
  wire \u2_Display/lt92_c7 ;
  wire \u2_Display/lt92_c8 ;
  wire \u2_Display/lt92_c9 ;
  wire \u2_Display/lt93_c0 ;
  wire \u2_Display/lt93_c1 ;
  wire \u2_Display/lt93_c10 ;
  wire \u2_Display/lt93_c11 ;
  wire \u2_Display/lt93_c12 ;
  wire \u2_Display/lt93_c13 ;
  wire \u2_Display/lt93_c14 ;
  wire \u2_Display/lt93_c15 ;
  wire \u2_Display/lt93_c16 ;
  wire \u2_Display/lt93_c17 ;
  wire \u2_Display/lt93_c18 ;
  wire \u2_Display/lt93_c19 ;
  wire \u2_Display/lt93_c2 ;
  wire \u2_Display/lt93_c20 ;
  wire \u2_Display/lt93_c21 ;
  wire \u2_Display/lt93_c22 ;
  wire \u2_Display/lt93_c23 ;
  wire \u2_Display/lt93_c24 ;
  wire \u2_Display/lt93_c25 ;
  wire \u2_Display/lt93_c26 ;
  wire \u2_Display/lt93_c27 ;
  wire \u2_Display/lt93_c28 ;
  wire \u2_Display/lt93_c29 ;
  wire \u2_Display/lt93_c3 ;
  wire \u2_Display/lt93_c30 ;
  wire \u2_Display/lt93_c31 ;
  wire \u2_Display/lt93_c32 ;
  wire \u2_Display/lt93_c4 ;
  wire \u2_Display/lt93_c5 ;
  wire \u2_Display/lt93_c6 ;
  wire \u2_Display/lt93_c7 ;
  wire \u2_Display/lt93_c8 ;
  wire \u2_Display/lt93_c9 ;
  wire \u2_Display/lt94_c0 ;
  wire \u2_Display/lt94_c1 ;
  wire \u2_Display/lt94_c10 ;
  wire \u2_Display/lt94_c11 ;
  wire \u2_Display/lt94_c12 ;
  wire \u2_Display/lt94_c13 ;
  wire \u2_Display/lt94_c14 ;
  wire \u2_Display/lt94_c15 ;
  wire \u2_Display/lt94_c16 ;
  wire \u2_Display/lt94_c17 ;
  wire \u2_Display/lt94_c18 ;
  wire \u2_Display/lt94_c19 ;
  wire \u2_Display/lt94_c2 ;
  wire \u2_Display/lt94_c20 ;
  wire \u2_Display/lt94_c21 ;
  wire \u2_Display/lt94_c22 ;
  wire \u2_Display/lt94_c23 ;
  wire \u2_Display/lt94_c24 ;
  wire \u2_Display/lt94_c25 ;
  wire \u2_Display/lt94_c26 ;
  wire \u2_Display/lt94_c27 ;
  wire \u2_Display/lt94_c28 ;
  wire \u2_Display/lt94_c29 ;
  wire \u2_Display/lt94_c3 ;
  wire \u2_Display/lt94_c30 ;
  wire \u2_Display/lt94_c31 ;
  wire \u2_Display/lt94_c32 ;
  wire \u2_Display/lt94_c4 ;
  wire \u2_Display/lt94_c5 ;
  wire \u2_Display/lt94_c6 ;
  wire \u2_Display/lt94_c7 ;
  wire \u2_Display/lt94_c8 ;
  wire \u2_Display/lt94_c9 ;
  wire \u2_Display/lt95_c0 ;
  wire \u2_Display/lt95_c1 ;
  wire \u2_Display/lt95_c10 ;
  wire \u2_Display/lt95_c11 ;
  wire \u2_Display/lt95_c12 ;
  wire \u2_Display/lt95_c13 ;
  wire \u2_Display/lt95_c14 ;
  wire \u2_Display/lt95_c15 ;
  wire \u2_Display/lt95_c16 ;
  wire \u2_Display/lt95_c17 ;
  wire \u2_Display/lt95_c18 ;
  wire \u2_Display/lt95_c19 ;
  wire \u2_Display/lt95_c2 ;
  wire \u2_Display/lt95_c20 ;
  wire \u2_Display/lt95_c21 ;
  wire \u2_Display/lt95_c22 ;
  wire \u2_Display/lt95_c23 ;
  wire \u2_Display/lt95_c24 ;
  wire \u2_Display/lt95_c25 ;
  wire \u2_Display/lt95_c26 ;
  wire \u2_Display/lt95_c27 ;
  wire \u2_Display/lt95_c28 ;
  wire \u2_Display/lt95_c29 ;
  wire \u2_Display/lt95_c3 ;
  wire \u2_Display/lt95_c30 ;
  wire \u2_Display/lt95_c31 ;
  wire \u2_Display/lt95_c32 ;
  wire \u2_Display/lt95_c4 ;
  wire \u2_Display/lt95_c5 ;
  wire \u2_Display/lt95_c6 ;
  wire \u2_Display/lt95_c7 ;
  wire \u2_Display/lt95_c8 ;
  wire \u2_Display/lt95_c9 ;
  wire \u2_Display/lt96_c0 ;
  wire \u2_Display/lt96_c1 ;
  wire \u2_Display/lt96_c10 ;
  wire \u2_Display/lt96_c11 ;
  wire \u2_Display/lt96_c12 ;
  wire \u2_Display/lt96_c13 ;
  wire \u2_Display/lt96_c14 ;
  wire \u2_Display/lt96_c15 ;
  wire \u2_Display/lt96_c16 ;
  wire \u2_Display/lt96_c17 ;
  wire \u2_Display/lt96_c18 ;
  wire \u2_Display/lt96_c19 ;
  wire \u2_Display/lt96_c2 ;
  wire \u2_Display/lt96_c20 ;
  wire \u2_Display/lt96_c21 ;
  wire \u2_Display/lt96_c22 ;
  wire \u2_Display/lt96_c23 ;
  wire \u2_Display/lt96_c24 ;
  wire \u2_Display/lt96_c25 ;
  wire \u2_Display/lt96_c26 ;
  wire \u2_Display/lt96_c27 ;
  wire \u2_Display/lt96_c28 ;
  wire \u2_Display/lt96_c29 ;
  wire \u2_Display/lt96_c3 ;
  wire \u2_Display/lt96_c30 ;
  wire \u2_Display/lt96_c31 ;
  wire \u2_Display/lt96_c32 ;
  wire \u2_Display/lt96_c4 ;
  wire \u2_Display/lt96_c5 ;
  wire \u2_Display/lt96_c6 ;
  wire \u2_Display/lt96_c7 ;
  wire \u2_Display/lt96_c8 ;
  wire \u2_Display/lt96_c9 ;
  wire \u2_Display/lt97_c0 ;
  wire \u2_Display/lt97_c1 ;
  wire \u2_Display/lt97_c10 ;
  wire \u2_Display/lt97_c11 ;
  wire \u2_Display/lt97_c12 ;
  wire \u2_Display/lt97_c13 ;
  wire \u2_Display/lt97_c14 ;
  wire \u2_Display/lt97_c15 ;
  wire \u2_Display/lt97_c16 ;
  wire \u2_Display/lt97_c17 ;
  wire \u2_Display/lt97_c18 ;
  wire \u2_Display/lt97_c19 ;
  wire \u2_Display/lt97_c2 ;
  wire \u2_Display/lt97_c20 ;
  wire \u2_Display/lt97_c21 ;
  wire \u2_Display/lt97_c22 ;
  wire \u2_Display/lt97_c23 ;
  wire \u2_Display/lt97_c24 ;
  wire \u2_Display/lt97_c25 ;
  wire \u2_Display/lt97_c26 ;
  wire \u2_Display/lt97_c27 ;
  wire \u2_Display/lt97_c28 ;
  wire \u2_Display/lt97_c29 ;
  wire \u2_Display/lt97_c3 ;
  wire \u2_Display/lt97_c30 ;
  wire \u2_Display/lt97_c31 ;
  wire \u2_Display/lt97_c32 ;
  wire \u2_Display/lt97_c4 ;
  wire \u2_Display/lt97_c5 ;
  wire \u2_Display/lt97_c6 ;
  wire \u2_Display/lt97_c7 ;
  wire \u2_Display/lt97_c8 ;
  wire \u2_Display/lt97_c9 ;
  wire \u2_Display/lt98_c0 ;
  wire \u2_Display/lt98_c1 ;
  wire \u2_Display/lt98_c10 ;
  wire \u2_Display/lt98_c11 ;
  wire \u2_Display/lt98_c12 ;
  wire \u2_Display/lt98_c13 ;
  wire \u2_Display/lt98_c14 ;
  wire \u2_Display/lt98_c15 ;
  wire \u2_Display/lt98_c16 ;
  wire \u2_Display/lt98_c17 ;
  wire \u2_Display/lt98_c18 ;
  wire \u2_Display/lt98_c19 ;
  wire \u2_Display/lt98_c2 ;
  wire \u2_Display/lt98_c20 ;
  wire \u2_Display/lt98_c21 ;
  wire \u2_Display/lt98_c22 ;
  wire \u2_Display/lt98_c23 ;
  wire \u2_Display/lt98_c24 ;
  wire \u2_Display/lt98_c25 ;
  wire \u2_Display/lt98_c26 ;
  wire \u2_Display/lt98_c27 ;
  wire \u2_Display/lt98_c28 ;
  wire \u2_Display/lt98_c29 ;
  wire \u2_Display/lt98_c3 ;
  wire \u2_Display/lt98_c30 ;
  wire \u2_Display/lt98_c31 ;
  wire \u2_Display/lt98_c32 ;
  wire \u2_Display/lt98_c4 ;
  wire \u2_Display/lt98_c5 ;
  wire \u2_Display/lt98_c6 ;
  wire \u2_Display/lt98_c7 ;
  wire \u2_Display/lt98_c8 ;
  wire \u2_Display/lt98_c9 ;
  wire \u2_Display/lt99_c0 ;
  wire \u2_Display/lt99_c1 ;
  wire \u2_Display/lt99_c10 ;
  wire \u2_Display/lt99_c11 ;
  wire \u2_Display/lt99_c12 ;
  wire \u2_Display/lt99_c13 ;
  wire \u2_Display/lt99_c14 ;
  wire \u2_Display/lt99_c15 ;
  wire \u2_Display/lt99_c16 ;
  wire \u2_Display/lt99_c17 ;
  wire \u2_Display/lt99_c18 ;
  wire \u2_Display/lt99_c19 ;
  wire \u2_Display/lt99_c2 ;
  wire \u2_Display/lt99_c20 ;
  wire \u2_Display/lt99_c21 ;
  wire \u2_Display/lt99_c22 ;
  wire \u2_Display/lt99_c23 ;
  wire \u2_Display/lt99_c24 ;
  wire \u2_Display/lt99_c25 ;
  wire \u2_Display/lt99_c26 ;
  wire \u2_Display/lt99_c27 ;
  wire \u2_Display/lt99_c28 ;
  wire \u2_Display/lt99_c29 ;
  wire \u2_Display/lt99_c3 ;
  wire \u2_Display/lt99_c30 ;
  wire \u2_Display/lt99_c31 ;
  wire \u2_Display/lt99_c32 ;
  wire \u2_Display/lt99_c4 ;
  wire \u2_Display/lt99_c5 ;
  wire \u2_Display/lt99_c6 ;
  wire \u2_Display/lt99_c7 ;
  wire \u2_Display/lt99_c8 ;
  wire \u2_Display/lt99_c9 ;
  wire \u2_Display/lt9_2_c0 ;
  wire \u2_Display/lt9_2_c1 ;
  wire \u2_Display/lt9_2_c10 ;
  wire \u2_Display/lt9_2_c11 ;
  wire \u2_Display/lt9_2_c12 ;
  wire \u2_Display/lt9_2_c13 ;
  wire \u2_Display/lt9_2_c2 ;
  wire \u2_Display/lt9_2_c3 ;
  wire \u2_Display/lt9_2_c4 ;
  wire \u2_Display/lt9_2_c5 ;
  wire \u2_Display/lt9_2_c6 ;
  wire \u2_Display/lt9_2_c7 ;
  wire \u2_Display/lt9_2_c8 ;
  wire \u2_Display/lt9_2_c9 ;
  wire \u2_Display/mux11_b0_sel_is_0_o ;
  wire \u2_Display/mux19_b0_sel_is_0_o ;
  wire \u2_Display/mux21_b0_sel_is_0_o ;
  wire \u2_Display/mux5_b0_sel_is_0_o ;
  wire \u2_Display/n100 ;
  wire \u2_Display/n1000 ;
  wire \u2_Display/n1001 ;
  wire \u2_Display/n1002 ;
  wire \u2_Display/n1003 ;
  wire \u2_Display/n1004 ;
  wire \u2_Display/n1005 ;
  wire \u2_Display/n1006 ;
  wire \u2_Display/n1007 ;
  wire \u2_Display/n1008 ;
  wire \u2_Display/n1009 ;
  wire \u2_Display/n1010 ;
  wire \u2_Display/n1011 ;
  wire \u2_Display/n1012 ;
  wire \u2_Display/n1015 ;
  wire \u2_Display/n1016 ;
  wire \u2_Display/n1017 ;
  wire \u2_Display/n1018 ;
  wire \u2_Display/n1019 ;
  wire \u2_Display/n1020 ;
  wire \u2_Display/n1021 ;
  wire \u2_Display/n1022 ;
  wire \u2_Display/n1023 ;
  wire \u2_Display/n1024 ;
  wire \u2_Display/n1025 ;
  wire \u2_Display/n1026 ;
  wire \u2_Display/n1027 ;
  wire \u2_Display/n1028 ;
  wire \u2_Display/n1029 ;
  wire \u2_Display/n103 ;
  wire \u2_Display/n1030 ;
  wire \u2_Display/n1031 ;
  wire \u2_Display/n1032 ;
  wire \u2_Display/n1033 ;
  wire \u2_Display/n1034 ;
  wire \u2_Display/n1035 ;
  wire \u2_Display/n1036 ;
  wire \u2_Display/n1037 ;
  wire \u2_Display/n1038 ;
  wire \u2_Display/n1039 ;
  wire \u2_Display/n104 ;
  wire \u2_Display/n1040 ;
  wire \u2_Display/n1041 ;
  wire \u2_Display/n1042 ;
  wire \u2_Display/n1043 ;
  wire \u2_Display/n1044 ;
  wire \u2_Display/n1045 ;
  wire \u2_Display/n1046 ;
  wire \u2_Display/n1047 ;
  wire \u2_Display/n1050 ;
  wire \u2_Display/n1051 ;
  wire \u2_Display/n1052 ;
  wire \u2_Display/n1053 ;
  wire \u2_Display/n1054 ;
  wire \u2_Display/n1055 ;
  wire \u2_Display/n1056 ;
  wire \u2_Display/n1057 ;
  wire \u2_Display/n1058 ;
  wire \u2_Display/n1059 ;
  wire \u2_Display/n1060 ;
  wire \u2_Display/n1061 ;
  wire \u2_Display/n1062 ;
  wire \u2_Display/n1063 ;
  wire \u2_Display/n1064 ;
  wire \u2_Display/n1065 ;
  wire \u2_Display/n1066 ;
  wire \u2_Display/n1067 ;
  wire \u2_Display/n1068 ;
  wire \u2_Display/n1069 ;
  wire \u2_Display/n1070 ;
  wire \u2_Display/n1071 ;
  wire \u2_Display/n1072 ;
  wire \u2_Display/n1073 ;
  wire \u2_Display/n1074 ;
  wire \u2_Display/n1075 ;
  wire \u2_Display/n1076 ;
  wire \u2_Display/n1077 ;
  wire \u2_Display/n1078 ;
  wire \u2_Display/n1079 ;
  wire \u2_Display/n1080 ;
  wire \u2_Display/n1081 ;
  wire \u2_Display/n1082 ;
  wire \u2_Display/n1085 ;
  wire \u2_Display/n1086 ;
  wire \u2_Display/n1087 ;
  wire \u2_Display/n1088 ;
  wire \u2_Display/n1089 ;
  wire \u2_Display/n1090 ;
  wire \u2_Display/n1091 ;
  wire \u2_Display/n1092 ;
  wire \u2_Display/n1093 ;
  wire \u2_Display/n1094 ;
  wire \u2_Display/n1095 ;
  wire \u2_Display/n1096 ;
  wire \u2_Display/n1097 ;
  wire \u2_Display/n1098 ;
  wire \u2_Display/n1099 ;
  wire \u2_Display/n1100 ;
  wire \u2_Display/n1101 ;
  wire \u2_Display/n1102 ;
  wire \u2_Display/n1103 ;
  wire \u2_Display/n1104 ;
  wire \u2_Display/n1105 ;
  wire \u2_Display/n1106 ;
  wire \u2_Display/n1107 ;
  wire \u2_Display/n1108 ;
  wire \u2_Display/n1109 ;
  wire \u2_Display/n1110 ;
  wire \u2_Display/n1111 ;
  wire \u2_Display/n1112 ;
  wire \u2_Display/n1113 ;
  wire \u2_Display/n1114 ;
  wire \u2_Display/n1115 ;
  wire \u2_Display/n1116 ;
  wire \u2_Display/n1117 ;
  wire \u2_Display/n1120 ;
  wire \u2_Display/n1121 ;
  wire \u2_Display/n1122 ;
  wire \u2_Display/n1123 ;
  wire \u2_Display/n1124 ;
  wire \u2_Display/n1125 ;
  wire \u2_Display/n1126 ;
  wire \u2_Display/n1127 ;
  wire \u2_Display/n1128 ;
  wire \u2_Display/n1129 ;
  wire \u2_Display/n1130 ;
  wire \u2_Display/n1131 ;
  wire \u2_Display/n1132 ;
  wire \u2_Display/n1133 ;
  wire \u2_Display/n1134 ;
  wire \u2_Display/n1135 ;
  wire \u2_Display/n1136 ;
  wire \u2_Display/n1137 ;
  wire \u2_Display/n1138 ;
  wire \u2_Display/n1139 ;
  wire \u2_Display/n1140 ;
  wire \u2_Display/n1141 ;
  wire \u2_Display/n1142 ;
  wire \u2_Display/n1143 ;
  wire \u2_Display/n1144 ;
  wire \u2_Display/n1145 ;
  wire \u2_Display/n1146 ;
  wire \u2_Display/n1147 ;
  wire \u2_Display/n1148 ;
  wire \u2_Display/n1149 ;
  wire \u2_Display/n1150 ;
  wire \u2_Display/n1151 ;
  wire \u2_Display/n1152 ;
  wire \u2_Display/n1155 ;
  wire \u2_Display/n1156 ;
  wire \u2_Display/n1157 ;
  wire \u2_Display/n1158 ;
  wire \u2_Display/n1159 ;
  wire \u2_Display/n1160 ;
  wire \u2_Display/n1161 ;
  wire \u2_Display/n1162 ;
  wire \u2_Display/n1163 ;
  wire \u2_Display/n1164 ;
  wire \u2_Display/n1165 ;
  wire \u2_Display/n1166 ;
  wire \u2_Display/n1167 ;
  wire \u2_Display/n1168 ;
  wire \u2_Display/n1169 ;
  wire \u2_Display/n1170 ;
  wire \u2_Display/n1171 ;
  wire \u2_Display/n1172 ;
  wire \u2_Display/n1173 ;
  wire \u2_Display/n1174 ;
  wire \u2_Display/n1175 ;
  wire \u2_Display/n1176 ;
  wire \u2_Display/n1177 ;
  wire \u2_Display/n1178 ;
  wire \u2_Display/n1179 ;
  wire \u2_Display/n1180 ;
  wire \u2_Display/n1181 ;
  wire \u2_Display/n1182 ;
  wire \u2_Display/n1183 ;
  wire \u2_Display/n1184 ;
  wire \u2_Display/n1185 ;
  wire \u2_Display/n1186 ;
  wire \u2_Display/n1187 ;
  wire \u2_Display/n136 ;
  wire \u2_Display/n138 ;
  wire \u2_Display/n141 ;
  wire \u2_Display/n144 ;
  wire \u2_Display/n145 ;
  wire \u2_Display/n1540 ;
  wire \u2_Display/n1543 ;
  wire \u2_Display/n1544 ;
  wire \u2_Display/n1545 ;
  wire \u2_Display/n1546 ;
  wire \u2_Display/n1547 ;
  wire \u2_Display/n1548 ;
  wire \u2_Display/n1549 ;
  wire \u2_Display/n1550 ;
  wire \u2_Display/n1551 ;
  wire \u2_Display/n1552 ;
  wire \u2_Display/n1553 ;
  wire \u2_Display/n1554 ;
  wire \u2_Display/n1555 ;
  wire \u2_Display/n1556 ;
  wire \u2_Display/n1557 ;
  wire \u2_Display/n1558 ;
  wire \u2_Display/n1559 ;
  wire \u2_Display/n1560 ;
  wire \u2_Display/n1561 ;
  wire \u2_Display/n1562 ;
  wire \u2_Display/n1563 ;
  wire \u2_Display/n1564 ;
  wire \u2_Display/n1565 ;
  wire \u2_Display/n1566 ;
  wire \u2_Display/n1567 ;
  wire \u2_Display/n1568 ;
  wire \u2_Display/n1569 ;
  wire \u2_Display/n1570 ;
  wire \u2_Display/n1571 ;
  wire \u2_Display/n1572 ;
  wire \u2_Display/n1573 ;
  wire \u2_Display/n1574 ;
  wire \u2_Display/n1575 ;
  wire \u2_Display/n1578 ;
  wire \u2_Display/n1579 ;
  wire \u2_Display/n1580 ;
  wire \u2_Display/n1581 ;
  wire \u2_Display/n1582 ;
  wire \u2_Display/n1583 ;
  wire \u2_Display/n1584 ;
  wire \u2_Display/n1585 ;
  wire \u2_Display/n1586 ;
  wire \u2_Display/n1587 ;
  wire \u2_Display/n1588 ;
  wire \u2_Display/n1589 ;
  wire \u2_Display/n1590 ;
  wire \u2_Display/n1591 ;
  wire \u2_Display/n1592 ;
  wire \u2_Display/n1593 ;
  wire \u2_Display/n1594 ;
  wire \u2_Display/n1595 ;
  wire \u2_Display/n1596 ;
  wire \u2_Display/n1597 ;
  wire \u2_Display/n1598 ;
  wire \u2_Display/n1599 ;
  wire \u2_Display/n1600 ;
  wire \u2_Display/n1601 ;
  wire \u2_Display/n1602 ;
  wire \u2_Display/n1603 ;
  wire \u2_Display/n1604 ;
  wire \u2_Display/n1605 ;
  wire \u2_Display/n1606 ;
  wire \u2_Display/n1607 ;
  wire \u2_Display/n1608 ;
  wire \u2_Display/n1609 ;
  wire \u2_Display/n1610 ;
  wire \u2_Display/n1613 ;
  wire \u2_Display/n1614 ;
  wire \u2_Display/n1615 ;
  wire \u2_Display/n1616 ;
  wire \u2_Display/n1617 ;
  wire \u2_Display/n1618 ;
  wire \u2_Display/n1619 ;
  wire \u2_Display/n1620 ;
  wire \u2_Display/n1621 ;
  wire \u2_Display/n1622 ;
  wire \u2_Display/n1623 ;
  wire \u2_Display/n1624 ;
  wire \u2_Display/n1625 ;
  wire \u2_Display/n1626 ;
  wire \u2_Display/n1627 ;
  wire \u2_Display/n1628 ;
  wire \u2_Display/n1629 ;
  wire \u2_Display/n1630 ;
  wire \u2_Display/n1631 ;
  wire \u2_Display/n1632 ;
  wire \u2_Display/n1633 ;
  wire \u2_Display/n1634 ;
  wire \u2_Display/n1635 ;
  wire \u2_Display/n1636 ;
  wire \u2_Display/n1637 ;
  wire \u2_Display/n1638 ;
  wire \u2_Display/n1639 ;
  wire \u2_Display/n1640 ;
  wire \u2_Display/n1641 ;
  wire \u2_Display/n1642 ;
  wire \u2_Display/n1643 ;
  wire \u2_Display/n1644 ;
  wire \u2_Display/n1645 ;
  wire \u2_Display/n1648 ;
  wire \u2_Display/n1649 ;
  wire \u2_Display/n1650 ;
  wire \u2_Display/n1651 ;
  wire \u2_Display/n1652 ;
  wire \u2_Display/n1653 ;
  wire \u2_Display/n1654 ;
  wire \u2_Display/n1655 ;
  wire \u2_Display/n1656 ;
  wire \u2_Display/n1657 ;
  wire \u2_Display/n1658 ;
  wire \u2_Display/n1659 ;
  wire \u2_Display/n1660 ;
  wire \u2_Display/n1661 ;
  wire \u2_Display/n1662 ;
  wire \u2_Display/n1663 ;
  wire \u2_Display/n1664 ;
  wire \u2_Display/n1665 ;
  wire \u2_Display/n1666 ;
  wire \u2_Display/n1667 ;
  wire \u2_Display/n1668 ;
  wire \u2_Display/n1669 ;
  wire \u2_Display/n1670 ;
  wire \u2_Display/n1671 ;
  wire \u2_Display/n1672 ;
  wire \u2_Display/n1673 ;
  wire \u2_Display/n1674 ;
  wire \u2_Display/n1675 ;
  wire \u2_Display/n1676 ;
  wire \u2_Display/n1677 ;
  wire \u2_Display/n1678 ;
  wire \u2_Display/n1679 ;
  wire \u2_Display/n1680 ;
  wire \u2_Display/n1683 ;
  wire \u2_Display/n1684 ;
  wire \u2_Display/n1685 ;
  wire \u2_Display/n1686 ;
  wire \u2_Display/n1687 ;
  wire \u2_Display/n1688 ;
  wire \u2_Display/n1689 ;
  wire \u2_Display/n1690 ;
  wire \u2_Display/n1691 ;
  wire \u2_Display/n1692 ;
  wire \u2_Display/n1693 ;
  wire \u2_Display/n1694 ;
  wire \u2_Display/n1695 ;
  wire \u2_Display/n1696 ;
  wire \u2_Display/n1697 ;
  wire \u2_Display/n1698 ;
  wire \u2_Display/n1699 ;
  wire \u2_Display/n1700 ;
  wire \u2_Display/n1701 ;
  wire \u2_Display/n1702 ;
  wire \u2_Display/n1703 ;
  wire \u2_Display/n1704 ;
  wire \u2_Display/n1705 ;
  wire \u2_Display/n1706 ;
  wire \u2_Display/n1707 ;
  wire \u2_Display/n1708 ;
  wire \u2_Display/n1709 ;
  wire \u2_Display/n1710 ;
  wire \u2_Display/n1711 ;
  wire \u2_Display/n1712 ;
  wire \u2_Display/n1713 ;
  wire \u2_Display/n1714 ;
  wire \u2_Display/n1715 ;
  wire \u2_Display/n1718 ;
  wire \u2_Display/n1719 ;
  wire \u2_Display/n1720 ;
  wire \u2_Display/n1721 ;
  wire \u2_Display/n1722 ;
  wire \u2_Display/n1723 ;
  wire \u2_Display/n1724 ;
  wire \u2_Display/n1725 ;
  wire \u2_Display/n1726 ;
  wire \u2_Display/n1727 ;
  wire \u2_Display/n1728 ;
  wire \u2_Display/n1729 ;
  wire \u2_Display/n1730 ;
  wire \u2_Display/n1731 ;
  wire \u2_Display/n1732 ;
  wire \u2_Display/n1733 ;
  wire \u2_Display/n1734 ;
  wire \u2_Display/n1735 ;
  wire \u2_Display/n1736 ;
  wire \u2_Display/n1737 ;
  wire \u2_Display/n1738 ;
  wire \u2_Display/n1739 ;
  wire \u2_Display/n1740 ;
  wire \u2_Display/n1741 ;
  wire \u2_Display/n1742 ;
  wire \u2_Display/n1743 ;
  wire \u2_Display/n1744 ;
  wire \u2_Display/n1745 ;
  wire \u2_Display/n1746 ;
  wire \u2_Display/n1747 ;
  wire \u2_Display/n1748 ;
  wire \u2_Display/n1749 ;
  wire \u2_Display/n1750 ;
  wire \u2_Display/n1753 ;
  wire \u2_Display/n1754 ;
  wire \u2_Display/n1755 ;
  wire \u2_Display/n1756 ;
  wire \u2_Display/n1757 ;
  wire \u2_Display/n1758 ;
  wire \u2_Display/n1759 ;
  wire \u2_Display/n1760 ;
  wire \u2_Display/n1761 ;
  wire \u2_Display/n1762 ;
  wire \u2_Display/n1763 ;
  wire \u2_Display/n1764 ;
  wire \u2_Display/n1765 ;
  wire \u2_Display/n1766 ;
  wire \u2_Display/n1767 ;
  wire \u2_Display/n1768 ;
  wire \u2_Display/n1769 ;
  wire \u2_Display/n1770 ;
  wire \u2_Display/n1771 ;
  wire \u2_Display/n1772 ;
  wire \u2_Display/n1773 ;
  wire \u2_Display/n1774 ;
  wire \u2_Display/n1775 ;
  wire \u2_Display/n1776 ;
  wire \u2_Display/n1777 ;
  wire \u2_Display/n1778 ;
  wire \u2_Display/n1779 ;
  wire \u2_Display/n1780 ;
  wire \u2_Display/n1781 ;
  wire \u2_Display/n1782 ;
  wire \u2_Display/n1783 ;
  wire \u2_Display/n1784 ;
  wire \u2_Display/n1785 ;
  wire \u2_Display/n1788 ;
  wire \u2_Display/n1789 ;
  wire \u2_Display/n1790 ;
  wire \u2_Display/n1791 ;
  wire \u2_Display/n1792 ;
  wire \u2_Display/n1793 ;
  wire \u2_Display/n1794 ;
  wire \u2_Display/n1795 ;
  wire \u2_Display/n1796 ;
  wire \u2_Display/n1797 ;
  wire \u2_Display/n1798 ;
  wire \u2_Display/n1799 ;
  wire \u2_Display/n1800 ;
  wire \u2_Display/n1801 ;
  wire \u2_Display/n1802 ;
  wire \u2_Display/n1803 ;
  wire \u2_Display/n1804 ;
  wire \u2_Display/n1805 ;
  wire \u2_Display/n1806 ;
  wire \u2_Display/n1807 ;
  wire \u2_Display/n1808 ;
  wire \u2_Display/n1809 ;
  wire \u2_Display/n1810 ;
  wire \u2_Display/n1811 ;
  wire \u2_Display/n1812 ;
  wire \u2_Display/n1813 ;
  wire \u2_Display/n1814 ;
  wire \u2_Display/n1815 ;
  wire \u2_Display/n1816 ;
  wire \u2_Display/n1817 ;
  wire \u2_Display/n1818 ;
  wire \u2_Display/n1819 ;
  wire \u2_Display/n1820 ;
  wire \u2_Display/n1823 ;
  wire \u2_Display/n1824 ;
  wire \u2_Display/n1825 ;
  wire \u2_Display/n1826 ;
  wire \u2_Display/n1827 ;
  wire \u2_Display/n1828 ;
  wire \u2_Display/n1829 ;
  wire \u2_Display/n1830 ;
  wire \u2_Display/n1831 ;
  wire \u2_Display/n1832 ;
  wire \u2_Display/n1833 ;
  wire \u2_Display/n1834 ;
  wire \u2_Display/n1835 ;
  wire \u2_Display/n1836 ;
  wire \u2_Display/n1837 ;
  wire \u2_Display/n1838 ;
  wire \u2_Display/n1839 ;
  wire \u2_Display/n1840 ;
  wire \u2_Display/n1841 ;
  wire \u2_Display/n1842 ;
  wire \u2_Display/n1843 ;
  wire \u2_Display/n1844 ;
  wire \u2_Display/n1845 ;
  wire \u2_Display/n1846 ;
  wire \u2_Display/n1847 ;
  wire \u2_Display/n1848 ;
  wire \u2_Display/n1849 ;
  wire \u2_Display/n1850 ;
  wire \u2_Display/n1851 ;
  wire \u2_Display/n1852 ;
  wire \u2_Display/n1853 ;
  wire \u2_Display/n1854 ;
  wire \u2_Display/n1855 ;
  wire \u2_Display/n1858 ;
  wire \u2_Display/n1859 ;
  wire \u2_Display/n1860 ;
  wire \u2_Display/n1861 ;
  wire \u2_Display/n1862 ;
  wire \u2_Display/n1863 ;
  wire \u2_Display/n1864 ;
  wire \u2_Display/n1865 ;
  wire \u2_Display/n1866 ;
  wire \u2_Display/n1867 ;
  wire \u2_Display/n1868 ;
  wire \u2_Display/n1869 ;
  wire \u2_Display/n1870 ;
  wire \u2_Display/n1871 ;
  wire \u2_Display/n1872 ;
  wire \u2_Display/n1873 ;
  wire \u2_Display/n1874 ;
  wire \u2_Display/n1875 ;
  wire \u2_Display/n1876 ;
  wire \u2_Display/n1877 ;
  wire \u2_Display/n1878 ;
  wire \u2_Display/n1879 ;
  wire \u2_Display/n1880 ;
  wire \u2_Display/n1881 ;
  wire \u2_Display/n1882 ;
  wire \u2_Display/n1883 ;
  wire \u2_Display/n1884 ;
  wire \u2_Display/n1885 ;
  wire \u2_Display/n1886 ;
  wire \u2_Display/n1887 ;
  wire \u2_Display/n1888 ;
  wire \u2_Display/n1889 ;
  wire \u2_Display/n1890 ;
  wire \u2_Display/n1893 ;
  wire \u2_Display/n1894 ;
  wire \u2_Display/n1895 ;
  wire \u2_Display/n1896 ;
  wire \u2_Display/n1897 ;
  wire \u2_Display/n1898 ;
  wire \u2_Display/n1899 ;
  wire \u2_Display/n1900 ;
  wire \u2_Display/n1901 ;
  wire \u2_Display/n1902 ;
  wire \u2_Display/n1903 ;
  wire \u2_Display/n1904 ;
  wire \u2_Display/n1905 ;
  wire \u2_Display/n1906 ;
  wire \u2_Display/n1907 ;
  wire \u2_Display/n1908 ;
  wire \u2_Display/n1909 ;
  wire \u2_Display/n1910 ;
  wire \u2_Display/n1911 ;
  wire \u2_Display/n1912 ;
  wire \u2_Display/n1913 ;
  wire \u2_Display/n1914 ;
  wire \u2_Display/n1915 ;
  wire \u2_Display/n1916 ;
  wire \u2_Display/n1917 ;
  wire \u2_Display/n1918 ;
  wire \u2_Display/n1919 ;
  wire \u2_Display/n1920 ;
  wire \u2_Display/n1921 ;
  wire \u2_Display/n1922 ;
  wire \u2_Display/n1923 ;
  wire \u2_Display/n1924 ;
  wire \u2_Display/n1925 ;
  wire \u2_Display/n1928 ;
  wire \u2_Display/n1929 ;
  wire \u2_Display/n1930 ;
  wire \u2_Display/n1931 ;
  wire \u2_Display/n1932 ;
  wire \u2_Display/n1933 ;
  wire \u2_Display/n1934 ;
  wire \u2_Display/n1935 ;
  wire \u2_Display/n1936 ;
  wire \u2_Display/n1937 ;
  wire \u2_Display/n1938 ;
  wire \u2_Display/n1939 ;
  wire \u2_Display/n1940 ;
  wire \u2_Display/n1941 ;
  wire \u2_Display/n1942 ;
  wire \u2_Display/n1943 ;
  wire \u2_Display/n1944 ;
  wire \u2_Display/n1945 ;
  wire \u2_Display/n1946 ;
  wire \u2_Display/n1947 ;
  wire \u2_Display/n1948 ;
  wire \u2_Display/n1949 ;
  wire \u2_Display/n1950 ;
  wire \u2_Display/n1951 ;
  wire \u2_Display/n1952 ;
  wire \u2_Display/n1953 ;
  wire \u2_Display/n1954 ;
  wire \u2_Display/n1955 ;
  wire \u2_Display/n1956 ;
  wire \u2_Display/n1957 ;
  wire \u2_Display/n1958 ;
  wire \u2_Display/n1959 ;
  wire \u2_Display/n1960 ;
  wire \u2_Display/n1963 ;
  wire \u2_Display/n1964 ;
  wire \u2_Display/n1965 ;
  wire \u2_Display/n1966 ;
  wire \u2_Display/n1967 ;
  wire \u2_Display/n1968 ;
  wire \u2_Display/n1969 ;
  wire \u2_Display/n1970 ;
  wire \u2_Display/n1971 ;
  wire \u2_Display/n1972 ;
  wire \u2_Display/n1973 ;
  wire \u2_Display/n1974 ;
  wire \u2_Display/n1975 ;
  wire \u2_Display/n1976 ;
  wire \u2_Display/n1977 ;
  wire \u2_Display/n1978 ;
  wire \u2_Display/n1979 ;
  wire \u2_Display/n1980 ;
  wire \u2_Display/n1981 ;
  wire \u2_Display/n1982 ;
  wire \u2_Display/n1983 ;
  wire \u2_Display/n1984 ;
  wire \u2_Display/n1985 ;
  wire \u2_Display/n1986 ;
  wire \u2_Display/n1987 ;
  wire \u2_Display/n1988 ;
  wire \u2_Display/n1989 ;
  wire \u2_Display/n1990 ;
  wire \u2_Display/n1991 ;
  wire \u2_Display/n1992 ;
  wire \u2_Display/n1993 ;
  wire \u2_Display/n1994 ;
  wire \u2_Display/n1995 ;
  wire \u2_Display/n1998 ;
  wire \u2_Display/n1999 ;
  wire \u2_Display/n2000 ;
  wire \u2_Display/n2001 ;
  wire \u2_Display/n2002 ;
  wire \u2_Display/n2003 ;
  wire \u2_Display/n2004 ;
  wire \u2_Display/n2005 ;
  wire \u2_Display/n2006 ;
  wire \u2_Display/n2007 ;
  wire \u2_Display/n2008 ;
  wire \u2_Display/n2009 ;
  wire \u2_Display/n2010 ;
  wire \u2_Display/n2011 ;
  wire \u2_Display/n2012 ;
  wire \u2_Display/n2013 ;
  wire \u2_Display/n2014 ;
  wire \u2_Display/n2015 ;
  wire \u2_Display/n2016 ;
  wire \u2_Display/n2017 ;
  wire \u2_Display/n2018 ;
  wire \u2_Display/n2019 ;
  wire \u2_Display/n2020 ;
  wire \u2_Display/n2021 ;
  wire \u2_Display/n2022 ;
  wire \u2_Display/n2023 ;
  wire \u2_Display/n2024 ;
  wire \u2_Display/n2025 ;
  wire \u2_Display/n2026 ;
  wire \u2_Display/n2027 ;
  wire \u2_Display/n2028 ;
  wire \u2_Display/n2029 ;
  wire \u2_Display/n2030 ;
  wire \u2_Display/n2033 ;
  wire \u2_Display/n2034 ;
  wire \u2_Display/n2035 ;
  wire \u2_Display/n2036 ;
  wire \u2_Display/n2037 ;
  wire \u2_Display/n2038 ;
  wire \u2_Display/n2039 ;
  wire \u2_Display/n2040 ;
  wire \u2_Display/n2041 ;
  wire \u2_Display/n2042 ;
  wire \u2_Display/n2043 ;
  wire \u2_Display/n2044 ;
  wire \u2_Display/n2045 ;
  wire \u2_Display/n2046 ;
  wire \u2_Display/n2047 ;
  wire \u2_Display/n2048 ;
  wire \u2_Display/n2049 ;
  wire \u2_Display/n2050 ;
  wire \u2_Display/n2051 ;
  wire \u2_Display/n2052 ;
  wire \u2_Display/n2053 ;
  wire \u2_Display/n2054 ;
  wire \u2_Display/n2055 ;
  wire \u2_Display/n2056 ;
  wire \u2_Display/n2057 ;
  wire \u2_Display/n2058 ;
  wire \u2_Display/n2059 ;
  wire \u2_Display/n2060 ;
  wire \u2_Display/n2061 ;
  wire \u2_Display/n2062 ;
  wire \u2_Display/n2063 ;
  wire \u2_Display/n2064 ;
  wire \u2_Display/n2065 ;
  wire \u2_Display/n2068 ;
  wire \u2_Display/n2069 ;
  wire \u2_Display/n2070 ;
  wire \u2_Display/n2071 ;
  wire \u2_Display/n2072 ;
  wire \u2_Display/n2073 ;
  wire \u2_Display/n2074 ;
  wire \u2_Display/n2075 ;
  wire \u2_Display/n2076 ;
  wire \u2_Display/n2077 ;
  wire \u2_Display/n2078 ;
  wire \u2_Display/n2079 ;
  wire \u2_Display/n2080 ;
  wire \u2_Display/n2081 ;
  wire \u2_Display/n2082 ;
  wire \u2_Display/n2083 ;
  wire \u2_Display/n2084 ;
  wire \u2_Display/n2085 ;
  wire \u2_Display/n2086 ;
  wire \u2_Display/n2087 ;
  wire \u2_Display/n2088 ;
  wire \u2_Display/n2089 ;
  wire \u2_Display/n2090 ;
  wire \u2_Display/n2091 ;
  wire \u2_Display/n2092 ;
  wire \u2_Display/n2093 ;
  wire \u2_Display/n2094 ;
  wire \u2_Display/n2095 ;
  wire \u2_Display/n2096 ;
  wire \u2_Display/n2097 ;
  wire \u2_Display/n2098 ;
  wire \u2_Display/n2099 ;
  wire \u2_Display/n2100 ;
  wire \u2_Display/n2103 ;
  wire \u2_Display/n2104 ;
  wire \u2_Display/n2105 ;
  wire \u2_Display/n2106 ;
  wire \u2_Display/n2107 ;
  wire \u2_Display/n2108 ;
  wire \u2_Display/n2109 ;
  wire \u2_Display/n2110 ;
  wire \u2_Display/n2111 ;
  wire \u2_Display/n2112 ;
  wire \u2_Display/n2113 ;
  wire \u2_Display/n2114 ;
  wire \u2_Display/n2115 ;
  wire \u2_Display/n2116 ;
  wire \u2_Display/n2117 ;
  wire \u2_Display/n2118 ;
  wire \u2_Display/n2119 ;
  wire \u2_Display/n2120 ;
  wire \u2_Display/n2121 ;
  wire \u2_Display/n2122 ;
  wire \u2_Display/n2123 ;
  wire \u2_Display/n2124 ;
  wire \u2_Display/n2125 ;
  wire \u2_Display/n2126 ;
  wire \u2_Display/n2127 ;
  wire \u2_Display/n2128 ;
  wire \u2_Display/n2129 ;
  wire \u2_Display/n2130 ;
  wire \u2_Display/n2131 ;
  wire \u2_Display/n2132 ;
  wire \u2_Display/n2133 ;
  wire \u2_Display/n2134 ;
  wire \u2_Display/n2135 ;
  wire \u2_Display/n2138 ;
  wire \u2_Display/n2139 ;
  wire \u2_Display/n2140 ;
  wire \u2_Display/n2141 ;
  wire \u2_Display/n2142 ;
  wire \u2_Display/n2143 ;
  wire \u2_Display/n2144 ;
  wire \u2_Display/n2145 ;
  wire \u2_Display/n2146 ;
  wire \u2_Display/n2147 ;
  wire \u2_Display/n2148 ;
  wire \u2_Display/n2149 ;
  wire \u2_Display/n2150 ;
  wire \u2_Display/n2151 ;
  wire \u2_Display/n2152 ;
  wire \u2_Display/n2153 ;
  wire \u2_Display/n2154 ;
  wire \u2_Display/n2155 ;
  wire \u2_Display/n2156 ;
  wire \u2_Display/n2157 ;
  wire \u2_Display/n2158 ;
  wire \u2_Display/n2159 ;
  wire \u2_Display/n2160 ;
  wire \u2_Display/n2161 ;
  wire \u2_Display/n2162 ;
  wire \u2_Display/n2163 ;
  wire \u2_Display/n2164 ;
  wire \u2_Display/n2165 ;
  wire \u2_Display/n2166 ;
  wire \u2_Display/n2167 ;
  wire \u2_Display/n2168 ;
  wire \u2_Display/n2169 ;
  wire \u2_Display/n2170 ;
  wire \u2_Display/n2173 ;
  wire \u2_Display/n2174 ;
  wire \u2_Display/n2175 ;
  wire \u2_Display/n2176 ;
  wire \u2_Display/n2177 ;
  wire \u2_Display/n2178 ;
  wire \u2_Display/n2179 ;
  wire \u2_Display/n2180 ;
  wire \u2_Display/n2181 ;
  wire \u2_Display/n2182 ;
  wire \u2_Display/n2183 ;
  wire \u2_Display/n2184 ;
  wire \u2_Display/n2185 ;
  wire \u2_Display/n2186 ;
  wire \u2_Display/n2187 ;
  wire \u2_Display/n2188 ;
  wire \u2_Display/n2189 ;
  wire \u2_Display/n2190 ;
  wire \u2_Display/n2191 ;
  wire \u2_Display/n2192 ;
  wire \u2_Display/n2193 ;
  wire \u2_Display/n2194 ;
  wire \u2_Display/n2195 ;
  wire \u2_Display/n2196 ;
  wire \u2_Display/n2197 ;
  wire \u2_Display/n2198 ;
  wire \u2_Display/n2199 ;
  wire \u2_Display/n2200 ;
  wire \u2_Display/n2201 ;
  wire \u2_Display/n2202 ;
  wire \u2_Display/n2203 ;
  wire \u2_Display/n2204 ;
  wire \u2_Display/n2205 ;
  wire \u2_Display/n2208 ;
  wire \u2_Display/n2209 ;
  wire \u2_Display/n2210 ;
  wire \u2_Display/n2211 ;
  wire \u2_Display/n2212 ;
  wire \u2_Display/n2213 ;
  wire \u2_Display/n2214 ;
  wire \u2_Display/n2215 ;
  wire \u2_Display/n2216 ;
  wire \u2_Display/n2217 ;
  wire \u2_Display/n2218 ;
  wire \u2_Display/n2219 ;
  wire \u2_Display/n2220 ;
  wire \u2_Display/n2221 ;
  wire \u2_Display/n2222 ;
  wire \u2_Display/n2223 ;
  wire \u2_Display/n2224 ;
  wire \u2_Display/n2225 ;
  wire \u2_Display/n2226 ;
  wire \u2_Display/n2227 ;
  wire \u2_Display/n2228 ;
  wire \u2_Display/n2229 ;
  wire \u2_Display/n2230 ;
  wire \u2_Display/n2231 ;
  wire \u2_Display/n2232 ;
  wire \u2_Display/n2233 ;
  wire \u2_Display/n2234 ;
  wire \u2_Display/n2235 ;
  wire \u2_Display/n2236 ;
  wire \u2_Display/n2237 ;
  wire \u2_Display/n2238 ;
  wire \u2_Display/n2239 ;
  wire \u2_Display/n2240 ;
  wire \u2_Display/n2243 ;
  wire \u2_Display/n2244 ;
  wire \u2_Display/n2245 ;
  wire \u2_Display/n2246 ;
  wire \u2_Display/n2247 ;
  wire \u2_Display/n2248 ;
  wire \u2_Display/n2249 ;
  wire \u2_Display/n2250 ;
  wire \u2_Display/n2251 ;
  wire \u2_Display/n2252 ;
  wire \u2_Display/n2253 ;
  wire \u2_Display/n2254 ;
  wire \u2_Display/n2255 ;
  wire \u2_Display/n2256 ;
  wire \u2_Display/n2257 ;
  wire \u2_Display/n2258 ;
  wire \u2_Display/n2259 ;
  wire \u2_Display/n2260 ;
  wire \u2_Display/n2261 ;
  wire \u2_Display/n2262 ;
  wire \u2_Display/n2263 ;
  wire \u2_Display/n2264 ;
  wire \u2_Display/n2265 ;
  wire \u2_Display/n2266 ;
  wire \u2_Display/n2267 ;
  wire \u2_Display/n2268 ;
  wire \u2_Display/n2269 ;
  wire \u2_Display/n2270 ;
  wire \u2_Display/n2271 ;
  wire \u2_Display/n2272 ;
  wire \u2_Display/n2273 ;
  wire \u2_Display/n2274 ;
  wire \u2_Display/n2275 ;
  wire \u2_Display/n2278 ;
  wire \u2_Display/n2279 ;
  wire \u2_Display/n2280 ;
  wire \u2_Display/n2281 ;
  wire \u2_Display/n2282 ;
  wire \u2_Display/n2283 ;
  wire \u2_Display/n2284 ;
  wire \u2_Display/n2285 ;
  wire \u2_Display/n2286 ;
  wire \u2_Display/n2287 ;
  wire \u2_Display/n2288 ;
  wire \u2_Display/n2289 ;
  wire \u2_Display/n2290 ;
  wire \u2_Display/n2291 ;
  wire \u2_Display/n2292 ;
  wire \u2_Display/n2293 ;
  wire \u2_Display/n2294 ;
  wire \u2_Display/n2295 ;
  wire \u2_Display/n2296 ;
  wire \u2_Display/n2297 ;
  wire \u2_Display/n2298 ;
  wire \u2_Display/n2299 ;
  wire \u2_Display/n2300 ;
  wire \u2_Display/n2301 ;
  wire \u2_Display/n2302 ;
  wire \u2_Display/n2303 ;
  wire \u2_Display/n2304 ;
  wire \u2_Display/n2305 ;
  wire \u2_Display/n2306 ;
  wire \u2_Display/n2307 ;
  wire \u2_Display/n2308 ;
  wire \u2_Display/n2309 ;
  wire \u2_Display/n2310 ;
  wire \u2_Display/n2663 ;
  wire \u2_Display/n2666 ;
  wire \u2_Display/n2667 ;
  wire \u2_Display/n2668 ;
  wire \u2_Display/n2669 ;
  wire \u2_Display/n2670 ;
  wire \u2_Display/n2671 ;
  wire \u2_Display/n2672 ;
  wire \u2_Display/n2673 ;
  wire \u2_Display/n2674 ;
  wire \u2_Display/n2675 ;
  wire \u2_Display/n2676 ;
  wire \u2_Display/n2677 ;
  wire \u2_Display/n2678 ;
  wire \u2_Display/n2679 ;
  wire \u2_Display/n2680 ;
  wire \u2_Display/n2681 ;
  wire \u2_Display/n2682 ;
  wire \u2_Display/n2683 ;
  wire \u2_Display/n2684 ;
  wire \u2_Display/n2685 ;
  wire \u2_Display/n2686 ;
  wire \u2_Display/n2687 ;
  wire \u2_Display/n2688 ;
  wire \u2_Display/n2689 ;
  wire \u2_Display/n2690 ;
  wire \u2_Display/n2691 ;
  wire \u2_Display/n2692 ;
  wire \u2_Display/n2693 ;
  wire \u2_Display/n2694 ;
  wire \u2_Display/n2695 ;
  wire \u2_Display/n2696 ;
  wire \u2_Display/n2697 ;
  wire \u2_Display/n2698 ;
  wire \u2_Display/n2701 ;
  wire \u2_Display/n2702 ;
  wire \u2_Display/n2703 ;
  wire \u2_Display/n2704 ;
  wire \u2_Display/n2705 ;
  wire \u2_Display/n2706 ;
  wire \u2_Display/n2707 ;
  wire \u2_Display/n2708 ;
  wire \u2_Display/n2709 ;
  wire \u2_Display/n2710 ;
  wire \u2_Display/n2711 ;
  wire \u2_Display/n2712 ;
  wire \u2_Display/n2713 ;
  wire \u2_Display/n2714 ;
  wire \u2_Display/n2715 ;
  wire \u2_Display/n2716 ;
  wire \u2_Display/n2717 ;
  wire \u2_Display/n2718 ;
  wire \u2_Display/n2719 ;
  wire \u2_Display/n2720 ;
  wire \u2_Display/n2721 ;
  wire \u2_Display/n2722 ;
  wire \u2_Display/n2723 ;
  wire \u2_Display/n2724 ;
  wire \u2_Display/n2725 ;
  wire \u2_Display/n2726 ;
  wire \u2_Display/n2727 ;
  wire \u2_Display/n2728 ;
  wire \u2_Display/n2729 ;
  wire \u2_Display/n2730 ;
  wire \u2_Display/n2731 ;
  wire \u2_Display/n2732 ;
  wire \u2_Display/n2733 ;
  wire \u2_Display/n2736 ;
  wire \u2_Display/n2737 ;
  wire \u2_Display/n2738 ;
  wire \u2_Display/n2739 ;
  wire \u2_Display/n2740 ;
  wire \u2_Display/n2741 ;
  wire \u2_Display/n2742 ;
  wire \u2_Display/n2743 ;
  wire \u2_Display/n2744 ;
  wire \u2_Display/n2745 ;
  wire \u2_Display/n2746 ;
  wire \u2_Display/n2747 ;
  wire \u2_Display/n2748 ;
  wire \u2_Display/n2749 ;
  wire \u2_Display/n2750 ;
  wire \u2_Display/n2751 ;
  wire \u2_Display/n2752 ;
  wire \u2_Display/n2753 ;
  wire \u2_Display/n2754 ;
  wire \u2_Display/n2755 ;
  wire \u2_Display/n2756 ;
  wire \u2_Display/n2757 ;
  wire \u2_Display/n2758 ;
  wire \u2_Display/n2759 ;
  wire \u2_Display/n2760 ;
  wire \u2_Display/n2761 ;
  wire \u2_Display/n2762 ;
  wire \u2_Display/n2763 ;
  wire \u2_Display/n2764 ;
  wire \u2_Display/n2765 ;
  wire \u2_Display/n2766 ;
  wire \u2_Display/n2767 ;
  wire \u2_Display/n2768 ;
  wire \u2_Display/n2771 ;
  wire \u2_Display/n2772 ;
  wire \u2_Display/n2773 ;
  wire \u2_Display/n2774 ;
  wire \u2_Display/n2775 ;
  wire \u2_Display/n2776 ;
  wire \u2_Display/n2777 ;
  wire \u2_Display/n2778 ;
  wire \u2_Display/n2779 ;
  wire \u2_Display/n2780 ;
  wire \u2_Display/n2781 ;
  wire \u2_Display/n2782 ;
  wire \u2_Display/n2783 ;
  wire \u2_Display/n2784 ;
  wire \u2_Display/n2785 ;
  wire \u2_Display/n2786 ;
  wire \u2_Display/n2787 ;
  wire \u2_Display/n2788 ;
  wire \u2_Display/n2789 ;
  wire \u2_Display/n2790 ;
  wire \u2_Display/n2791 ;
  wire \u2_Display/n2792 ;
  wire \u2_Display/n2793 ;
  wire \u2_Display/n2794 ;
  wire \u2_Display/n2795 ;
  wire \u2_Display/n2796 ;
  wire \u2_Display/n2797 ;
  wire \u2_Display/n2798 ;
  wire \u2_Display/n2799 ;
  wire \u2_Display/n2800 ;
  wire \u2_Display/n2801 ;
  wire \u2_Display/n2802 ;
  wire \u2_Display/n2803 ;
  wire \u2_Display/n2806 ;
  wire \u2_Display/n2807 ;
  wire \u2_Display/n2808 ;
  wire \u2_Display/n2809 ;
  wire \u2_Display/n2810 ;
  wire \u2_Display/n2811 ;
  wire \u2_Display/n2812 ;
  wire \u2_Display/n2813 ;
  wire \u2_Display/n2814 ;
  wire \u2_Display/n2815 ;
  wire \u2_Display/n2816 ;
  wire \u2_Display/n2817 ;
  wire \u2_Display/n2818 ;
  wire \u2_Display/n2819 ;
  wire \u2_Display/n2820 ;
  wire \u2_Display/n2821 ;
  wire \u2_Display/n2822 ;
  wire \u2_Display/n2823 ;
  wire \u2_Display/n2824 ;
  wire \u2_Display/n2825 ;
  wire \u2_Display/n2826 ;
  wire \u2_Display/n2827 ;
  wire \u2_Display/n2828 ;
  wire \u2_Display/n2829 ;
  wire \u2_Display/n2830 ;
  wire \u2_Display/n2831 ;
  wire \u2_Display/n2832 ;
  wire \u2_Display/n2833 ;
  wire \u2_Display/n2834 ;
  wire \u2_Display/n2835 ;
  wire \u2_Display/n2836 ;
  wire \u2_Display/n2837 ;
  wire \u2_Display/n2838 ;
  wire \u2_Display/n2841 ;
  wire \u2_Display/n2842 ;
  wire \u2_Display/n2843 ;
  wire \u2_Display/n2844 ;
  wire \u2_Display/n2845 ;
  wire \u2_Display/n2846 ;
  wire \u2_Display/n2847 ;
  wire \u2_Display/n2848 ;
  wire \u2_Display/n2849 ;
  wire \u2_Display/n2850 ;
  wire \u2_Display/n2851 ;
  wire \u2_Display/n2852 ;
  wire \u2_Display/n2853 ;
  wire \u2_Display/n2854 ;
  wire \u2_Display/n2855 ;
  wire \u2_Display/n2856 ;
  wire \u2_Display/n2857 ;
  wire \u2_Display/n2858 ;
  wire \u2_Display/n2859 ;
  wire \u2_Display/n2860 ;
  wire \u2_Display/n2861 ;
  wire \u2_Display/n2862 ;
  wire \u2_Display/n2863 ;
  wire \u2_Display/n2864 ;
  wire \u2_Display/n2865 ;
  wire \u2_Display/n2866 ;
  wire \u2_Display/n2867 ;
  wire \u2_Display/n2868 ;
  wire \u2_Display/n2869 ;
  wire \u2_Display/n2870 ;
  wire \u2_Display/n2871 ;
  wire \u2_Display/n2872 ;
  wire \u2_Display/n2873 ;
  wire \u2_Display/n2876 ;
  wire \u2_Display/n2877 ;
  wire \u2_Display/n2878 ;
  wire \u2_Display/n2879 ;
  wire \u2_Display/n2880 ;
  wire \u2_Display/n2881 ;
  wire \u2_Display/n2882 ;
  wire \u2_Display/n2883 ;
  wire \u2_Display/n2884 ;
  wire \u2_Display/n2885 ;
  wire \u2_Display/n2886 ;
  wire \u2_Display/n2887 ;
  wire \u2_Display/n2888 ;
  wire \u2_Display/n2889 ;
  wire \u2_Display/n2890 ;
  wire \u2_Display/n2891 ;
  wire \u2_Display/n2892 ;
  wire \u2_Display/n2893 ;
  wire \u2_Display/n2894 ;
  wire \u2_Display/n2895 ;
  wire \u2_Display/n2896 ;
  wire \u2_Display/n2897 ;
  wire \u2_Display/n2898 ;
  wire \u2_Display/n2899 ;
  wire \u2_Display/n2900 ;
  wire \u2_Display/n2901 ;
  wire \u2_Display/n2902 ;
  wire \u2_Display/n2903 ;
  wire \u2_Display/n2904 ;
  wire \u2_Display/n2905 ;
  wire \u2_Display/n2906 ;
  wire \u2_Display/n2907 ;
  wire \u2_Display/n2908 ;
  wire \u2_Display/n2911 ;
  wire \u2_Display/n2912 ;
  wire \u2_Display/n2913 ;
  wire \u2_Display/n2914 ;
  wire \u2_Display/n2915 ;
  wire \u2_Display/n2916 ;
  wire \u2_Display/n2917 ;
  wire \u2_Display/n2918 ;
  wire \u2_Display/n2919 ;
  wire \u2_Display/n2920 ;
  wire \u2_Display/n2921 ;
  wire \u2_Display/n2922 ;
  wire \u2_Display/n2923 ;
  wire \u2_Display/n2924 ;
  wire \u2_Display/n2925 ;
  wire \u2_Display/n2926 ;
  wire \u2_Display/n2927 ;
  wire \u2_Display/n2928 ;
  wire \u2_Display/n2929 ;
  wire \u2_Display/n2930 ;
  wire \u2_Display/n2931 ;
  wire \u2_Display/n2932 ;
  wire \u2_Display/n2933 ;
  wire \u2_Display/n2934 ;
  wire \u2_Display/n2935 ;
  wire \u2_Display/n2936 ;
  wire \u2_Display/n2937 ;
  wire \u2_Display/n2938 ;
  wire \u2_Display/n2939 ;
  wire \u2_Display/n2940 ;
  wire \u2_Display/n2941 ;
  wire \u2_Display/n2942 ;
  wire \u2_Display/n2943 ;
  wire \u2_Display/n2946 ;
  wire \u2_Display/n2947 ;
  wire \u2_Display/n2948 ;
  wire \u2_Display/n2949 ;
  wire \u2_Display/n2950 ;
  wire \u2_Display/n2951 ;
  wire \u2_Display/n2952 ;
  wire \u2_Display/n2953 ;
  wire \u2_Display/n2954 ;
  wire \u2_Display/n2955 ;
  wire \u2_Display/n2956 ;
  wire \u2_Display/n2957 ;
  wire \u2_Display/n2958 ;
  wire \u2_Display/n2959 ;
  wire \u2_Display/n2960 ;
  wire \u2_Display/n2961 ;
  wire \u2_Display/n2962 ;
  wire \u2_Display/n2963 ;
  wire \u2_Display/n2964 ;
  wire \u2_Display/n2965 ;
  wire \u2_Display/n2966 ;
  wire \u2_Display/n2967 ;
  wire \u2_Display/n2968 ;
  wire \u2_Display/n2969 ;
  wire \u2_Display/n2970 ;
  wire \u2_Display/n2971 ;
  wire \u2_Display/n2972 ;
  wire \u2_Display/n2973 ;
  wire \u2_Display/n2974 ;
  wire \u2_Display/n2975 ;
  wire \u2_Display/n2976 ;
  wire \u2_Display/n2977 ;
  wire \u2_Display/n2978 ;
  wire \u2_Display/n2981 ;
  wire \u2_Display/n2982 ;
  wire \u2_Display/n2983 ;
  wire \u2_Display/n2984 ;
  wire \u2_Display/n2985 ;
  wire \u2_Display/n2986 ;
  wire \u2_Display/n2987 ;
  wire \u2_Display/n2988 ;
  wire \u2_Display/n2989 ;
  wire \u2_Display/n2990 ;
  wire \u2_Display/n2991 ;
  wire \u2_Display/n2992 ;
  wire \u2_Display/n2993 ;
  wire \u2_Display/n2994 ;
  wire \u2_Display/n2995 ;
  wire \u2_Display/n2996 ;
  wire \u2_Display/n2997 ;
  wire \u2_Display/n2998 ;
  wire \u2_Display/n2999 ;
  wire \u2_Display/n3000 ;
  wire \u2_Display/n3001 ;
  wire \u2_Display/n3002 ;
  wire \u2_Display/n3003 ;
  wire \u2_Display/n3004 ;
  wire \u2_Display/n3005 ;
  wire \u2_Display/n3006 ;
  wire \u2_Display/n3007 ;
  wire \u2_Display/n3008 ;
  wire \u2_Display/n3009 ;
  wire \u2_Display/n3010 ;
  wire \u2_Display/n3011 ;
  wire \u2_Display/n3012 ;
  wire \u2_Display/n3013 ;
  wire \u2_Display/n3016 ;
  wire \u2_Display/n3017 ;
  wire \u2_Display/n3018 ;
  wire \u2_Display/n3019 ;
  wire \u2_Display/n3020 ;
  wire \u2_Display/n3021 ;
  wire \u2_Display/n3022 ;
  wire \u2_Display/n3023 ;
  wire \u2_Display/n3024 ;
  wire \u2_Display/n3025 ;
  wire \u2_Display/n3026 ;
  wire \u2_Display/n3027 ;
  wire \u2_Display/n3028 ;
  wire \u2_Display/n3029 ;
  wire \u2_Display/n3030 ;
  wire \u2_Display/n3031 ;
  wire \u2_Display/n3032 ;
  wire \u2_Display/n3033 ;
  wire \u2_Display/n3034 ;
  wire \u2_Display/n3035 ;
  wire \u2_Display/n3036 ;
  wire \u2_Display/n3037 ;
  wire \u2_Display/n3038 ;
  wire \u2_Display/n3039 ;
  wire \u2_Display/n3040 ;
  wire \u2_Display/n3041 ;
  wire \u2_Display/n3042 ;
  wire \u2_Display/n3043 ;
  wire \u2_Display/n3044 ;
  wire \u2_Display/n3045 ;
  wire \u2_Display/n3046 ;
  wire \u2_Display/n3047 ;
  wire \u2_Display/n3048 ;
  wire \u2_Display/n3051 ;
  wire \u2_Display/n3052 ;
  wire \u2_Display/n3053 ;
  wire \u2_Display/n3054 ;
  wire \u2_Display/n3055 ;
  wire \u2_Display/n3056 ;
  wire \u2_Display/n3057 ;
  wire \u2_Display/n3058 ;
  wire \u2_Display/n3059 ;
  wire \u2_Display/n3060 ;
  wire \u2_Display/n3061 ;
  wire \u2_Display/n3062 ;
  wire \u2_Display/n3063 ;
  wire \u2_Display/n3064 ;
  wire \u2_Display/n3065 ;
  wire \u2_Display/n3066 ;
  wire \u2_Display/n3067 ;
  wire \u2_Display/n3068 ;
  wire \u2_Display/n3069 ;
  wire \u2_Display/n3070 ;
  wire \u2_Display/n3071 ;
  wire \u2_Display/n3072 ;
  wire \u2_Display/n3073 ;
  wire \u2_Display/n3074 ;
  wire \u2_Display/n3075 ;
  wire \u2_Display/n3076 ;
  wire \u2_Display/n3077 ;
  wire \u2_Display/n3078 ;
  wire \u2_Display/n3079 ;
  wire \u2_Display/n3080 ;
  wire \u2_Display/n3081 ;
  wire \u2_Display/n3082 ;
  wire \u2_Display/n3083 ;
  wire \u2_Display/n3086 ;
  wire \u2_Display/n3087 ;
  wire \u2_Display/n3088 ;
  wire \u2_Display/n3089 ;
  wire \u2_Display/n3090 ;
  wire \u2_Display/n3091 ;
  wire \u2_Display/n3092 ;
  wire \u2_Display/n3093 ;
  wire \u2_Display/n3094 ;
  wire \u2_Display/n3095 ;
  wire \u2_Display/n3096 ;
  wire \u2_Display/n3097 ;
  wire \u2_Display/n3098 ;
  wire \u2_Display/n3099 ;
  wire \u2_Display/n3100 ;
  wire \u2_Display/n3101 ;
  wire \u2_Display/n3102 ;
  wire \u2_Display/n3103 ;
  wire \u2_Display/n3104 ;
  wire \u2_Display/n3105 ;
  wire \u2_Display/n3106 ;
  wire \u2_Display/n3107 ;
  wire \u2_Display/n3108 ;
  wire \u2_Display/n3109 ;
  wire \u2_Display/n3110 ;
  wire \u2_Display/n3111 ;
  wire \u2_Display/n3112 ;
  wire \u2_Display/n3113 ;
  wire \u2_Display/n3114 ;
  wire \u2_Display/n3115 ;
  wire \u2_Display/n3116 ;
  wire \u2_Display/n3117 ;
  wire \u2_Display/n3118 ;
  wire \u2_Display/n3121 ;
  wire \u2_Display/n3122 ;
  wire \u2_Display/n3123 ;
  wire \u2_Display/n3124 ;
  wire \u2_Display/n3125 ;
  wire \u2_Display/n3126 ;
  wire \u2_Display/n3127 ;
  wire \u2_Display/n3128 ;
  wire \u2_Display/n3129 ;
  wire \u2_Display/n3130 ;
  wire \u2_Display/n3131 ;
  wire \u2_Display/n3132 ;
  wire \u2_Display/n3133 ;
  wire \u2_Display/n3134 ;
  wire \u2_Display/n3135 ;
  wire \u2_Display/n3136 ;
  wire \u2_Display/n3137 ;
  wire \u2_Display/n3138 ;
  wire \u2_Display/n3139 ;
  wire \u2_Display/n3140 ;
  wire \u2_Display/n3141 ;
  wire \u2_Display/n3142 ;
  wire \u2_Display/n3143 ;
  wire \u2_Display/n3144 ;
  wire \u2_Display/n3145 ;
  wire \u2_Display/n3146 ;
  wire \u2_Display/n3147 ;
  wire \u2_Display/n3148 ;
  wire \u2_Display/n3149 ;
  wire \u2_Display/n3150 ;
  wire \u2_Display/n3151 ;
  wire \u2_Display/n3152 ;
  wire \u2_Display/n3153 ;
  wire \u2_Display/n3156 ;
  wire \u2_Display/n3157 ;
  wire \u2_Display/n3158 ;
  wire \u2_Display/n3159 ;
  wire \u2_Display/n3160 ;
  wire \u2_Display/n3161 ;
  wire \u2_Display/n3162 ;
  wire \u2_Display/n3163 ;
  wire \u2_Display/n3164 ;
  wire \u2_Display/n3165 ;
  wire \u2_Display/n3166 ;
  wire \u2_Display/n3167 ;
  wire \u2_Display/n3168 ;
  wire \u2_Display/n3169 ;
  wire \u2_Display/n3170 ;
  wire \u2_Display/n3171 ;
  wire \u2_Display/n3172 ;
  wire \u2_Display/n3173 ;
  wire \u2_Display/n3174 ;
  wire \u2_Display/n3175 ;
  wire \u2_Display/n3176 ;
  wire \u2_Display/n3177 ;
  wire \u2_Display/n3178 ;
  wire \u2_Display/n3179 ;
  wire \u2_Display/n3180 ;
  wire \u2_Display/n3181 ;
  wire \u2_Display/n3182 ;
  wire \u2_Display/n3183 ;
  wire \u2_Display/n3184 ;
  wire \u2_Display/n3185 ;
  wire \u2_Display/n3186 ;
  wire \u2_Display/n3187 ;
  wire \u2_Display/n3188 ;
  wire \u2_Display/n3191 ;
  wire \u2_Display/n3192 ;
  wire \u2_Display/n3193 ;
  wire \u2_Display/n3194 ;
  wire \u2_Display/n3195 ;
  wire \u2_Display/n3196 ;
  wire \u2_Display/n3197 ;
  wire \u2_Display/n3198 ;
  wire \u2_Display/n3199 ;
  wire \u2_Display/n3200 ;
  wire \u2_Display/n3201 ;
  wire \u2_Display/n3202 ;
  wire \u2_Display/n3203 ;
  wire \u2_Display/n3204 ;
  wire \u2_Display/n3205 ;
  wire \u2_Display/n3206 ;
  wire \u2_Display/n3207 ;
  wire \u2_Display/n3208 ;
  wire \u2_Display/n3209 ;
  wire \u2_Display/n3210 ;
  wire \u2_Display/n3211 ;
  wire \u2_Display/n3212 ;
  wire \u2_Display/n3213 ;
  wire \u2_Display/n3214 ;
  wire \u2_Display/n3215 ;
  wire \u2_Display/n3216 ;
  wire \u2_Display/n3217 ;
  wire \u2_Display/n3218 ;
  wire \u2_Display/n3219 ;
  wire \u2_Display/n3220 ;
  wire \u2_Display/n3221 ;
  wire \u2_Display/n3222 ;
  wire \u2_Display/n3223 ;
  wire \u2_Display/n3226 ;
  wire \u2_Display/n3227 ;
  wire \u2_Display/n3228 ;
  wire \u2_Display/n3229 ;
  wire \u2_Display/n3230 ;
  wire \u2_Display/n3231 ;
  wire \u2_Display/n3232 ;
  wire \u2_Display/n3233 ;
  wire \u2_Display/n3234 ;
  wire \u2_Display/n3235 ;
  wire \u2_Display/n3236 ;
  wire \u2_Display/n3237 ;
  wire \u2_Display/n3238 ;
  wire \u2_Display/n3239 ;
  wire \u2_Display/n3240 ;
  wire \u2_Display/n3241 ;
  wire \u2_Display/n3242 ;
  wire \u2_Display/n3243 ;
  wire \u2_Display/n3244 ;
  wire \u2_Display/n3245 ;
  wire \u2_Display/n3246 ;
  wire \u2_Display/n3247 ;
  wire \u2_Display/n3248 ;
  wire \u2_Display/n3249 ;
  wire \u2_Display/n3250 ;
  wire \u2_Display/n3251 ;
  wire \u2_Display/n3252 ;
  wire \u2_Display/n3253 ;
  wire \u2_Display/n3254 ;
  wire \u2_Display/n3255 ;
  wire \u2_Display/n3256 ;
  wire \u2_Display/n3257 ;
  wire \u2_Display/n3258 ;
  wire \u2_Display/n3261 ;
  wire \u2_Display/n3262 ;
  wire \u2_Display/n3263 ;
  wire \u2_Display/n3264 ;
  wire \u2_Display/n3265 ;
  wire \u2_Display/n3266 ;
  wire \u2_Display/n3267 ;
  wire \u2_Display/n3268 ;
  wire \u2_Display/n3269 ;
  wire \u2_Display/n3270 ;
  wire \u2_Display/n3271 ;
  wire \u2_Display/n3272 ;
  wire \u2_Display/n3273 ;
  wire \u2_Display/n3274 ;
  wire \u2_Display/n3275 ;
  wire \u2_Display/n3276 ;
  wire \u2_Display/n3277 ;
  wire \u2_Display/n3278 ;
  wire \u2_Display/n3279 ;
  wire \u2_Display/n3280 ;
  wire \u2_Display/n3281 ;
  wire \u2_Display/n3282 ;
  wire \u2_Display/n3283 ;
  wire \u2_Display/n3284 ;
  wire \u2_Display/n3285 ;
  wire \u2_Display/n3286 ;
  wire \u2_Display/n3287 ;
  wire \u2_Display/n3288 ;
  wire \u2_Display/n3289 ;
  wire \u2_Display/n3290 ;
  wire \u2_Display/n3291 ;
  wire \u2_Display/n3292 ;
  wire \u2_Display/n3293 ;
  wire \u2_Display/n3296 ;
  wire \u2_Display/n3297 ;
  wire \u2_Display/n3298 ;
  wire \u2_Display/n3299 ;
  wire \u2_Display/n3300 ;
  wire \u2_Display/n3301 ;
  wire \u2_Display/n3302 ;
  wire \u2_Display/n3303 ;
  wire \u2_Display/n3304 ;
  wire \u2_Display/n3305 ;
  wire \u2_Display/n3306 ;
  wire \u2_Display/n3307 ;
  wire \u2_Display/n3308 ;
  wire \u2_Display/n3309 ;
  wire \u2_Display/n3310 ;
  wire \u2_Display/n3311 ;
  wire \u2_Display/n3312 ;
  wire \u2_Display/n3313 ;
  wire \u2_Display/n3314 ;
  wire \u2_Display/n3315 ;
  wire \u2_Display/n3316 ;
  wire \u2_Display/n3317 ;
  wire \u2_Display/n3318 ;
  wire \u2_Display/n3319 ;
  wire \u2_Display/n3320 ;
  wire \u2_Display/n3321 ;
  wire \u2_Display/n3322 ;
  wire \u2_Display/n3323 ;
  wire \u2_Display/n3324 ;
  wire \u2_Display/n3325 ;
  wire \u2_Display/n3326 ;
  wire \u2_Display/n3327 ;
  wire \u2_Display/n3328 ;
  wire \u2_Display/n3331 ;
  wire \u2_Display/n3332 ;
  wire \u2_Display/n3333 ;
  wire \u2_Display/n3334 ;
  wire \u2_Display/n3335 ;
  wire \u2_Display/n3336 ;
  wire \u2_Display/n3337 ;
  wire \u2_Display/n3338 ;
  wire \u2_Display/n3339 ;
  wire \u2_Display/n3340 ;
  wire \u2_Display/n3341 ;
  wire \u2_Display/n3342 ;
  wire \u2_Display/n3343 ;
  wire \u2_Display/n3344 ;
  wire \u2_Display/n3345 ;
  wire \u2_Display/n3346 ;
  wire \u2_Display/n3347 ;
  wire \u2_Display/n3348 ;
  wire \u2_Display/n3349 ;
  wire \u2_Display/n3350 ;
  wire \u2_Display/n3351 ;
  wire \u2_Display/n3352 ;
  wire \u2_Display/n3353 ;
  wire \u2_Display/n3354 ;
  wire \u2_Display/n3355 ;
  wire \u2_Display/n3356 ;
  wire \u2_Display/n3357 ;
  wire \u2_Display/n3358 ;
  wire \u2_Display/n3359 ;
  wire \u2_Display/n3360 ;
  wire \u2_Display/n3361 ;
  wire \u2_Display/n3362 ;
  wire \u2_Display/n3363 ;
  wire \u2_Display/n3366 ;
  wire \u2_Display/n3367 ;
  wire \u2_Display/n3368 ;
  wire \u2_Display/n3369 ;
  wire \u2_Display/n3370 ;
  wire \u2_Display/n3371 ;
  wire \u2_Display/n3372 ;
  wire \u2_Display/n3373 ;
  wire \u2_Display/n3374 ;
  wire \u2_Display/n3375 ;
  wire \u2_Display/n3376 ;
  wire \u2_Display/n3377 ;
  wire \u2_Display/n3378 ;
  wire \u2_Display/n3379 ;
  wire \u2_Display/n3380 ;
  wire \u2_Display/n3381 ;
  wire \u2_Display/n3382 ;
  wire \u2_Display/n3383 ;
  wire \u2_Display/n3384 ;
  wire \u2_Display/n3385 ;
  wire \u2_Display/n3386 ;
  wire \u2_Display/n3387 ;
  wire \u2_Display/n3388 ;
  wire \u2_Display/n3389 ;
  wire \u2_Display/n3390 ;
  wire \u2_Display/n3391 ;
  wire \u2_Display/n3392 ;
  wire \u2_Display/n3393 ;
  wire \u2_Display/n3394 ;
  wire \u2_Display/n3395 ;
  wire \u2_Display/n3396 ;
  wire \u2_Display/n3397 ;
  wire \u2_Display/n3398 ;
  wire \u2_Display/n3401 ;
  wire \u2_Display/n3402 ;
  wire \u2_Display/n3403 ;
  wire \u2_Display/n3404 ;
  wire \u2_Display/n3405 ;
  wire \u2_Display/n3406 ;
  wire \u2_Display/n3407 ;
  wire \u2_Display/n3408 ;
  wire \u2_Display/n3409 ;
  wire \u2_Display/n3410 ;
  wire \u2_Display/n3411 ;
  wire \u2_Display/n3412 ;
  wire \u2_Display/n3413 ;
  wire \u2_Display/n3414 ;
  wire \u2_Display/n3415 ;
  wire \u2_Display/n3416 ;
  wire \u2_Display/n3417 ;
  wire \u2_Display/n3418 ;
  wire \u2_Display/n3419 ;
  wire \u2_Display/n3420 ;
  wire \u2_Display/n3421 ;
  wire \u2_Display/n3422 ;
  wire \u2_Display/n3423 ;
  wire \u2_Display/n3424 ;
  wire \u2_Display/n3425 ;
  wire \u2_Display/n3426 ;
  wire \u2_Display/n3427 ;
  wire \u2_Display/n3428 ;
  wire \u2_Display/n3429 ;
  wire \u2_Display/n3430 ;
  wire \u2_Display/n3431 ;
  wire \u2_Display/n3432 ;
  wire \u2_Display/n3433 ;
  wire \u2_Display/n35 ;
  wire \u2_Display/n36 ;
  wire \u2_Display/n3786 ;
  wire \u2_Display/n3789 ;
  wire \u2_Display/n3790 ;
  wire \u2_Display/n3791 ;
  wire \u2_Display/n3792 ;
  wire \u2_Display/n3793 ;
  wire \u2_Display/n3794 ;
  wire \u2_Display/n3795 ;
  wire \u2_Display/n3796 ;
  wire \u2_Display/n3797 ;
  wire \u2_Display/n3798 ;
  wire \u2_Display/n3799 ;
  wire \u2_Display/n3800 ;
  wire \u2_Display/n3801 ;
  wire \u2_Display/n3802 ;
  wire \u2_Display/n3803 ;
  wire \u2_Display/n3804 ;
  wire \u2_Display/n3805 ;
  wire \u2_Display/n3806 ;
  wire \u2_Display/n3807 ;
  wire \u2_Display/n3808 ;
  wire \u2_Display/n3809 ;
  wire \u2_Display/n3810 ;
  wire \u2_Display/n3811 ;
  wire \u2_Display/n3812 ;
  wire \u2_Display/n3813 ;
  wire \u2_Display/n3814 ;
  wire \u2_Display/n3815 ;
  wire \u2_Display/n3816 ;
  wire \u2_Display/n3817 ;
  wire \u2_Display/n3818 ;
  wire \u2_Display/n3819 ;
  wire \u2_Display/n3820 ;
  wire \u2_Display/n3821 ;
  wire \u2_Display/n3824 ;
  wire \u2_Display/n3825 ;
  wire \u2_Display/n3826 ;
  wire \u2_Display/n3827 ;
  wire \u2_Display/n3828 ;
  wire \u2_Display/n3829 ;
  wire \u2_Display/n3830 ;
  wire \u2_Display/n3831 ;
  wire \u2_Display/n3832 ;
  wire \u2_Display/n3833 ;
  wire \u2_Display/n3834 ;
  wire \u2_Display/n3835 ;
  wire \u2_Display/n3836 ;
  wire \u2_Display/n3837 ;
  wire \u2_Display/n3838 ;
  wire \u2_Display/n3839 ;
  wire \u2_Display/n3840 ;
  wire \u2_Display/n3841 ;
  wire \u2_Display/n3842 ;
  wire \u2_Display/n3843 ;
  wire \u2_Display/n3844 ;
  wire \u2_Display/n3845 ;
  wire \u2_Display/n3846 ;
  wire \u2_Display/n3847 ;
  wire \u2_Display/n3848 ;
  wire \u2_Display/n3849 ;
  wire \u2_Display/n3850 ;
  wire \u2_Display/n3851 ;
  wire \u2_Display/n3852 ;
  wire \u2_Display/n3853 ;
  wire \u2_Display/n3854 ;
  wire \u2_Display/n3855 ;
  wire \u2_Display/n3856 ;
  wire \u2_Display/n3859 ;
  wire \u2_Display/n3860 ;
  wire \u2_Display/n3861 ;
  wire \u2_Display/n3862 ;
  wire \u2_Display/n3863 ;
  wire \u2_Display/n3864 ;
  wire \u2_Display/n3865 ;
  wire \u2_Display/n3866 ;
  wire \u2_Display/n3867 ;
  wire \u2_Display/n3868 ;
  wire \u2_Display/n3869 ;
  wire \u2_Display/n3870 ;
  wire \u2_Display/n3871 ;
  wire \u2_Display/n3872 ;
  wire \u2_Display/n3873 ;
  wire \u2_Display/n3874 ;
  wire \u2_Display/n3875 ;
  wire \u2_Display/n3876 ;
  wire \u2_Display/n3877 ;
  wire \u2_Display/n3878 ;
  wire \u2_Display/n3879 ;
  wire \u2_Display/n3880 ;
  wire \u2_Display/n3881 ;
  wire \u2_Display/n3882 ;
  wire \u2_Display/n3883 ;
  wire \u2_Display/n3884 ;
  wire \u2_Display/n3885 ;
  wire \u2_Display/n3886 ;
  wire \u2_Display/n3887 ;
  wire \u2_Display/n3888 ;
  wire \u2_Display/n3889 ;
  wire \u2_Display/n3890 ;
  wire \u2_Display/n3891 ;
  wire \u2_Display/n3894 ;
  wire \u2_Display/n3895 ;
  wire \u2_Display/n3896 ;
  wire \u2_Display/n3897 ;
  wire \u2_Display/n3898 ;
  wire \u2_Display/n3899 ;
  wire \u2_Display/n3900 ;
  wire \u2_Display/n3901 ;
  wire \u2_Display/n3902 ;
  wire \u2_Display/n3903 ;
  wire \u2_Display/n3904 ;
  wire \u2_Display/n3905 ;
  wire \u2_Display/n3906 ;
  wire \u2_Display/n3907 ;
  wire \u2_Display/n3908 ;
  wire \u2_Display/n3909 ;
  wire \u2_Display/n3910 ;
  wire \u2_Display/n3911 ;
  wire \u2_Display/n3912 ;
  wire \u2_Display/n3913 ;
  wire \u2_Display/n3914 ;
  wire \u2_Display/n3915 ;
  wire \u2_Display/n3916 ;
  wire \u2_Display/n3917 ;
  wire \u2_Display/n3918 ;
  wire \u2_Display/n3919 ;
  wire \u2_Display/n3920 ;
  wire \u2_Display/n3921 ;
  wire \u2_Display/n3922 ;
  wire \u2_Display/n3923 ;
  wire \u2_Display/n3924 ;
  wire \u2_Display/n3925 ;
  wire \u2_Display/n3926 ;
  wire \u2_Display/n3929 ;
  wire \u2_Display/n3930 ;
  wire \u2_Display/n3931 ;
  wire \u2_Display/n3932 ;
  wire \u2_Display/n3933 ;
  wire \u2_Display/n3934 ;
  wire \u2_Display/n3935 ;
  wire \u2_Display/n3936 ;
  wire \u2_Display/n3937 ;
  wire \u2_Display/n3938 ;
  wire \u2_Display/n3939 ;
  wire \u2_Display/n3940 ;
  wire \u2_Display/n3941 ;
  wire \u2_Display/n3942 ;
  wire \u2_Display/n3943 ;
  wire \u2_Display/n3944 ;
  wire \u2_Display/n3945 ;
  wire \u2_Display/n3946 ;
  wire \u2_Display/n3947 ;
  wire \u2_Display/n3948 ;
  wire \u2_Display/n3949 ;
  wire \u2_Display/n3950 ;
  wire \u2_Display/n3951 ;
  wire \u2_Display/n3952 ;
  wire \u2_Display/n3953 ;
  wire \u2_Display/n3954 ;
  wire \u2_Display/n3955 ;
  wire \u2_Display/n3956 ;
  wire \u2_Display/n3957 ;
  wire \u2_Display/n3958 ;
  wire \u2_Display/n3959 ;
  wire \u2_Display/n3960 ;
  wire \u2_Display/n3961 ;
  wire \u2_Display/n3964 ;
  wire \u2_Display/n3965 ;
  wire \u2_Display/n3966 ;
  wire \u2_Display/n3967 ;
  wire \u2_Display/n3968 ;
  wire \u2_Display/n3969 ;
  wire \u2_Display/n3970 ;
  wire \u2_Display/n3971 ;
  wire \u2_Display/n3972 ;
  wire \u2_Display/n3973 ;
  wire \u2_Display/n3974 ;
  wire \u2_Display/n3975 ;
  wire \u2_Display/n3976 ;
  wire \u2_Display/n3977 ;
  wire \u2_Display/n3978 ;
  wire \u2_Display/n3979 ;
  wire \u2_Display/n3980 ;
  wire \u2_Display/n3981 ;
  wire \u2_Display/n3982 ;
  wire \u2_Display/n3983 ;
  wire \u2_Display/n3984 ;
  wire \u2_Display/n3985 ;
  wire \u2_Display/n3986 ;
  wire \u2_Display/n3987 ;
  wire \u2_Display/n3988 ;
  wire \u2_Display/n3989 ;
  wire \u2_Display/n3990 ;
  wire \u2_Display/n3991 ;
  wire \u2_Display/n3992 ;
  wire \u2_Display/n3993 ;
  wire \u2_Display/n3994 ;
  wire \u2_Display/n3995 ;
  wire \u2_Display/n3996 ;
  wire \u2_Display/n3999 ;
  wire \u2_Display/n4000 ;
  wire \u2_Display/n4001 ;
  wire \u2_Display/n4002 ;
  wire \u2_Display/n4003 ;
  wire \u2_Display/n4004 ;
  wire \u2_Display/n4005 ;
  wire \u2_Display/n4006 ;
  wire \u2_Display/n4007 ;
  wire \u2_Display/n4008 ;
  wire \u2_Display/n4009 ;
  wire \u2_Display/n4010 ;
  wire \u2_Display/n4011 ;
  wire \u2_Display/n4012 ;
  wire \u2_Display/n4013 ;
  wire \u2_Display/n4014 ;
  wire \u2_Display/n4015 ;
  wire \u2_Display/n4016 ;
  wire \u2_Display/n4017 ;
  wire \u2_Display/n4018 ;
  wire \u2_Display/n4019 ;
  wire \u2_Display/n4020 ;
  wire \u2_Display/n4021 ;
  wire \u2_Display/n4022 ;
  wire \u2_Display/n4023 ;
  wire \u2_Display/n4024 ;
  wire \u2_Display/n4025 ;
  wire \u2_Display/n4026 ;
  wire \u2_Display/n4027 ;
  wire \u2_Display/n4028 ;
  wire \u2_Display/n4029 ;
  wire \u2_Display/n4030 ;
  wire \u2_Display/n4031 ;
  wire \u2_Display/n4034 ;
  wire \u2_Display/n4035 ;
  wire \u2_Display/n4036 ;
  wire \u2_Display/n4037 ;
  wire \u2_Display/n4038 ;
  wire \u2_Display/n4039 ;
  wire \u2_Display/n4040 ;
  wire \u2_Display/n4041 ;
  wire \u2_Display/n4042 ;
  wire \u2_Display/n4043 ;
  wire \u2_Display/n4044 ;
  wire \u2_Display/n4045 ;
  wire \u2_Display/n4046 ;
  wire \u2_Display/n4047 ;
  wire \u2_Display/n4048 ;
  wire \u2_Display/n4049 ;
  wire \u2_Display/n4050 ;
  wire \u2_Display/n4051 ;
  wire \u2_Display/n4052 ;
  wire \u2_Display/n4053 ;
  wire \u2_Display/n4054 ;
  wire \u2_Display/n4055 ;
  wire \u2_Display/n4056 ;
  wire \u2_Display/n4057 ;
  wire \u2_Display/n4058 ;
  wire \u2_Display/n4059 ;
  wire \u2_Display/n4060 ;
  wire \u2_Display/n4061 ;
  wire \u2_Display/n4062 ;
  wire \u2_Display/n4063 ;
  wire \u2_Display/n4064 ;
  wire \u2_Display/n4065 ;
  wire \u2_Display/n4066 ;
  wire \u2_Display/n4069 ;
  wire \u2_Display/n4070 ;
  wire \u2_Display/n4071 ;
  wire \u2_Display/n4072 ;
  wire \u2_Display/n4073 ;
  wire \u2_Display/n4074 ;
  wire \u2_Display/n4075 ;
  wire \u2_Display/n4076 ;
  wire \u2_Display/n4077 ;
  wire \u2_Display/n4078 ;
  wire \u2_Display/n4079 ;
  wire \u2_Display/n4080 ;
  wire \u2_Display/n4081 ;
  wire \u2_Display/n4082 ;
  wire \u2_Display/n4083 ;
  wire \u2_Display/n4084 ;
  wire \u2_Display/n4085 ;
  wire \u2_Display/n4086 ;
  wire \u2_Display/n4087 ;
  wire \u2_Display/n4088 ;
  wire \u2_Display/n4089 ;
  wire \u2_Display/n4090 ;
  wire \u2_Display/n4091 ;
  wire \u2_Display/n4092 ;
  wire \u2_Display/n4093 ;
  wire \u2_Display/n4094 ;
  wire \u2_Display/n4095 ;
  wire \u2_Display/n4096 ;
  wire \u2_Display/n4097 ;
  wire \u2_Display/n4098 ;
  wire \u2_Display/n4099 ;
  wire \u2_Display/n4100 ;
  wire \u2_Display/n4101 ;
  wire \u2_Display/n4104 ;
  wire \u2_Display/n4105 ;
  wire \u2_Display/n4106 ;
  wire \u2_Display/n4107 ;
  wire \u2_Display/n4108 ;
  wire \u2_Display/n4109 ;
  wire \u2_Display/n4110 ;
  wire \u2_Display/n4111 ;
  wire \u2_Display/n4112 ;
  wire \u2_Display/n4113 ;
  wire \u2_Display/n4114 ;
  wire \u2_Display/n4115 ;
  wire \u2_Display/n4116 ;
  wire \u2_Display/n4117 ;
  wire \u2_Display/n4118 ;
  wire \u2_Display/n4119 ;
  wire \u2_Display/n4120 ;
  wire \u2_Display/n4121 ;
  wire \u2_Display/n4122 ;
  wire \u2_Display/n4123 ;
  wire \u2_Display/n4124 ;
  wire \u2_Display/n4125 ;
  wire \u2_Display/n4126 ;
  wire \u2_Display/n4127 ;
  wire \u2_Display/n4128 ;
  wire \u2_Display/n4129 ;
  wire \u2_Display/n4130 ;
  wire \u2_Display/n4131 ;
  wire \u2_Display/n4132 ;
  wire \u2_Display/n4133 ;
  wire \u2_Display/n4134 ;
  wire \u2_Display/n4135 ;
  wire \u2_Display/n4136 ;
  wire \u2_Display/n4139 ;
  wire \u2_Display/n4140 ;
  wire \u2_Display/n4141 ;
  wire \u2_Display/n4142 ;
  wire \u2_Display/n4143 ;
  wire \u2_Display/n4144 ;
  wire \u2_Display/n4145 ;
  wire \u2_Display/n4146 ;
  wire \u2_Display/n4147 ;
  wire \u2_Display/n4148 ;
  wire \u2_Display/n4149 ;
  wire \u2_Display/n4150 ;
  wire \u2_Display/n4151 ;
  wire \u2_Display/n4152 ;
  wire \u2_Display/n4153 ;
  wire \u2_Display/n4154 ;
  wire \u2_Display/n4155 ;
  wire \u2_Display/n4156 ;
  wire \u2_Display/n4157 ;
  wire \u2_Display/n4158 ;
  wire \u2_Display/n4159 ;
  wire \u2_Display/n4160 ;
  wire \u2_Display/n4161 ;
  wire \u2_Display/n4162 ;
  wire \u2_Display/n4163 ;
  wire \u2_Display/n4164 ;
  wire \u2_Display/n4165 ;
  wire \u2_Display/n4166 ;
  wire \u2_Display/n4167 ;
  wire \u2_Display/n4168 ;
  wire \u2_Display/n4169 ;
  wire \u2_Display/n417 ;
  wire \u2_Display/n4170 ;
  wire \u2_Display/n4171 ;
  wire \u2_Display/n4174 ;
  wire \u2_Display/n4175 ;
  wire \u2_Display/n4176 ;
  wire \u2_Display/n4177 ;
  wire \u2_Display/n4178 ;
  wire \u2_Display/n4179 ;
  wire \u2_Display/n4180 ;
  wire \u2_Display/n4181 ;
  wire \u2_Display/n4182 ;
  wire \u2_Display/n4183 ;
  wire \u2_Display/n4184 ;
  wire \u2_Display/n4185 ;
  wire \u2_Display/n4186 ;
  wire \u2_Display/n4187 ;
  wire \u2_Display/n4188 ;
  wire \u2_Display/n4189 ;
  wire \u2_Display/n4190 ;
  wire \u2_Display/n4191 ;
  wire \u2_Display/n4192 ;
  wire \u2_Display/n4193 ;
  wire \u2_Display/n4194 ;
  wire \u2_Display/n4195 ;
  wire \u2_Display/n4196 ;
  wire \u2_Display/n4197 ;
  wire \u2_Display/n4198 ;
  wire \u2_Display/n4199 ;
  wire \u2_Display/n420 ;
  wire \u2_Display/n4200 ;
  wire \u2_Display/n4201 ;
  wire \u2_Display/n4202 ;
  wire \u2_Display/n4203 ;
  wire \u2_Display/n4204 ;
  wire \u2_Display/n4205 ;
  wire \u2_Display/n4206 ;
  wire \u2_Display/n4209 ;
  wire \u2_Display/n421 ;
  wire \u2_Display/n4210 ;
  wire \u2_Display/n4211 ;
  wire \u2_Display/n4212 ;
  wire \u2_Display/n4213 ;
  wire \u2_Display/n4214 ;
  wire \u2_Display/n4215 ;
  wire \u2_Display/n4216 ;
  wire \u2_Display/n4217 ;
  wire \u2_Display/n4218 ;
  wire \u2_Display/n4219 ;
  wire \u2_Display/n422 ;
  wire \u2_Display/n4220 ;
  wire \u2_Display/n4221 ;
  wire \u2_Display/n4222 ;
  wire \u2_Display/n4223 ;
  wire \u2_Display/n4224 ;
  wire \u2_Display/n4225 ;
  wire \u2_Display/n4226 ;
  wire \u2_Display/n4227 ;
  wire \u2_Display/n4228 ;
  wire \u2_Display/n4229 ;
  wire \u2_Display/n423 ;
  wire \u2_Display/n4230 ;
  wire \u2_Display/n4231 ;
  wire \u2_Display/n4232 ;
  wire \u2_Display/n4233 ;
  wire \u2_Display/n4234 ;
  wire \u2_Display/n4235 ;
  wire \u2_Display/n4236 ;
  wire \u2_Display/n4237 ;
  wire \u2_Display/n4238 ;
  wire \u2_Display/n4239 ;
  wire \u2_Display/n424 ;
  wire \u2_Display/n4240 ;
  wire \u2_Display/n4241 ;
  wire \u2_Display/n4244 ;
  wire \u2_Display/n4245 ;
  wire \u2_Display/n4246 ;
  wire \u2_Display/n4247 ;
  wire \u2_Display/n4248 ;
  wire \u2_Display/n4249 ;
  wire \u2_Display/n425 ;
  wire \u2_Display/n4250 ;
  wire \u2_Display/n4251 ;
  wire \u2_Display/n4252 ;
  wire \u2_Display/n4253 ;
  wire \u2_Display/n4254 ;
  wire \u2_Display/n4255 ;
  wire \u2_Display/n4256 ;
  wire \u2_Display/n4257 ;
  wire \u2_Display/n4258 ;
  wire \u2_Display/n4259 ;
  wire \u2_Display/n426 ;
  wire \u2_Display/n4260 ;
  wire \u2_Display/n4261 ;
  wire \u2_Display/n4262 ;
  wire \u2_Display/n4263 ;
  wire \u2_Display/n4264 ;
  wire \u2_Display/n4265 ;
  wire \u2_Display/n4266 ;
  wire \u2_Display/n4267 ;
  wire \u2_Display/n4268 ;
  wire \u2_Display/n4269 ;
  wire \u2_Display/n427 ;
  wire \u2_Display/n4270 ;
  wire \u2_Display/n4271 ;
  wire \u2_Display/n4272 ;
  wire \u2_Display/n4273 ;
  wire \u2_Display/n4274 ;
  wire \u2_Display/n4275 ;
  wire \u2_Display/n4276 ;
  wire \u2_Display/n4279 ;
  wire \u2_Display/n428 ;
  wire \u2_Display/n4280 ;
  wire \u2_Display/n4281 ;
  wire \u2_Display/n4282 ;
  wire \u2_Display/n4283 ;
  wire \u2_Display/n4284 ;
  wire \u2_Display/n4285 ;
  wire \u2_Display/n4286 ;
  wire \u2_Display/n4287 ;
  wire \u2_Display/n4288 ;
  wire \u2_Display/n4289 ;
  wire \u2_Display/n429 ;
  wire \u2_Display/n4290 ;
  wire \u2_Display/n4291 ;
  wire \u2_Display/n4292 ;
  wire \u2_Display/n4293 ;
  wire \u2_Display/n4294 ;
  wire \u2_Display/n4295 ;
  wire \u2_Display/n4296 ;
  wire \u2_Display/n4297 ;
  wire \u2_Display/n4298 ;
  wire \u2_Display/n4299 ;
  wire \u2_Display/n430 ;
  wire \u2_Display/n4300 ;
  wire \u2_Display/n4301 ;
  wire \u2_Display/n4302 ;
  wire \u2_Display/n4303 ;
  wire \u2_Display/n4304 ;
  wire \u2_Display/n4305 ;
  wire \u2_Display/n4306 ;
  wire \u2_Display/n4307 ;
  wire \u2_Display/n4308 ;
  wire \u2_Display/n4309 ;
  wire \u2_Display/n431 ;
  wire \u2_Display/n4310 ;
  wire \u2_Display/n4311 ;
  wire \u2_Display/n4314 ;
  wire \u2_Display/n4315 ;
  wire \u2_Display/n4316 ;
  wire \u2_Display/n4317 ;
  wire \u2_Display/n4318 ;
  wire \u2_Display/n4319 ;
  wire \u2_Display/n432 ;
  wire \u2_Display/n4320 ;
  wire \u2_Display/n4321 ;
  wire \u2_Display/n4322 ;
  wire \u2_Display/n4323 ;
  wire \u2_Display/n4324 ;
  wire \u2_Display/n4325 ;
  wire \u2_Display/n4326 ;
  wire \u2_Display/n4327 ;
  wire \u2_Display/n4328 ;
  wire \u2_Display/n4329 ;
  wire \u2_Display/n433 ;
  wire \u2_Display/n4330 ;
  wire \u2_Display/n4331 ;
  wire \u2_Display/n4332 ;
  wire \u2_Display/n4333 ;
  wire \u2_Display/n4334 ;
  wire \u2_Display/n4335 ;
  wire \u2_Display/n4336 ;
  wire \u2_Display/n4337 ;
  wire \u2_Display/n4338 ;
  wire \u2_Display/n4339 ;
  wire \u2_Display/n434 ;
  wire \u2_Display/n4340 ;
  wire \u2_Display/n4341 ;
  wire \u2_Display/n4342 ;
  wire \u2_Display/n4343 ;
  wire \u2_Display/n4344 ;
  wire \u2_Display/n4345 ;
  wire \u2_Display/n4346 ;
  wire \u2_Display/n4349 ;
  wire \u2_Display/n435 ;
  wire \u2_Display/n4350 ;
  wire \u2_Display/n4351 ;
  wire \u2_Display/n4352 ;
  wire \u2_Display/n4353 ;
  wire \u2_Display/n4354 ;
  wire \u2_Display/n4355 ;
  wire \u2_Display/n4356 ;
  wire \u2_Display/n4357 ;
  wire \u2_Display/n4358 ;
  wire \u2_Display/n4359 ;
  wire \u2_Display/n436 ;
  wire \u2_Display/n4360 ;
  wire \u2_Display/n4361 ;
  wire \u2_Display/n4362 ;
  wire \u2_Display/n4363 ;
  wire \u2_Display/n4364 ;
  wire \u2_Display/n4365 ;
  wire \u2_Display/n4366 ;
  wire \u2_Display/n4367 ;
  wire \u2_Display/n4368 ;
  wire \u2_Display/n4369 ;
  wire \u2_Display/n437 ;
  wire \u2_Display/n4370 ;
  wire \u2_Display/n4371 ;
  wire \u2_Display/n4372 ;
  wire \u2_Display/n4373 ;
  wire \u2_Display/n4374 ;
  wire \u2_Display/n4375 ;
  wire \u2_Display/n4376 ;
  wire \u2_Display/n4377 ;
  wire \u2_Display/n4378 ;
  wire \u2_Display/n4379 ;
  wire \u2_Display/n438 ;
  wire \u2_Display/n4380 ;
  wire \u2_Display/n4381 ;
  wire \u2_Display/n4384 ;
  wire \u2_Display/n4385 ;
  wire \u2_Display/n4386 ;
  wire \u2_Display/n4387 ;
  wire \u2_Display/n4388 ;
  wire \u2_Display/n4389 ;
  wire \u2_Display/n439 ;
  wire \u2_Display/n4390 ;
  wire \u2_Display/n4391 ;
  wire \u2_Display/n4392 ;
  wire \u2_Display/n4393 ;
  wire \u2_Display/n4394 ;
  wire \u2_Display/n4395 ;
  wire \u2_Display/n4396 ;
  wire \u2_Display/n4397 ;
  wire \u2_Display/n4398 ;
  wire \u2_Display/n4399 ;
  wire \u2_Display/n44 ;
  wire \u2_Display/n440 ;
  wire \u2_Display/n4400 ;
  wire \u2_Display/n4401 ;
  wire \u2_Display/n4402 ;
  wire \u2_Display/n4403 ;
  wire \u2_Display/n4404 ;
  wire \u2_Display/n4405 ;
  wire \u2_Display/n4406 ;
  wire \u2_Display/n4407 ;
  wire \u2_Display/n4408 ;
  wire \u2_Display/n4409 ;
  wire \u2_Display/n441 ;
  wire \u2_Display/n4410 ;
  wire \u2_Display/n4411 ;
  wire \u2_Display/n4412 ;
  wire \u2_Display/n4413 ;
  wire \u2_Display/n4414 ;
  wire \u2_Display/n4415 ;
  wire \u2_Display/n4416 ;
  wire \u2_Display/n4419 ;
  wire \u2_Display/n442 ;
  wire \u2_Display/n4420 ;
  wire \u2_Display/n4421 ;
  wire \u2_Display/n4422 ;
  wire \u2_Display/n4423 ;
  wire \u2_Display/n4424 ;
  wire \u2_Display/n4425 ;
  wire \u2_Display/n4426 ;
  wire \u2_Display/n4427 ;
  wire \u2_Display/n4428 ;
  wire \u2_Display/n4429 ;
  wire \u2_Display/n443 ;
  wire \u2_Display/n4430 ;
  wire \u2_Display/n4431 ;
  wire \u2_Display/n4432 ;
  wire \u2_Display/n4433 ;
  wire \u2_Display/n4434 ;
  wire \u2_Display/n4435 ;
  wire \u2_Display/n4436 ;
  wire \u2_Display/n4437 ;
  wire \u2_Display/n4438 ;
  wire \u2_Display/n4439 ;
  wire \u2_Display/n444 ;
  wire \u2_Display/n4440 ;
  wire \u2_Display/n4441 ;
  wire \u2_Display/n4442 ;
  wire \u2_Display/n4443 ;
  wire \u2_Display/n4444 ;
  wire \u2_Display/n4445 ;
  wire \u2_Display/n4446 ;
  wire \u2_Display/n4447 ;
  wire \u2_Display/n4448 ;
  wire \u2_Display/n4449 ;
  wire \u2_Display/n445 ;
  wire \u2_Display/n4450 ;
  wire \u2_Display/n4451 ;
  wire \u2_Display/n4454 ;
  wire \u2_Display/n4455 ;
  wire \u2_Display/n4456 ;
  wire \u2_Display/n4457 ;
  wire \u2_Display/n4458 ;
  wire \u2_Display/n4459 ;
  wire \u2_Display/n446 ;
  wire \u2_Display/n4460 ;
  wire \u2_Display/n4461 ;
  wire \u2_Display/n4462 ;
  wire \u2_Display/n4463 ;
  wire \u2_Display/n4464 ;
  wire \u2_Display/n4465 ;
  wire \u2_Display/n4466 ;
  wire \u2_Display/n4467 ;
  wire \u2_Display/n4468 ;
  wire \u2_Display/n4469 ;
  wire \u2_Display/n447 ;
  wire \u2_Display/n4470 ;
  wire \u2_Display/n4471 ;
  wire \u2_Display/n4472 ;
  wire \u2_Display/n4473 ;
  wire \u2_Display/n4474 ;
  wire \u2_Display/n4475 ;
  wire \u2_Display/n4476 ;
  wire \u2_Display/n4477 ;
  wire \u2_Display/n4478 ;
  wire \u2_Display/n4479 ;
  wire \u2_Display/n448 ;
  wire \u2_Display/n4480 ;
  wire \u2_Display/n4481 ;
  wire \u2_Display/n4482 ;
  wire \u2_Display/n4483 ;
  wire \u2_Display/n4484 ;
  wire \u2_Display/n4485 ;
  wire \u2_Display/n4486 ;
  wire \u2_Display/n4489 ;
  wire \u2_Display/n449 ;
  wire \u2_Display/n4490 ;
  wire \u2_Display/n4491 ;
  wire \u2_Display/n4492 ;
  wire \u2_Display/n4493 ;
  wire \u2_Display/n4494 ;
  wire \u2_Display/n4495 ;
  wire \u2_Display/n4496 ;
  wire \u2_Display/n4497 ;
  wire \u2_Display/n4498 ;
  wire \u2_Display/n4499 ;
  wire \u2_Display/n45 ;
  wire \u2_Display/n450 ;
  wire \u2_Display/n4500 ;
  wire \u2_Display/n4501 ;
  wire \u2_Display/n4502 ;
  wire \u2_Display/n4503 ;
  wire \u2_Display/n4504 ;
  wire \u2_Display/n4505 ;
  wire \u2_Display/n4506 ;
  wire \u2_Display/n4507 ;
  wire \u2_Display/n4508 ;
  wire \u2_Display/n4509 ;
  wire \u2_Display/n451 ;
  wire \u2_Display/n4510 ;
  wire \u2_Display/n4511 ;
  wire \u2_Display/n4512 ;
  wire \u2_Display/n4513 ;
  wire \u2_Display/n4514 ;
  wire \u2_Display/n4515 ;
  wire \u2_Display/n4516 ;
  wire \u2_Display/n4517 ;
  wire \u2_Display/n4518 ;
  wire \u2_Display/n4519 ;
  wire \u2_Display/n452 ;
  wire \u2_Display/n4520 ;
  wire \u2_Display/n4521 ;
  wire \u2_Display/n4524 ;
  wire \u2_Display/n4525 ;
  wire \u2_Display/n4526 ;
  wire \u2_Display/n4527 ;
  wire \u2_Display/n4528 ;
  wire \u2_Display/n4529 ;
  wire \u2_Display/n4530 ;
  wire \u2_Display/n4531 ;
  wire \u2_Display/n4532 ;
  wire \u2_Display/n4533 ;
  wire \u2_Display/n4534 ;
  wire \u2_Display/n4535 ;
  wire \u2_Display/n4536 ;
  wire \u2_Display/n4537 ;
  wire \u2_Display/n4538 ;
  wire \u2_Display/n4539 ;
  wire \u2_Display/n4540 ;
  wire \u2_Display/n4541 ;
  wire \u2_Display/n4542 ;
  wire \u2_Display/n4543 ;
  wire \u2_Display/n4544 ;
  wire \u2_Display/n4545 ;
  wire \u2_Display/n4546 ;
  wire \u2_Display/n4547 ;
  wire \u2_Display/n4548 ;
  wire \u2_Display/n4549 ;
  wire \u2_Display/n455 ;
  wire \u2_Display/n4550 ;
  wire \u2_Display/n4551 ;
  wire \u2_Display/n4552 ;
  wire \u2_Display/n4553 ;
  wire \u2_Display/n4554 ;
  wire \u2_Display/n4555 ;
  wire \u2_Display/n4556 ;
  wire \u2_Display/n456 ;
  wire \u2_Display/n457 ;
  wire \u2_Display/n458 ;
  wire \u2_Display/n459 ;
  wire \u2_Display/n460 ;
  wire \u2_Display/n461 ;
  wire \u2_Display/n462 ;
  wire \u2_Display/n463 ;
  wire \u2_Display/n464 ;
  wire \u2_Display/n465 ;
  wire \u2_Display/n466 ;
  wire \u2_Display/n467 ;
  wire \u2_Display/n468 ;
  wire \u2_Display/n469 ;
  wire \u2_Display/n470 ;
  wire \u2_Display/n471 ;
  wire \u2_Display/n472 ;
  wire \u2_Display/n473 ;
  wire \u2_Display/n474 ;
  wire \u2_Display/n475 ;
  wire \u2_Display/n476 ;
  wire \u2_Display/n477 ;
  wire \u2_Display/n478 ;
  wire \u2_Display/n479 ;
  wire \u2_Display/n48 ;
  wire \u2_Display/n480 ;
  wire \u2_Display/n481 ;
  wire \u2_Display/n482 ;
  wire \u2_Display/n483 ;
  wire \u2_Display/n484 ;
  wire \u2_Display/n485 ;
  wire \u2_Display/n486 ;
  wire \u2_Display/n487 ;
  wire \u2_Display/n490 ;
  wire \u2_Display/n4909 ;
  wire \u2_Display/n491 ;
  wire \u2_Display/n492 ;
  wire \u2_Display/n493 ;
  wire \u2_Display/n494 ;
  wire \u2_Display/n4944 ;
  wire \u2_Display/n495 ;
  wire \u2_Display/n496 ;
  wire \u2_Display/n497 ;
  wire \u2_Display/n4979 ;
  wire \u2_Display/n498 ;
  wire \u2_Display/n499 ;
  wire \u2_Display/n50 ;
  wire \u2_Display/n500 ;
  wire \u2_Display/n501 ;
  wire \u2_Display/n5014 ;
  wire \u2_Display/n502 ;
  wire \u2_Display/n503 ;
  wire \u2_Display/n504 ;
  wire \u2_Display/n5049 ;
  wire \u2_Display/n505 ;
  wire \u2_Display/n506 ;
  wire \u2_Display/n507 ;
  wire \u2_Display/n508 ;
  wire \u2_Display/n5084 ;
  wire \u2_Display/n509 ;
  wire \u2_Display/n51 ;
  wire \u2_Display/n510 ;
  wire \u2_Display/n511 ;
  wire \u2_Display/n5119 ;
  wire \u2_Display/n512 ;
  wire \u2_Display/n513 ;
  wire \u2_Display/n514 ;
  wire \u2_Display/n515 ;
  wire \u2_Display/n5154 ;
  wire \u2_Display/n516 ;
  wire \u2_Display/n517 ;
  wire \u2_Display/n518 ;
  wire \u2_Display/n5189 ;
  wire \u2_Display/n519 ;
  wire \u2_Display/n5196 ;
  wire \u2_Display/n5197 ;
  wire \u2_Display/n5198 ;
  wire \u2_Display/n5199 ;
  wire \u2_Display/n520 ;
  wire \u2_Display/n5200 ;
  wire \u2_Display/n5201 ;
  wire \u2_Display/n5202 ;
  wire \u2_Display/n5203 ;
  wire \u2_Display/n5204 ;
  wire \u2_Display/n5205 ;
  wire \u2_Display/n5206 ;
  wire \u2_Display/n5207 ;
  wire \u2_Display/n5208 ;
  wire \u2_Display/n5209 ;
  wire \u2_Display/n521 ;
  wire \u2_Display/n5210 ;
  wire \u2_Display/n5211 ;
  wire \u2_Display/n5212 ;
  wire \u2_Display/n5213 ;
  wire \u2_Display/n5214 ;
  wire \u2_Display/n5215 ;
  wire \u2_Display/n5216 ;
  wire \u2_Display/n5217 ;
  wire \u2_Display/n5218 ;
  wire \u2_Display/n5219 ;
  wire \u2_Display/n522 ;
  wire \u2_Display/n5220 ;
  wire \u2_Display/n5221 ;
  wire \u2_Display/n5222 ;
  wire \u2_Display/n5223 ;
  wire \u2_Display/n5224 ;
  wire \u2_Display/n5227 ;
  wire \u2_Display/n5228 ;
  wire \u2_Display/n5229 ;
  wire \u2_Display/n5230 ;
  wire \u2_Display/n5231 ;
  wire \u2_Display/n5232 ;
  wire \u2_Display/n5233 ;
  wire \u2_Display/n5234 ;
  wire \u2_Display/n5235 ;
  wire \u2_Display/n5236 ;
  wire \u2_Display/n5237 ;
  wire \u2_Display/n5238 ;
  wire \u2_Display/n5239 ;
  wire \u2_Display/n5240 ;
  wire \u2_Display/n5241 ;
  wire \u2_Display/n5242 ;
  wire \u2_Display/n5243 ;
  wire \u2_Display/n5244 ;
  wire \u2_Display/n5245 ;
  wire \u2_Display/n5246 ;
  wire \u2_Display/n5247 ;
  wire \u2_Display/n5248 ;
  wire \u2_Display/n5249 ;
  wire \u2_Display/n525 ;
  wire \u2_Display/n5250 ;
  wire \u2_Display/n5251 ;
  wire \u2_Display/n5252 ;
  wire \u2_Display/n5253 ;
  wire \u2_Display/n5254 ;
  wire \u2_Display/n5255 ;
  wire \u2_Display/n5256 ;
  wire \u2_Display/n5257 ;
  wire \u2_Display/n5258 ;
  wire \u2_Display/n5259 ;
  wire \u2_Display/n526 ;
  wire \u2_Display/n5262 ;
  wire \u2_Display/n5263 ;
  wire \u2_Display/n5264 ;
  wire \u2_Display/n5265 ;
  wire \u2_Display/n5266 ;
  wire \u2_Display/n5267 ;
  wire \u2_Display/n5268 ;
  wire \u2_Display/n5269 ;
  wire \u2_Display/n527 ;
  wire \u2_Display/n5270 ;
  wire \u2_Display/n5271 ;
  wire \u2_Display/n5272 ;
  wire \u2_Display/n5273 ;
  wire \u2_Display/n5274 ;
  wire \u2_Display/n5275 ;
  wire \u2_Display/n5276 ;
  wire \u2_Display/n5277 ;
  wire \u2_Display/n5278 ;
  wire \u2_Display/n5279 ;
  wire \u2_Display/n528 ;
  wire \u2_Display/n5280 ;
  wire \u2_Display/n5281 ;
  wire \u2_Display/n5282 ;
  wire \u2_Display/n5283 ;
  wire \u2_Display/n5284 ;
  wire \u2_Display/n5285 ;
  wire \u2_Display/n5286 ;
  wire \u2_Display/n5287 ;
  wire \u2_Display/n5288 ;
  wire \u2_Display/n5289 ;
  wire \u2_Display/n529 ;
  wire \u2_Display/n5290 ;
  wire \u2_Display/n5291 ;
  wire \u2_Display/n5292 ;
  wire \u2_Display/n5293 ;
  wire \u2_Display/n5294 ;
  wire \u2_Display/n5297 ;
  wire \u2_Display/n5298 ;
  wire \u2_Display/n5299 ;
  wire \u2_Display/n530 ;
  wire \u2_Display/n5300 ;
  wire \u2_Display/n5301 ;
  wire \u2_Display/n5302 ;
  wire \u2_Display/n5303 ;
  wire \u2_Display/n5304 ;
  wire \u2_Display/n5305 ;
  wire \u2_Display/n5306 ;
  wire \u2_Display/n5307 ;
  wire \u2_Display/n5308 ;
  wire \u2_Display/n5309 ;
  wire \u2_Display/n531 ;
  wire \u2_Display/n5310 ;
  wire \u2_Display/n5311 ;
  wire \u2_Display/n5312 ;
  wire \u2_Display/n5313 ;
  wire \u2_Display/n5314 ;
  wire \u2_Display/n5315 ;
  wire \u2_Display/n5316 ;
  wire \u2_Display/n5317 ;
  wire \u2_Display/n5318 ;
  wire \u2_Display/n5319 ;
  wire \u2_Display/n532 ;
  wire \u2_Display/n5320 ;
  wire \u2_Display/n5321 ;
  wire \u2_Display/n5322 ;
  wire \u2_Display/n5323 ;
  wire \u2_Display/n5324 ;
  wire \u2_Display/n5325 ;
  wire \u2_Display/n5326 ;
  wire \u2_Display/n5327 ;
  wire \u2_Display/n5328 ;
  wire \u2_Display/n5329 ;
  wire \u2_Display/n533 ;
  wire \u2_Display/n5332 ;
  wire \u2_Display/n5333 ;
  wire \u2_Display/n5334 ;
  wire \u2_Display/n5335 ;
  wire \u2_Display/n5336 ;
  wire \u2_Display/n5337 ;
  wire \u2_Display/n5338 ;
  wire \u2_Display/n5339 ;
  wire \u2_Display/n534 ;
  wire \u2_Display/n5340 ;
  wire \u2_Display/n5341 ;
  wire \u2_Display/n5342 ;
  wire \u2_Display/n5343 ;
  wire \u2_Display/n5344 ;
  wire \u2_Display/n5345 ;
  wire \u2_Display/n5346 ;
  wire \u2_Display/n5347 ;
  wire \u2_Display/n5348 ;
  wire \u2_Display/n5349 ;
  wire \u2_Display/n535 ;
  wire \u2_Display/n5350 ;
  wire \u2_Display/n5351 ;
  wire \u2_Display/n5352 ;
  wire \u2_Display/n5353 ;
  wire \u2_Display/n5354 ;
  wire \u2_Display/n5355 ;
  wire \u2_Display/n5356 ;
  wire \u2_Display/n5357 ;
  wire \u2_Display/n5358 ;
  wire \u2_Display/n5359 ;
  wire \u2_Display/n536 ;
  wire \u2_Display/n5360 ;
  wire \u2_Display/n5361 ;
  wire \u2_Display/n5362 ;
  wire \u2_Display/n5363 ;
  wire \u2_Display/n5364 ;
  wire \u2_Display/n5367 ;
  wire \u2_Display/n5368 ;
  wire \u2_Display/n5369 ;
  wire \u2_Display/n537 ;
  wire \u2_Display/n5370 ;
  wire \u2_Display/n5371 ;
  wire \u2_Display/n5372 ;
  wire \u2_Display/n5373 ;
  wire \u2_Display/n5374 ;
  wire \u2_Display/n5375 ;
  wire \u2_Display/n5376 ;
  wire \u2_Display/n5377 ;
  wire \u2_Display/n5378 ;
  wire \u2_Display/n5379 ;
  wire \u2_Display/n538 ;
  wire \u2_Display/n5380 ;
  wire \u2_Display/n5381 ;
  wire \u2_Display/n5382 ;
  wire \u2_Display/n5383 ;
  wire \u2_Display/n5384 ;
  wire \u2_Display/n5385 ;
  wire \u2_Display/n5386 ;
  wire \u2_Display/n5387 ;
  wire \u2_Display/n5388 ;
  wire \u2_Display/n5389 ;
  wire \u2_Display/n539 ;
  wire \u2_Display/n5390 ;
  wire \u2_Display/n5391 ;
  wire \u2_Display/n5392 ;
  wire \u2_Display/n5393 ;
  wire \u2_Display/n5394 ;
  wire \u2_Display/n5395 ;
  wire \u2_Display/n5396 ;
  wire \u2_Display/n5397 ;
  wire \u2_Display/n5398 ;
  wire \u2_Display/n5399 ;
  wire \u2_Display/n540 ;
  wire \u2_Display/n5402 ;
  wire \u2_Display/n5403 ;
  wire \u2_Display/n5404 ;
  wire \u2_Display/n5405 ;
  wire \u2_Display/n5406 ;
  wire \u2_Display/n5407 ;
  wire \u2_Display/n5408 ;
  wire \u2_Display/n5409 ;
  wire \u2_Display/n541 ;
  wire \u2_Display/n5410 ;
  wire \u2_Display/n5411 ;
  wire \u2_Display/n5412 ;
  wire \u2_Display/n5413 ;
  wire \u2_Display/n5414 ;
  wire \u2_Display/n5415 ;
  wire \u2_Display/n5416 ;
  wire \u2_Display/n5417 ;
  wire \u2_Display/n5418 ;
  wire \u2_Display/n5419 ;
  wire \u2_Display/n542 ;
  wire \u2_Display/n5420 ;
  wire \u2_Display/n5421 ;
  wire \u2_Display/n5422 ;
  wire \u2_Display/n5423 ;
  wire \u2_Display/n5424 ;
  wire \u2_Display/n5425 ;
  wire \u2_Display/n5426 ;
  wire \u2_Display/n5427 ;
  wire \u2_Display/n5428 ;
  wire \u2_Display/n5429 ;
  wire \u2_Display/n543 ;
  wire \u2_Display/n5430 ;
  wire \u2_Display/n5431 ;
  wire \u2_Display/n5432 ;
  wire \u2_Display/n5433 ;
  wire \u2_Display/n5434 ;
  wire \u2_Display/n5437 ;
  wire \u2_Display/n5438 ;
  wire \u2_Display/n5439 ;
  wire \u2_Display/n544 ;
  wire \u2_Display/n5440 ;
  wire \u2_Display/n5441 ;
  wire \u2_Display/n5442 ;
  wire \u2_Display/n5443 ;
  wire \u2_Display/n5444 ;
  wire \u2_Display/n5445 ;
  wire \u2_Display/n5446 ;
  wire \u2_Display/n5447 ;
  wire \u2_Display/n5448 ;
  wire \u2_Display/n5449 ;
  wire \u2_Display/n545 ;
  wire \u2_Display/n5450 ;
  wire \u2_Display/n5451 ;
  wire \u2_Display/n5452 ;
  wire \u2_Display/n5453 ;
  wire \u2_Display/n5454 ;
  wire \u2_Display/n5455 ;
  wire \u2_Display/n5456 ;
  wire \u2_Display/n5457 ;
  wire \u2_Display/n5458 ;
  wire \u2_Display/n5459 ;
  wire \u2_Display/n546 ;
  wire \u2_Display/n5460 ;
  wire \u2_Display/n5461 ;
  wire \u2_Display/n5462 ;
  wire \u2_Display/n5463 ;
  wire \u2_Display/n5464 ;
  wire \u2_Display/n5465 ;
  wire \u2_Display/n5466 ;
  wire \u2_Display/n5467 ;
  wire \u2_Display/n5468 ;
  wire \u2_Display/n5469 ;
  wire \u2_Display/n547 ;
  wire \u2_Display/n5472 ;
  wire \u2_Display/n5473 ;
  wire \u2_Display/n5474 ;
  wire \u2_Display/n5475 ;
  wire \u2_Display/n5476 ;
  wire \u2_Display/n5477 ;
  wire \u2_Display/n5478 ;
  wire \u2_Display/n5479 ;
  wire \u2_Display/n548 ;
  wire \u2_Display/n5480 ;
  wire \u2_Display/n5481 ;
  wire \u2_Display/n5482 ;
  wire \u2_Display/n5483 ;
  wire \u2_Display/n5484 ;
  wire \u2_Display/n5485 ;
  wire \u2_Display/n5486 ;
  wire \u2_Display/n5487 ;
  wire \u2_Display/n5488 ;
  wire \u2_Display/n5489 ;
  wire \u2_Display/n549 ;
  wire \u2_Display/n5490 ;
  wire \u2_Display/n5491 ;
  wire \u2_Display/n5492 ;
  wire \u2_Display/n5493 ;
  wire \u2_Display/n5494 ;
  wire \u2_Display/n5495 ;
  wire \u2_Display/n5496 ;
  wire \u2_Display/n5497 ;
  wire \u2_Display/n5498 ;
  wire \u2_Display/n5499 ;
  wire \u2_Display/n550 ;
  wire \u2_Display/n5500 ;
  wire \u2_Display/n5501 ;
  wire \u2_Display/n5502 ;
  wire \u2_Display/n5503 ;
  wire \u2_Display/n5504 ;
  wire \u2_Display/n5507 ;
  wire \u2_Display/n5508 ;
  wire \u2_Display/n5509 ;
  wire \u2_Display/n551 ;
  wire \u2_Display/n5510 ;
  wire \u2_Display/n5511 ;
  wire \u2_Display/n5512 ;
  wire \u2_Display/n5513 ;
  wire \u2_Display/n5514 ;
  wire \u2_Display/n5515 ;
  wire \u2_Display/n5516 ;
  wire \u2_Display/n5517 ;
  wire \u2_Display/n5518 ;
  wire \u2_Display/n5519 ;
  wire \u2_Display/n552 ;
  wire \u2_Display/n5520 ;
  wire \u2_Display/n5521 ;
  wire \u2_Display/n5522 ;
  wire \u2_Display/n5523 ;
  wire \u2_Display/n5524 ;
  wire \u2_Display/n5525 ;
  wire \u2_Display/n5526 ;
  wire \u2_Display/n5527 ;
  wire \u2_Display/n5528 ;
  wire \u2_Display/n5529 ;
  wire \u2_Display/n553 ;
  wire \u2_Display/n5530 ;
  wire \u2_Display/n5531 ;
  wire \u2_Display/n5532 ;
  wire \u2_Display/n5533 ;
  wire \u2_Display/n5534 ;
  wire \u2_Display/n5535 ;
  wire \u2_Display/n5536 ;
  wire \u2_Display/n5537 ;
  wire \u2_Display/n5538 ;
  wire \u2_Display/n5539 ;
  wire \u2_Display/n554 ;
  wire \u2_Display/n5542 ;
  wire \u2_Display/n5543 ;
  wire \u2_Display/n5544 ;
  wire \u2_Display/n5545 ;
  wire \u2_Display/n5546 ;
  wire \u2_Display/n5547 ;
  wire \u2_Display/n5548 ;
  wire \u2_Display/n5549 ;
  wire \u2_Display/n555 ;
  wire \u2_Display/n5550 ;
  wire \u2_Display/n5551 ;
  wire \u2_Display/n5552 ;
  wire \u2_Display/n5553 ;
  wire \u2_Display/n5554 ;
  wire \u2_Display/n5555 ;
  wire \u2_Display/n5556 ;
  wire \u2_Display/n5557 ;
  wire \u2_Display/n5558 ;
  wire \u2_Display/n5559 ;
  wire \u2_Display/n556 ;
  wire \u2_Display/n5560 ;
  wire \u2_Display/n5561 ;
  wire \u2_Display/n5562 ;
  wire \u2_Display/n5563 ;
  wire \u2_Display/n5564 ;
  wire \u2_Display/n5565 ;
  wire \u2_Display/n5566 ;
  wire \u2_Display/n5567 ;
  wire \u2_Display/n5568 ;
  wire \u2_Display/n5569 ;
  wire \u2_Display/n557 ;
  wire \u2_Display/n5570 ;
  wire \u2_Display/n5571 ;
  wire \u2_Display/n5572 ;
  wire \u2_Display/n5573 ;
  wire \u2_Display/n5574 ;
  wire \u2_Display/n5577 ;
  wire \u2_Display/n5578 ;
  wire \u2_Display/n5579 ;
  wire \u2_Display/n5580 ;
  wire \u2_Display/n5581 ;
  wire \u2_Display/n5582 ;
  wire \u2_Display/n5583 ;
  wire \u2_Display/n5584 ;
  wire \u2_Display/n5585 ;
  wire \u2_Display/n5586 ;
  wire \u2_Display/n5587 ;
  wire \u2_Display/n5588 ;
  wire \u2_Display/n5589 ;
  wire \u2_Display/n5590 ;
  wire \u2_Display/n5591 ;
  wire \u2_Display/n5592 ;
  wire \u2_Display/n5593 ;
  wire \u2_Display/n5594 ;
  wire \u2_Display/n5595 ;
  wire \u2_Display/n5596 ;
  wire \u2_Display/n5597 ;
  wire \u2_Display/n5598 ;
  wire \u2_Display/n5599 ;
  wire \u2_Display/n560 ;
  wire \u2_Display/n5600 ;
  wire \u2_Display/n5601 ;
  wire \u2_Display/n5602 ;
  wire \u2_Display/n5603 ;
  wire \u2_Display/n5604 ;
  wire \u2_Display/n5605 ;
  wire \u2_Display/n5606 ;
  wire \u2_Display/n5607 ;
  wire \u2_Display/n5608 ;
  wire \u2_Display/n5609 ;
  wire \u2_Display/n561 ;
  wire \u2_Display/n5612 ;
  wire \u2_Display/n5613 ;
  wire \u2_Display/n5614 ;
  wire \u2_Display/n5615 ;
  wire \u2_Display/n5616 ;
  wire \u2_Display/n5617 ;
  wire \u2_Display/n5618 ;
  wire \u2_Display/n5619 ;
  wire \u2_Display/n562 ;
  wire \u2_Display/n5620 ;
  wire \u2_Display/n5621 ;
  wire \u2_Display/n5622 ;
  wire \u2_Display/n5623 ;
  wire \u2_Display/n5624 ;
  wire \u2_Display/n5625 ;
  wire \u2_Display/n5626 ;
  wire \u2_Display/n5627 ;
  wire \u2_Display/n5628 ;
  wire \u2_Display/n5629 ;
  wire \u2_Display/n563 ;
  wire \u2_Display/n5630 ;
  wire \u2_Display/n5631 ;
  wire \u2_Display/n5632 ;
  wire \u2_Display/n5633 ;
  wire \u2_Display/n5634 ;
  wire \u2_Display/n5635 ;
  wire \u2_Display/n5636 ;
  wire \u2_Display/n5637 ;
  wire \u2_Display/n5638 ;
  wire \u2_Display/n5639 ;
  wire \u2_Display/n564 ;
  wire \u2_Display/n5640 ;
  wire \u2_Display/n5641 ;
  wire \u2_Display/n5642 ;
  wire \u2_Display/n5643 ;
  wire \u2_Display/n5644 ;
  wire \u2_Display/n5647 ;
  wire \u2_Display/n5648 ;
  wire \u2_Display/n5649 ;
  wire \u2_Display/n565 ;
  wire \u2_Display/n5650 ;
  wire \u2_Display/n5651 ;
  wire \u2_Display/n5652 ;
  wire \u2_Display/n5653 ;
  wire \u2_Display/n5654 ;
  wire \u2_Display/n5655 ;
  wire \u2_Display/n5656 ;
  wire \u2_Display/n5657 ;
  wire \u2_Display/n5658 ;
  wire \u2_Display/n5659 ;
  wire \u2_Display/n566 ;
  wire \u2_Display/n5660 ;
  wire \u2_Display/n5661 ;
  wire \u2_Display/n5662 ;
  wire \u2_Display/n5663 ;
  wire \u2_Display/n5664 ;
  wire \u2_Display/n5665 ;
  wire \u2_Display/n5666 ;
  wire \u2_Display/n5667 ;
  wire \u2_Display/n5668 ;
  wire \u2_Display/n5669 ;
  wire \u2_Display/n567 ;
  wire \u2_Display/n5670 ;
  wire \u2_Display/n5671 ;
  wire \u2_Display/n5672 ;
  wire \u2_Display/n5673 ;
  wire \u2_Display/n5674 ;
  wire \u2_Display/n5675 ;
  wire \u2_Display/n5676 ;
  wire \u2_Display/n5677 ;
  wire \u2_Display/n5678 ;
  wire \u2_Display/n5679 ;
  wire \u2_Display/n568 ;
  wire \u2_Display/n569 ;
  wire \u2_Display/n570 ;
  wire \u2_Display/n571 ;
  wire \u2_Display/n572 ;
  wire \u2_Display/n573 ;
  wire \u2_Display/n574 ;
  wire \u2_Display/n575 ;
  wire \u2_Display/n576 ;
  wire \u2_Display/n577 ;
  wire \u2_Display/n578 ;
  wire \u2_Display/n579 ;
  wire \u2_Display/n580 ;
  wire \u2_Display/n581 ;
  wire \u2_Display/n582 ;
  wire \u2_Display/n583 ;
  wire \u2_Display/n584 ;
  wire \u2_Display/n585 ;
  wire \u2_Display/n586 ;
  wire \u2_Display/n587 ;
  wire \u2_Display/n588 ;
  wire \u2_Display/n589 ;
  wire \u2_Display/n590 ;
  wire \u2_Display/n591 ;
  wire \u2_Display/n592 ;
  wire \u2_Display/n595 ;
  wire \u2_Display/n596 ;
  wire \u2_Display/n597 ;
  wire \u2_Display/n598 ;
  wire \u2_Display/n599 ;
  wire \u2_Display/n600 ;
  wire \u2_Display/n601 ;
  wire \u2_Display/n602 ;
  wire \u2_Display/n603 ;
  wire \u2_Display/n604 ;
  wire \u2_Display/n605 ;
  wire \u2_Display/n606 ;
  wire \u2_Display/n607 ;
  wire \u2_Display/n6070 ;
  wire \u2_Display/n6071 ;
  wire \u2_Display/n6072 ;
  wire \u2_Display/n6073 ;
  wire \u2_Display/n6074 ;
  wire \u2_Display/n6075 ;
  wire \u2_Display/n6076 ;
  wire \u2_Display/n6077 ;
  wire \u2_Display/n6078 ;
  wire \u2_Display/n6079 ;
  wire \u2_Display/n608 ;
  wire \u2_Display/n6080 ;
  wire \u2_Display/n6081 ;
  wire \u2_Display/n6082 ;
  wire \u2_Display/n6083 ;
  wire \u2_Display/n6084 ;
  wire \u2_Display/n6085 ;
  wire \u2_Display/n6086 ;
  wire \u2_Display/n6087 ;
  wire \u2_Display/n6088 ;
  wire \u2_Display/n6089 ;
  wire \u2_Display/n609 ;
  wire \u2_Display/n6090 ;
  wire \u2_Display/n6091 ;
  wire \u2_Display/n6092 ;
  wire \u2_Display/n6093 ;
  wire \u2_Display/n6094 ;
  wire \u2_Display/n6095 ;
  wire \u2_Display/n6096 ;
  wire \u2_Display/n6097 ;
  wire \u2_Display/n6098 ;
  wire \u2_Display/n6099 ;
  wire \u2_Display/n610 ;
  wire \u2_Display/n6100 ;
  wire \u2_Display/n6101 ;
  wire \u2_Display/n6105 ;
  wire \u2_Display/n6106 ;
  wire \u2_Display/n6107 ;
  wire \u2_Display/n6108 ;
  wire \u2_Display/n6109 ;
  wire \u2_Display/n611 ;
  wire \u2_Display/n6110 ;
  wire \u2_Display/n6111 ;
  wire \u2_Display/n6112 ;
  wire \u2_Display/n6113 ;
  wire \u2_Display/n6114 ;
  wire \u2_Display/n6115 ;
  wire \u2_Display/n6116 ;
  wire \u2_Display/n6117 ;
  wire \u2_Display/n6118 ;
  wire \u2_Display/n6119 ;
  wire \u2_Display/n612 ;
  wire \u2_Display/n6120 ;
  wire \u2_Display/n6121 ;
  wire \u2_Display/n6122 ;
  wire \u2_Display/n6123 ;
  wire \u2_Display/n6124 ;
  wire \u2_Display/n6125 ;
  wire \u2_Display/n6126 ;
  wire \u2_Display/n6127 ;
  wire \u2_Display/n6128 ;
  wire \u2_Display/n6129 ;
  wire \u2_Display/n613 ;
  wire \u2_Display/n6130 ;
  wire \u2_Display/n6131 ;
  wire \u2_Display/n6132 ;
  wire \u2_Display/n6133 ;
  wire \u2_Display/n6134 ;
  wire \u2_Display/n6135 ;
  wire \u2_Display/n6136 ;
  wire \u2_Display/n614 ;
  wire \u2_Display/n6140 ;
  wire \u2_Display/n6141 ;
  wire \u2_Display/n6142 ;
  wire \u2_Display/n6143 ;
  wire \u2_Display/n6144 ;
  wire \u2_Display/n6145 ;
  wire \u2_Display/n6146 ;
  wire \u2_Display/n6147 ;
  wire \u2_Display/n6148 ;
  wire \u2_Display/n6149 ;
  wire \u2_Display/n615 ;
  wire \u2_Display/n6150 ;
  wire \u2_Display/n6151 ;
  wire \u2_Display/n6152 ;
  wire \u2_Display/n6153 ;
  wire \u2_Display/n6154 ;
  wire \u2_Display/n6155 ;
  wire \u2_Display/n6156 ;
  wire \u2_Display/n6157 ;
  wire \u2_Display/n6158 ;
  wire \u2_Display/n6159 ;
  wire \u2_Display/n616 ;
  wire \u2_Display/n6160 ;
  wire \u2_Display/n6161 ;
  wire \u2_Display/n6162 ;
  wire \u2_Display/n6163 ;
  wire \u2_Display/n6164 ;
  wire \u2_Display/n6165 ;
  wire \u2_Display/n6166 ;
  wire \u2_Display/n6167 ;
  wire \u2_Display/n6168 ;
  wire \u2_Display/n6169 ;
  wire \u2_Display/n617 ;
  wire \u2_Display/n6170 ;
  wire \u2_Display/n6171 ;
  wire \u2_Display/n6175 ;
  wire \u2_Display/n6176 ;
  wire \u2_Display/n6177 ;
  wire \u2_Display/n6178 ;
  wire \u2_Display/n6179 ;
  wire \u2_Display/n618 ;
  wire \u2_Display/n6180 ;
  wire \u2_Display/n6181 ;
  wire \u2_Display/n6182 ;
  wire \u2_Display/n6183 ;
  wire \u2_Display/n6184 ;
  wire \u2_Display/n6185 ;
  wire \u2_Display/n6186 ;
  wire \u2_Display/n6187 ;
  wire \u2_Display/n6188 ;
  wire \u2_Display/n6189 ;
  wire \u2_Display/n619 ;
  wire \u2_Display/n6190 ;
  wire \u2_Display/n6191 ;
  wire \u2_Display/n6192 ;
  wire \u2_Display/n6193 ;
  wire \u2_Display/n6194 ;
  wire \u2_Display/n6195 ;
  wire \u2_Display/n6196 ;
  wire \u2_Display/n6197 ;
  wire \u2_Display/n6198 ;
  wire \u2_Display/n6199 ;
  wire \u2_Display/n620 ;
  wire \u2_Display/n6200 ;
  wire \u2_Display/n6201 ;
  wire \u2_Display/n6202 ;
  wire \u2_Display/n6203 ;
  wire \u2_Display/n6204 ;
  wire \u2_Display/n6205 ;
  wire \u2_Display/n6206 ;
  wire \u2_Display/n621 ;
  wire \u2_Display/n6210 ;
  wire \u2_Display/n6211 ;
  wire \u2_Display/n6212 ;
  wire \u2_Display/n6213 ;
  wire \u2_Display/n6214 ;
  wire \u2_Display/n6215 ;
  wire \u2_Display/n6216 ;
  wire \u2_Display/n6217 ;
  wire \u2_Display/n6218 ;
  wire \u2_Display/n6219 ;
  wire \u2_Display/n622 ;
  wire \u2_Display/n6220 ;
  wire \u2_Display/n6221 ;
  wire \u2_Display/n6222 ;
  wire \u2_Display/n6223 ;
  wire \u2_Display/n6224 ;
  wire \u2_Display/n6225 ;
  wire \u2_Display/n6226 ;
  wire \u2_Display/n6227 ;
  wire \u2_Display/n6228 ;
  wire \u2_Display/n6229 ;
  wire \u2_Display/n623 ;
  wire \u2_Display/n6230 ;
  wire \u2_Display/n6231 ;
  wire \u2_Display/n6232 ;
  wire \u2_Display/n6233 ;
  wire \u2_Display/n6234 ;
  wire \u2_Display/n6235 ;
  wire \u2_Display/n6236 ;
  wire \u2_Display/n6237 ;
  wire \u2_Display/n6238 ;
  wire \u2_Display/n6239 ;
  wire \u2_Display/n624 ;
  wire \u2_Display/n6240 ;
  wire \u2_Display/n6241 ;
  wire \u2_Display/n6245 ;
  wire \u2_Display/n6246 ;
  wire \u2_Display/n6247 ;
  wire \u2_Display/n6248 ;
  wire \u2_Display/n6249 ;
  wire \u2_Display/n625 ;
  wire \u2_Display/n6250 ;
  wire \u2_Display/n6251 ;
  wire \u2_Display/n6252 ;
  wire \u2_Display/n6253 ;
  wire \u2_Display/n6254 ;
  wire \u2_Display/n6255 ;
  wire \u2_Display/n6256 ;
  wire \u2_Display/n6257 ;
  wire \u2_Display/n6258 ;
  wire \u2_Display/n6259 ;
  wire \u2_Display/n626 ;
  wire \u2_Display/n6260 ;
  wire \u2_Display/n6261 ;
  wire \u2_Display/n6262 ;
  wire \u2_Display/n6263 ;
  wire \u2_Display/n6264 ;
  wire \u2_Display/n6265 ;
  wire \u2_Display/n6266 ;
  wire \u2_Display/n6267 ;
  wire \u2_Display/n6268 ;
  wire \u2_Display/n6269 ;
  wire \u2_Display/n627 ;
  wire \u2_Display/n6270 ;
  wire \u2_Display/n6271 ;
  wire \u2_Display/n6272 ;
  wire \u2_Display/n6273 ;
  wire \u2_Display/n6274 ;
  wire \u2_Display/n6275 ;
  wire \u2_Display/n6276 ;
  wire \u2_Display/n6280 ;
  wire \u2_Display/n6281 ;
  wire \u2_Display/n6282 ;
  wire \u2_Display/n6283 ;
  wire \u2_Display/n6284 ;
  wire \u2_Display/n6285 ;
  wire \u2_Display/n6286 ;
  wire \u2_Display/n6287 ;
  wire \u2_Display/n6288 ;
  wire \u2_Display/n6289 ;
  wire \u2_Display/n6290 ;
  wire \u2_Display/n6291 ;
  wire \u2_Display/n6292 ;
  wire \u2_Display/n6293 ;
  wire \u2_Display/n6294 ;
  wire \u2_Display/n6295 ;
  wire \u2_Display/n6296 ;
  wire \u2_Display/n6297 ;
  wire \u2_Display/n6298 ;
  wire \u2_Display/n6299 ;
  wire \u2_Display/n630 ;
  wire \u2_Display/n6300 ;
  wire \u2_Display/n6301 ;
  wire \u2_Display/n6302 ;
  wire \u2_Display/n6303 ;
  wire \u2_Display/n6304 ;
  wire \u2_Display/n6305 ;
  wire \u2_Display/n6306 ;
  wire \u2_Display/n6307 ;
  wire \u2_Display/n6308 ;
  wire \u2_Display/n6309 ;
  wire \u2_Display/n631 ;
  wire \u2_Display/n6310 ;
  wire \u2_Display/n6311 ;
  wire \u2_Display/n6315 ;
  wire \u2_Display/n6316 ;
  wire \u2_Display/n6317 ;
  wire \u2_Display/n6318 ;
  wire \u2_Display/n6319 ;
  wire \u2_Display/n632 ;
  wire \u2_Display/n6320 ;
  wire \u2_Display/n6321 ;
  wire \u2_Display/n6322 ;
  wire \u2_Display/n6323 ;
  wire \u2_Display/n6324 ;
  wire \u2_Display/n6325 ;
  wire \u2_Display/n6326 ;
  wire \u2_Display/n6327 ;
  wire \u2_Display/n6328 ;
  wire \u2_Display/n6329 ;
  wire \u2_Display/n633 ;
  wire \u2_Display/n6330 ;
  wire \u2_Display/n6331 ;
  wire \u2_Display/n6332 ;
  wire \u2_Display/n6333 ;
  wire \u2_Display/n6334 ;
  wire \u2_Display/n6335 ;
  wire \u2_Display/n6336 ;
  wire \u2_Display/n6337 ;
  wire \u2_Display/n6338 ;
  wire \u2_Display/n6339 ;
  wire \u2_Display/n634 ;
  wire \u2_Display/n6340 ;
  wire \u2_Display/n6341 ;
  wire \u2_Display/n6342 ;
  wire \u2_Display/n6343 ;
  wire \u2_Display/n6344 ;
  wire \u2_Display/n6345 ;
  wire \u2_Display/n6346 ;
  wire \u2_Display/n635 ;
  wire \u2_Display/n6350 ;
  wire \u2_Display/n6351 ;
  wire \u2_Display/n6352 ;
  wire \u2_Display/n6353 ;
  wire \u2_Display/n636 ;
  wire \u2_Display/n637 ;
  wire \u2_Display/n638 ;
  wire \u2_Display/n639 ;
  wire \u2_Display/n640 ;
  wire \u2_Display/n641 ;
  wire \u2_Display/n642 ;
  wire \u2_Display/n643 ;
  wire \u2_Display/n644 ;
  wire \u2_Display/n645 ;
  wire \u2_Display/n646 ;
  wire \u2_Display/n647 ;
  wire \u2_Display/n648 ;
  wire \u2_Display/n649 ;
  wire \u2_Display/n650 ;
  wire \u2_Display/n651 ;
  wire \u2_Display/n652 ;
  wire \u2_Display/n653 ;
  wire \u2_Display/n654 ;
  wire \u2_Display/n655 ;
  wire \u2_Display/n656 ;
  wire \u2_Display/n657 ;
  wire \u2_Display/n658 ;
  wire \u2_Display/n659 ;
  wire \u2_Display/n660 ;
  wire \u2_Display/n661 ;
  wire \u2_Display/n662 ;
  wire \u2_Display/n665 ;
  wire \u2_Display/n666 ;
  wire \u2_Display/n667 ;
  wire \u2_Display/n668 ;
  wire \u2_Display/n669 ;
  wire \u2_Display/n670 ;
  wire \u2_Display/n671 ;
  wire \u2_Display/n672 ;
  wire \u2_Display/n673 ;
  wire \u2_Display/n674 ;
  wire \u2_Display/n675 ;
  wire \u2_Display/n676 ;
  wire \u2_Display/n677 ;
  wire \u2_Display/n678 ;
  wire \u2_Display/n679 ;
  wire \u2_Display/n680 ;
  wire \u2_Display/n681 ;
  wire \u2_Display/n682 ;
  wire \u2_Display/n683 ;
  wire \u2_Display/n684 ;
  wire \u2_Display/n685 ;
  wire \u2_Display/n686 ;
  wire \u2_Display/n687 ;
  wire \u2_Display/n688 ;
  wire \u2_Display/n689 ;
  wire \u2_Display/n690 ;
  wire \u2_Display/n691 ;
  wire \u2_Display/n692 ;
  wire \u2_Display/n693 ;
  wire \u2_Display/n694 ;
  wire \u2_Display/n695 ;
  wire \u2_Display/n696 ;
  wire \u2_Display/n697 ;
  wire \u2_Display/n700 ;
  wire \u2_Display/n701 ;
  wire \u2_Display/n702 ;
  wire \u2_Display/n703 ;
  wire \u2_Display/n704 ;
  wire \u2_Display/n705 ;
  wire \u2_Display/n706 ;
  wire \u2_Display/n707 ;
  wire \u2_Display/n708 ;
  wire \u2_Display/n709 ;
  wire \u2_Display/n710 ;
  wire \u2_Display/n711 ;
  wire \u2_Display/n712 ;
  wire \u2_Display/n713 ;
  wire \u2_Display/n714 ;
  wire \u2_Display/n715 ;
  wire \u2_Display/n716 ;
  wire \u2_Display/n717 ;
  wire \u2_Display/n718 ;
  wire \u2_Display/n719 ;
  wire \u2_Display/n720 ;
  wire \u2_Display/n721 ;
  wire \u2_Display/n722 ;
  wire \u2_Display/n723 ;
  wire \u2_Display/n724 ;
  wire \u2_Display/n725 ;
  wire \u2_Display/n726 ;
  wire \u2_Display/n727 ;
  wire \u2_Display/n728 ;
  wire \u2_Display/n729 ;
  wire \u2_Display/n730 ;
  wire \u2_Display/n731 ;
  wire \u2_Display/n732 ;
  wire \u2_Display/n735 ;
  wire \u2_Display/n736 ;
  wire \u2_Display/n737 ;
  wire \u2_Display/n738 ;
  wire \u2_Display/n739 ;
  wire \u2_Display/n740 ;
  wire \u2_Display/n741 ;
  wire \u2_Display/n742 ;
  wire \u2_Display/n743 ;
  wire \u2_Display/n744 ;
  wire \u2_Display/n745 ;
  wire \u2_Display/n746 ;
  wire \u2_Display/n747 ;
  wire \u2_Display/n748 ;
  wire \u2_Display/n749 ;
  wire \u2_Display/n750 ;
  wire \u2_Display/n751 ;
  wire \u2_Display/n752 ;
  wire \u2_Display/n753 ;
  wire \u2_Display/n754 ;
  wire \u2_Display/n755 ;
  wire \u2_Display/n756 ;
  wire \u2_Display/n757 ;
  wire \u2_Display/n758 ;
  wire \u2_Display/n759 ;
  wire \u2_Display/n760 ;
  wire \u2_Display/n761 ;
  wire \u2_Display/n762 ;
  wire \u2_Display/n763 ;
  wire \u2_Display/n764 ;
  wire \u2_Display/n765 ;
  wire \u2_Display/n766 ;
  wire \u2_Display/n767 ;
  wire \u2_Display/n770 ;
  wire \u2_Display/n771 ;
  wire \u2_Display/n772 ;
  wire \u2_Display/n773 ;
  wire \u2_Display/n774 ;
  wire \u2_Display/n775 ;
  wire \u2_Display/n776 ;
  wire \u2_Display/n777 ;
  wire \u2_Display/n778 ;
  wire \u2_Display/n779 ;
  wire \u2_Display/n780 ;
  wire \u2_Display/n781 ;
  wire \u2_Display/n782 ;
  wire \u2_Display/n783 ;
  wire \u2_Display/n784 ;
  wire \u2_Display/n785 ;
  wire \u2_Display/n786 ;
  wire \u2_Display/n787 ;
  wire \u2_Display/n788 ;
  wire \u2_Display/n789 ;
  wire \u2_Display/n790 ;
  wire \u2_Display/n791 ;
  wire \u2_Display/n792 ;
  wire \u2_Display/n793 ;
  wire \u2_Display/n794 ;
  wire \u2_Display/n795 ;
  wire \u2_Display/n796 ;
  wire \u2_Display/n797 ;
  wire \u2_Display/n798 ;
  wire \u2_Display/n799 ;
  wire \u2_Display/n800 ;
  wire \u2_Display/n801 ;
  wire \u2_Display/n802 ;
  wire \u2_Display/n805 ;
  wire \u2_Display/n806 ;
  wire \u2_Display/n807 ;
  wire \u2_Display/n808 ;
  wire \u2_Display/n809 ;
  wire \u2_Display/n810 ;
  wire \u2_Display/n811 ;
  wire \u2_Display/n812 ;
  wire \u2_Display/n813 ;
  wire \u2_Display/n814 ;
  wire \u2_Display/n815 ;
  wire \u2_Display/n816 ;
  wire \u2_Display/n817 ;
  wire \u2_Display/n818 ;
  wire \u2_Display/n819 ;
  wire \u2_Display/n820 ;
  wire \u2_Display/n821 ;
  wire \u2_Display/n822 ;
  wire \u2_Display/n823 ;
  wire \u2_Display/n824 ;
  wire \u2_Display/n825 ;
  wire \u2_Display/n826 ;
  wire \u2_Display/n827 ;
  wire \u2_Display/n828 ;
  wire \u2_Display/n829 ;
  wire \u2_Display/n830 ;
  wire \u2_Display/n831 ;
  wire \u2_Display/n832 ;
  wire \u2_Display/n833 ;
  wire \u2_Display/n834 ;
  wire \u2_Display/n835 ;
  wire \u2_Display/n836 ;
  wire \u2_Display/n837 ;
  wire \u2_Display/n840 ;
  wire \u2_Display/n841 ;
  wire \u2_Display/n842 ;
  wire \u2_Display/n843 ;
  wire \u2_Display/n844 ;
  wire \u2_Display/n845 ;
  wire \u2_Display/n846 ;
  wire \u2_Display/n847 ;
  wire \u2_Display/n848 ;
  wire \u2_Display/n849 ;
  wire \u2_Display/n850 ;
  wire \u2_Display/n851 ;
  wire \u2_Display/n852 ;
  wire \u2_Display/n853 ;
  wire \u2_Display/n854 ;
  wire \u2_Display/n855 ;
  wire \u2_Display/n856 ;
  wire \u2_Display/n857 ;
  wire \u2_Display/n858 ;
  wire \u2_Display/n859 ;
  wire \u2_Display/n860 ;
  wire \u2_Display/n861 ;
  wire \u2_Display/n862 ;
  wire \u2_Display/n863 ;
  wire \u2_Display/n864 ;
  wire \u2_Display/n865 ;
  wire \u2_Display/n866 ;
  wire \u2_Display/n867 ;
  wire \u2_Display/n868 ;
  wire \u2_Display/n869 ;
  wire \u2_Display/n870 ;
  wire \u2_Display/n871 ;
  wire \u2_Display/n872 ;
  wire \u2_Display/n875 ;
  wire \u2_Display/n876 ;
  wire \u2_Display/n877 ;
  wire \u2_Display/n878 ;
  wire \u2_Display/n879 ;
  wire \u2_Display/n880 ;
  wire \u2_Display/n881 ;
  wire \u2_Display/n882 ;
  wire \u2_Display/n883 ;
  wire \u2_Display/n884 ;
  wire \u2_Display/n885 ;
  wire \u2_Display/n886 ;
  wire \u2_Display/n887 ;
  wire \u2_Display/n888 ;
  wire \u2_Display/n889 ;
  wire \u2_Display/n890 ;
  wire \u2_Display/n891 ;
  wire \u2_Display/n892 ;
  wire \u2_Display/n893 ;
  wire \u2_Display/n894 ;
  wire \u2_Display/n895 ;
  wire \u2_Display/n896 ;
  wire \u2_Display/n897 ;
  wire \u2_Display/n898 ;
  wire \u2_Display/n899 ;
  wire \u2_Display/n900 ;
  wire \u2_Display/n901 ;
  wire \u2_Display/n902 ;
  wire \u2_Display/n903 ;
  wire \u2_Display/n904 ;
  wire \u2_Display/n905 ;
  wire \u2_Display/n906 ;
  wire \u2_Display/n907 ;
  wire \u2_Display/n910 ;
  wire \u2_Display/n911 ;
  wire \u2_Display/n912 ;
  wire \u2_Display/n913 ;
  wire \u2_Display/n914 ;
  wire \u2_Display/n915 ;
  wire \u2_Display/n916 ;
  wire \u2_Display/n917 ;
  wire \u2_Display/n918 ;
  wire \u2_Display/n919 ;
  wire \u2_Display/n920 ;
  wire \u2_Display/n921 ;
  wire \u2_Display/n922 ;
  wire \u2_Display/n923 ;
  wire \u2_Display/n924 ;
  wire \u2_Display/n925 ;
  wire \u2_Display/n926 ;
  wire \u2_Display/n927 ;
  wire \u2_Display/n928 ;
  wire \u2_Display/n929 ;
  wire \u2_Display/n930 ;
  wire \u2_Display/n931 ;
  wire \u2_Display/n932 ;
  wire \u2_Display/n933 ;
  wire \u2_Display/n934 ;
  wire \u2_Display/n935 ;
  wire \u2_Display/n936 ;
  wire \u2_Display/n937 ;
  wire \u2_Display/n938 ;
  wire \u2_Display/n939 ;
  wire \u2_Display/n940 ;
  wire \u2_Display/n941 ;
  wire \u2_Display/n942 ;
  wire \u2_Display/n945 ;
  wire \u2_Display/n946 ;
  wire \u2_Display/n947 ;
  wire \u2_Display/n948 ;
  wire \u2_Display/n949 ;
  wire \u2_Display/n95 ;
  wire \u2_Display/n950 ;
  wire \u2_Display/n951 ;
  wire \u2_Display/n952 ;
  wire \u2_Display/n953 ;
  wire \u2_Display/n954 ;
  wire \u2_Display/n955 ;
  wire \u2_Display/n956 ;
  wire \u2_Display/n957 ;
  wire \u2_Display/n958 ;
  wire \u2_Display/n959 ;
  wire \u2_Display/n960 ;
  wire \u2_Display/n961 ;
  wire \u2_Display/n962 ;
  wire \u2_Display/n963 ;
  wire \u2_Display/n964 ;
  wire \u2_Display/n965 ;
  wire \u2_Display/n966 ;
  wire \u2_Display/n967 ;
  wire \u2_Display/n968 ;
  wire \u2_Display/n969 ;
  wire \u2_Display/n97 ;
  wire \u2_Display/n970 ;
  wire \u2_Display/n971 ;
  wire \u2_Display/n972 ;
  wire \u2_Display/n973 ;
  wire \u2_Display/n974 ;
  wire \u2_Display/n975 ;
  wire \u2_Display/n976 ;
  wire \u2_Display/n977 ;
  wire \u2_Display/n980 ;
  wire \u2_Display/n981 ;
  wire \u2_Display/n982 ;
  wire \u2_Display/n983 ;
  wire \u2_Display/n984 ;
  wire \u2_Display/n985 ;
  wire \u2_Display/n986 ;
  wire \u2_Display/n987 ;
  wire \u2_Display/n988 ;
  wire \u2_Display/n989 ;
  wire \u2_Display/n990 ;
  wire \u2_Display/n991 ;
  wire \u2_Display/n992 ;
  wire \u2_Display/n993 ;
  wire \u2_Display/n994 ;
  wire \u2_Display/n995 ;
  wire \u2_Display/n996 ;
  wire \u2_Display/n997 ;
  wire \u2_Display/n998 ;
  wire \u2_Display/n999 ;
  wire \u2_Display/sub0_2/c0 ;
  wire \u2_Display/sub0_2/c1 ;
  wire \u2_Display/sub0_2/c10 ;
  wire \u2_Display/sub0_2/c11 ;
  wire \u2_Display/sub0_2/c2 ;
  wire \u2_Display/sub0_2/c3 ;
  wire \u2_Display/sub0_2/c4 ;
  wire \u2_Display/sub0_2/c5 ;
  wire \u2_Display/sub0_2/c6 ;
  wire \u2_Display/sub0_2/c7 ;
  wire \u2_Display/sub0_2/c8 ;
  wire \u2_Display/sub0_2/c9 ;
  wire \u2_Display/sub1_2/c0 ;
  wire \u2_Display/sub1_2/c1 ;
  wire \u2_Display/sub1_2/c10 ;
  wire \u2_Display/sub1_2/c2 ;
  wire \u2_Display/sub1_2/c3 ;
  wire \u2_Display/sub1_2/c4 ;
  wire \u2_Display/sub1_2/c5 ;
  wire \u2_Display/sub1_2/c6 ;
  wire \u2_Display/sub1_2/c7 ;
  wire \u2_Display/sub1_2/c8 ;
  wire \u2_Display/sub1_2/c9 ;
  wire \u2_Display/sub2_2/c0 ;
  wire \u2_Display/sub2_2/c1 ;
  wire \u2_Display/sub2_2/c10 ;
  wire \u2_Display/sub2_2/c2 ;
  wire \u2_Display/sub2_2/c3 ;
  wire \u2_Display/sub2_2/c4 ;
  wire \u2_Display/sub2_2/c5 ;
  wire \u2_Display/sub2_2/c6 ;
  wire \u2_Display/sub2_2/c7 ;
  wire \u2_Display/sub2_2/c8 ;
  wire \u2_Display/sub2_2/c9 ;
  wire \u2_Display/sub3_2/c0 ;
  wire \u2_Display/sub3_2/c1 ;
  wire \u2_Display/sub3_2/c10 ;
  wire \u2_Display/sub3_2/c11 ;
  wire \u2_Display/sub3_2/c2 ;
  wire \u2_Display/sub3_2/c3 ;
  wire \u2_Display/sub3_2/c4 ;
  wire \u2_Display/sub3_2/c5 ;
  wire \u2_Display/sub3_2/c6 ;
  wire \u2_Display/sub3_2/c7 ;
  wire \u2_Display/sub3_2/c8 ;
  wire \u2_Display/sub3_2/c9 ;
  wire vga_clk_pad;  // source/rtl/VGA_Demo.v(9)
  wire vga_de_pad;  // source/rtl/VGA_Demo.v(13)
  wire vga_hs_pad;  // source/rtl/VGA_Demo.v(10)
  wire vga_vs_pad;  // source/rtl/VGA_Demo.v(11)

  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1000 (
    .a(\u2_Display/n3925 ),
    .b(\u2_Display/n3928 [0]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3960 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1001 (
    .a(\u2_Display/n3924 ),
    .b(\u2_Display/n3928 [1]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3959 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1002 (
    .a(\u2_Display/n3923 ),
    .b(\u2_Display/n3928 [2]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3958 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1003 (
    .a(\u2_Display/n3922 ),
    .b(\u2_Display/n3928 [3]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3957 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1004 (
    .a(\u2_Display/n3921 ),
    .b(\u2_Display/n3928 [4]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3956 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1005 (
    .a(\u2_Display/n3920 ),
    .b(\u2_Display/n3928 [5]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3955 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1006 (
    .a(\u2_Display/n3919 ),
    .b(\u2_Display/n3928 [6]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3954 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1007 (
    .a(\u2_Display/n3918 ),
    .b(\u2_Display/n3928 [7]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3953 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1008 (
    .a(\u2_Display/n3917 ),
    .b(\u2_Display/n3928 [8]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3952 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1009 (
    .a(\u2_Display/n3916 ),
    .b(\u2_Display/n3928 [9]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3951 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1010 (
    .a(\u2_Display/n3915 ),
    .b(\u2_Display/n3928 [10]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3950 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1011 (
    .a(\u2_Display/n3914 ),
    .b(\u2_Display/n3928 [11]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3949 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1012 (
    .a(\u2_Display/n3913 ),
    .b(\u2_Display/n3928 [12]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3948 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1013 (
    .a(\u2_Display/n3912 ),
    .b(\u2_Display/n3928 [13]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3947 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1014 (
    .a(\u2_Display/n3911 ),
    .b(\u2_Display/n3928 [14]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3946 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1015 (
    .a(\u2_Display/n3910 ),
    .b(\u2_Display/n3928 [15]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3945 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1016 (
    .a(\u2_Display/n3909 ),
    .b(\u2_Display/n3928 [16]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3944 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1017 (
    .a(\u2_Display/n3908 ),
    .b(\u2_Display/n3928 [17]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3943 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1018 (
    .a(\u2_Display/n3907 ),
    .b(\u2_Display/n3928 [18]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3942 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1019 (
    .a(\u2_Display/n3906 ),
    .b(\u2_Display/n3928 [19]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3941 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1020 (
    .a(\u2_Display/n3905 ),
    .b(\u2_Display/n3928 [20]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3940 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1021 (
    .a(\u2_Display/n3904 ),
    .b(\u2_Display/n3928 [21]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3939 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1022 (
    .a(\u2_Display/n3903 ),
    .b(\u2_Display/n3928 [22]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3938 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1023 (
    .a(\u2_Display/n3902 ),
    .b(\u2_Display/n3928 [23]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3937 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1024 (
    .a(\u2_Display/n3901 ),
    .b(\u2_Display/n3928 [24]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3936 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1025 (
    .a(\u2_Display/n3900 ),
    .b(\u2_Display/n3928 [25]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3935 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1026 (
    .a(\u2_Display/n3899 ),
    .b(\u2_Display/n3928 [26]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3934 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1027 (
    .a(\u2_Display/n3898 ),
    .b(\u2_Display/n3928 [27]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3933 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1028 (
    .a(\u2_Display/n3897 ),
    .b(\u2_Display/n3928 [28]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3932 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1029 (
    .a(\u2_Display/n3896 ),
    .b(\u2_Display/n3928 [29]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3931 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1030 (
    .a(\u2_Display/n3895 ),
    .b(\u2_Display/n3928 [30]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3930 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1031 (
    .a(\u2_Display/n3894 ),
    .b(\u2_Display/n3928 [31]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3929 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1032 (
    .a(\u2_Display/n6206 ),
    .b(\u2_Display/n5051 [0]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6241 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1033 (
    .a(\u2_Display/n6205 ),
    .b(\u2_Display/n5051 [1]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6240 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1034 (
    .a(\u2_Display/n6204 ),
    .b(\u2_Display/n5051 [2]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6239 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1035 (
    .a(\u2_Display/n6203 ),
    .b(\u2_Display/n5051 [3]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6238 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1036 (
    .a(\u2_Display/n6202 ),
    .b(\u2_Display/n5051 [4]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6237 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1037 (
    .a(\u2_Display/n6201 ),
    .b(\u2_Display/n5051 [5]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6236 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1038 (
    .a(\u2_Display/n6200 ),
    .b(\u2_Display/n5051 [6]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6235 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1039 (
    .a(\u2_Display/n6199 ),
    .b(\u2_Display/n5051 [7]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6234 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1040 (
    .a(\u2_Display/n6198 ),
    .b(\u2_Display/n5051 [8]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6233 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1041 (
    .a(\u2_Display/n6197 ),
    .b(\u2_Display/n5051 [9]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6232 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1042 (
    .a(\u2_Display/n6196 ),
    .b(\u2_Display/n5051 [10]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6231 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1043 (
    .a(\u2_Display/n6195 ),
    .b(\u2_Display/n5051 [11]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6230 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1044 (
    .a(\u2_Display/n6194 ),
    .b(\u2_Display/n5051 [12]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6229 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1045 (
    .a(\u2_Display/n6193 ),
    .b(\u2_Display/n5051 [13]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6228 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1046 (
    .a(\u2_Display/n6192 ),
    .b(\u2_Display/n5051 [14]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6227 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1047 (
    .a(\u2_Display/n6191 ),
    .b(\u2_Display/n5051 [15]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6226 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1048 (
    .a(\u2_Display/n6190 ),
    .b(\u2_Display/n5051 [16]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6225 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1049 (
    .a(\u2_Display/n6189 ),
    .b(\u2_Display/n5051 [17]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6224 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1050 (
    .a(\u2_Display/n6188 ),
    .b(\u2_Display/n5051 [18]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6223 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1051 (
    .a(\u2_Display/n6187 ),
    .b(\u2_Display/n5051 [19]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6222 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1052 (
    .a(\u2_Display/n6186 ),
    .b(\u2_Display/n5051 [20]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6221 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1053 (
    .a(\u2_Display/n6185 ),
    .b(\u2_Display/n5051 [21]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6220 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1054 (
    .a(\u2_Display/n6184 ),
    .b(\u2_Display/n5051 [22]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6219 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1055 (
    .a(\u2_Display/n6183 ),
    .b(\u2_Display/n5051 [23]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6218 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1056 (
    .a(\u2_Display/n6182 ),
    .b(\u2_Display/n5051 [24]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6217 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1057 (
    .a(\u2_Display/n6181 ),
    .b(\u2_Display/n5051 [25]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6216 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1058 (
    .a(\u2_Display/n6180 ),
    .b(\u2_Display/n5051 [26]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6215 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1059 (
    .a(\u2_Display/n6179 ),
    .b(\u2_Display/n5051 [27]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6214 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1060 (
    .a(\u2_Display/n6178 ),
    .b(\u2_Display/n5051 [28]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6213 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1061 (
    .a(\u2_Display/n6177 ),
    .b(\u2_Display/n5051 [29]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6212 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1062 (
    .a(\u2_Display/n6176 ),
    .b(\u2_Display/n5051 [30]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6211 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1063 (
    .a(\u2_Display/n6175 ),
    .b(\u2_Display/n5051 [31]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6210 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1064 (
    .a(\u2_Display/n556 ),
    .b(\u2_Display/n559 [0]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n591 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1065 (
    .a(\u2_Display/n555 ),
    .b(\u2_Display/n559 [1]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n590 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1066 (
    .a(\u2_Display/n554 ),
    .b(\u2_Display/n559 [2]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n589 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1067 (
    .a(\u2_Display/n553 ),
    .b(\u2_Display/n559 [3]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n588 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1068 (
    .a(\u2_Display/n552 ),
    .b(\u2_Display/n559 [4]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n587 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1069 (
    .a(\u2_Display/n551 ),
    .b(\u2_Display/n559 [5]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n586 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1070 (
    .a(\u2_Display/n550 ),
    .b(\u2_Display/n559 [6]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n585 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1071 (
    .a(\u2_Display/n549 ),
    .b(\u2_Display/n559 [7]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n584 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1072 (
    .a(\u2_Display/n548 ),
    .b(\u2_Display/n559 [8]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n583 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1073 (
    .a(\u2_Display/n547 ),
    .b(\u2_Display/n559 [9]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n582 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1074 (
    .a(\u2_Display/n546 ),
    .b(\u2_Display/n559 [10]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n581 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1075 (
    .a(\u2_Display/n545 ),
    .b(\u2_Display/n559 [11]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n580 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1076 (
    .a(\u2_Display/n544 ),
    .b(\u2_Display/n559 [12]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n579 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1077 (
    .a(\u2_Display/n543 ),
    .b(\u2_Display/n559 [13]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n578 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1078 (
    .a(\u2_Display/n542 ),
    .b(\u2_Display/n559 [14]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n577 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1079 (
    .a(\u2_Display/n541 ),
    .b(\u2_Display/n559 [15]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n576 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1080 (
    .a(\u2_Display/n540 ),
    .b(\u2_Display/n559 [16]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n575 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1081 (
    .a(\u2_Display/n539 ),
    .b(\u2_Display/n559 [17]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n574 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1082 (
    .a(\u2_Display/n538 ),
    .b(\u2_Display/n559 [18]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n573 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1083 (
    .a(\u2_Display/n537 ),
    .b(\u2_Display/n559 [19]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n572 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1084 (
    .a(\u2_Display/n536 ),
    .b(\u2_Display/n559 [20]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n571 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1085 (
    .a(\u2_Display/n535 ),
    .b(\u2_Display/n559 [21]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n570 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1086 (
    .a(\u2_Display/n534 ),
    .b(\u2_Display/n559 [22]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n569 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1087 (
    .a(\u2_Display/n533 ),
    .b(\u2_Display/n559 [23]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n568 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1088 (
    .a(\u2_Display/n532 ),
    .b(\u2_Display/n559 [24]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n567 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1089 (
    .a(\u2_Display/n531 ),
    .b(\u2_Display/n559 [25]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n566 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1090 (
    .a(\u2_Display/n530 ),
    .b(\u2_Display/n559 [26]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n565 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1091 (
    .a(\u2_Display/n529 ),
    .b(\u2_Display/n559 [27]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n564 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1092 (
    .a(\u2_Display/n528 ),
    .b(\u2_Display/n559 [28]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n563 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1093 (
    .a(\u2_Display/n527 ),
    .b(\u2_Display/n559 [29]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n562 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1094 (
    .a(\u2_Display/n526 ),
    .b(\u2_Display/n559 [30]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n561 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1095 (
    .a(\u2_Display/n525 ),
    .b(\u2_Display/n559 [31]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n560 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1096 (
    .a(\u2_Display/n1679 ),
    .b(\u2_Display/n1682 [0]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1714 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1097 (
    .a(\u2_Display/n1678 ),
    .b(\u2_Display/n1682 [1]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1713 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1098 (
    .a(\u2_Display/n1677 ),
    .b(\u2_Display/n1682 [2]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1712 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1099 (
    .a(\u2_Display/n1676 ),
    .b(\u2_Display/n1682 [3]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1711 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1100 (
    .a(\u2_Display/n1675 ),
    .b(\u2_Display/n1682 [4]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1710 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1101 (
    .a(\u2_Display/n1674 ),
    .b(\u2_Display/n1682 [5]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1709 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1102 (
    .a(\u2_Display/n1673 ),
    .b(\u2_Display/n1682 [6]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1708 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1103 (
    .a(\u2_Display/n1672 ),
    .b(\u2_Display/n1682 [7]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1707 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1104 (
    .a(\u2_Display/n1671 ),
    .b(\u2_Display/n1682 [8]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1706 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1105 (
    .a(\u2_Display/n1670 ),
    .b(\u2_Display/n1682 [9]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1705 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1106 (
    .a(\u2_Display/n1669 ),
    .b(\u2_Display/n1682 [10]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1704 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1107 (
    .a(\u2_Display/n1668 ),
    .b(\u2_Display/n1682 [11]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1703 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1108 (
    .a(\u2_Display/n1667 ),
    .b(\u2_Display/n1682 [12]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1702 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1109 (
    .a(\u2_Display/n1666 ),
    .b(\u2_Display/n1682 [13]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1701 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1110 (
    .a(\u2_Display/n1665 ),
    .b(\u2_Display/n1682 [14]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1700 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1111 (
    .a(\u2_Display/n1664 ),
    .b(\u2_Display/n1682 [15]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1699 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1112 (
    .a(\u2_Display/n1663 ),
    .b(\u2_Display/n1682 [16]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1698 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1113 (
    .a(\u2_Display/n1662 ),
    .b(\u2_Display/n1682 [17]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1697 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1114 (
    .a(\u2_Display/n1661 ),
    .b(\u2_Display/n1682 [18]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1696 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1115 (
    .a(\u2_Display/n1660 ),
    .b(\u2_Display/n1682 [19]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1695 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1116 (
    .a(\u2_Display/n1659 ),
    .b(\u2_Display/n1682 [20]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1694 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1117 (
    .a(\u2_Display/n1658 ),
    .b(\u2_Display/n1682 [21]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1693 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1118 (
    .a(\u2_Display/n1657 ),
    .b(\u2_Display/n1682 [22]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1692 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1119 (
    .a(\u2_Display/n1656 ),
    .b(\u2_Display/n1682 [23]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1691 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1120 (
    .a(\u2_Display/n1655 ),
    .b(\u2_Display/n1682 [24]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1690 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1121 (
    .a(\u2_Display/n1654 ),
    .b(\u2_Display/n1682 [25]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1689 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1122 (
    .a(\u2_Display/n1653 ),
    .b(\u2_Display/n1682 [26]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1688 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1123 (
    .a(\u2_Display/n1652 ),
    .b(\u2_Display/n1682 [27]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1687 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1124 (
    .a(\u2_Display/n1651 ),
    .b(\u2_Display/n1682 [28]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1686 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1125 (
    .a(\u2_Display/n1650 ),
    .b(\u2_Display/n1682 [29]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1685 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1126 (
    .a(\u2_Display/n1649 ),
    .b(\u2_Display/n1682 [30]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1684 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1127 (
    .a(\u2_Display/n1648 ),
    .b(\u2_Display/n1682 [31]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1683 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1128 (
    .a(\u2_Display/n2802 ),
    .b(\u2_Display/n2805 [0]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2837 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1129 (
    .a(\u2_Display/n2801 ),
    .b(\u2_Display/n2805 [1]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2836 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1130 (
    .a(\u2_Display/n2800 ),
    .b(\u2_Display/n2805 [2]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2835 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1131 (
    .a(\u2_Display/n2799 ),
    .b(\u2_Display/n2805 [3]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2834 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1132 (
    .a(\u2_Display/n2798 ),
    .b(\u2_Display/n2805 [4]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2833 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1133 (
    .a(\u2_Display/n2797 ),
    .b(\u2_Display/n2805 [5]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2832 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1134 (
    .a(\u2_Display/n2796 ),
    .b(\u2_Display/n2805 [6]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2831 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1135 (
    .a(\u2_Display/n2795 ),
    .b(\u2_Display/n2805 [7]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2830 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1136 (
    .a(\u2_Display/n2794 ),
    .b(\u2_Display/n2805 [8]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2829 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1137 (
    .a(\u2_Display/n2793 ),
    .b(\u2_Display/n2805 [9]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2828 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1138 (
    .a(\u2_Display/n2792 ),
    .b(\u2_Display/n2805 [10]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2827 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1139 (
    .a(\u2_Display/n2791 ),
    .b(\u2_Display/n2805 [11]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2826 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1140 (
    .a(\u2_Display/n2790 ),
    .b(\u2_Display/n2805 [12]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2825 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1141 (
    .a(\u2_Display/n2789 ),
    .b(\u2_Display/n2805 [13]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2824 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1142 (
    .a(\u2_Display/n2788 ),
    .b(\u2_Display/n2805 [14]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2823 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1143 (
    .a(\u2_Display/n2787 ),
    .b(\u2_Display/n2805 [15]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2822 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1144 (
    .a(\u2_Display/n2786 ),
    .b(\u2_Display/n2805 [16]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2821 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1145 (
    .a(\u2_Display/n2785 ),
    .b(\u2_Display/n2805 [17]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2820 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1146 (
    .a(\u2_Display/n2784 ),
    .b(\u2_Display/n2805 [18]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2819 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1147 (
    .a(\u2_Display/n2783 ),
    .b(\u2_Display/n2805 [19]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2818 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1148 (
    .a(\u2_Display/n2782 ),
    .b(\u2_Display/n2805 [20]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2817 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1149 (
    .a(\u2_Display/n2781 ),
    .b(\u2_Display/n2805 [21]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2816 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1150 (
    .a(\u2_Display/n2780 ),
    .b(\u2_Display/n2805 [22]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2815 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1151 (
    .a(\u2_Display/n2779 ),
    .b(\u2_Display/n2805 [23]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2814 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1152 (
    .a(\u2_Display/n2778 ),
    .b(\u2_Display/n2805 [24]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2813 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1153 (
    .a(\u2_Display/n2777 ),
    .b(\u2_Display/n2805 [25]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2812 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1154 (
    .a(\u2_Display/n2776 ),
    .b(\u2_Display/n2805 [26]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2811 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1155 (
    .a(\u2_Display/n2775 ),
    .b(\u2_Display/n2805 [27]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2810 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1156 (
    .a(\u2_Display/n2774 ),
    .b(\u2_Display/n2805 [28]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2809 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1157 (
    .a(\u2_Display/n2773 ),
    .b(\u2_Display/n2805 [29]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2808 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1158 (
    .a(\u2_Display/n2772 ),
    .b(\u2_Display/n2805 [30]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2807 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1159 (
    .a(\u2_Display/n2771 ),
    .b(\u2_Display/n2805 [31]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2806 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1160 (
    .a(on_off_pad[3]),
    .b(on_off_pad[2]),
    .o(\u2_Display/mux11_b0_sel_is_0_o ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1161 (
    .a(on_off_pad[4]),
    .b(on_off_pad[3]),
    .o(\u2_Display/mux5_b0_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1162 (
    .a(\u2_Display/n141 ),
    .b(\u2_Display/n144 ),
    .c(\u2_Display/n136 ),
    .d(\u2_Display/n138 ),
    .o(\u2_Display/n145 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1163 (
    .a(on_off_pad[1]),
    .b(on_off_pad[0]),
    .o(\u2_Display/mux19_b0_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1164 (
    .a(\u2_Display/n44 ),
    .b(\u2_Display/n45 ),
    .c(\u2_Display/n48 ),
    .d(\u2_Display/n50 ),
    .o(\u2_Display/n51 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1165 (
    .a(\u2_Display/n95 ),
    .b(\u2_Display/n97 ),
    .c(\u2_Display/n100 ),
    .d(\u2_Display/n103 ),
    .o(\u2_Display/n104 ));
  AL_MAP_LUT5 #(
    .EQN("((A*~(~D*C))*~(B)*~(E)+(A*~(~D*C))*B*~(E)+~((A*~(~D*C)))*B*E+(A*~(~D*C))*B*E)"),
    .INIT(32'hccccaa0a))
    _al_u1166 (
    .a(\u2_Display/n145 ),
    .b(\u2_Display/n104 ),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(on_off_pad[1]),
    .o(\u2_Display/n236 [0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u1167 (
    .a(\u2_Display/n236 [0]),
    .b(\u2_Display/n51 ),
    .c(on_off_pad[0]),
    .o(\u2_Display/n240 [0]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1168 (
    .a(\u2_Display/mux11_b0_sel_is_0_o ),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(on_off_pad[4]),
    .o(_al_u1168_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1169 (
    .a(_al_u1168_o),
    .b(rst_n_pad),
    .o(\u2_Display/mux21_b0_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1170 (
    .a(\u1_Driver/vcnt [6]),
    .b(\u1_Driver/vcnt [7]),
    .c(\u1_Driver/vcnt [8]),
    .d(\u1_Driver/vcnt [9]),
    .o(_al_u1170_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    _al_u1171 (
    .a(_al_u1170_o),
    .b(\u1_Driver/vcnt [0]),
    .c(\u1_Driver/vcnt [10]),
    .d(\u1_Driver/vcnt [2]),
    .e(\u1_Driver/vcnt [4]),
    .o(_al_u1171_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*A)"),
    .INIT(32'h02000000))
    _al_u1172 (
    .a(_al_u1171_o),
    .b(\u1_Driver/vcnt [1]),
    .c(\u1_Driver/vcnt [11]),
    .d(\u1_Driver/vcnt [3]),
    .e(\u1_Driver/vcnt [5]),
    .o(\u1_Driver/n6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1173 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [9]),
    .o(\u1_Driver/n8 [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1174 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [8]),
    .o(\u1_Driver/n8 [8]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1175 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [7]),
    .o(\u1_Driver/n8 [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1176 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [6]),
    .o(\u1_Driver/n8 [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1177 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [5]),
    .o(\u1_Driver/n8 [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1178 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [4]),
    .o(\u1_Driver/n8 [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1179 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [3]),
    .o(\u1_Driver/n8 [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1180 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [2]),
    .o(\u1_Driver/n8 [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1181 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [11]),
    .o(\u1_Driver/n8 [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1182 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [10]),
    .o(\u1_Driver/n8 [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1183 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [1]),
    .o(\u1_Driver/n8 [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1184 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [0]),
    .o(\u1_Driver/n8 [0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1185 (
    .a(\u2_Display/n3960 ),
    .b(\u2_Display/n3963 [0]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3995 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1186 (
    .a(\u2_Display/n3959 ),
    .b(\u2_Display/n3963 [1]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3994 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1187 (
    .a(\u2_Display/n3958 ),
    .b(\u2_Display/n3963 [2]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3993 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1188 (
    .a(\u2_Display/n3957 ),
    .b(\u2_Display/n3963 [3]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3992 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1189 (
    .a(\u2_Display/n3956 ),
    .b(\u2_Display/n3963 [4]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3991 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1190 (
    .a(\u2_Display/n3955 ),
    .b(\u2_Display/n3963 [5]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3990 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1191 (
    .a(\u2_Display/n3954 ),
    .b(\u2_Display/n3963 [6]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3989 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1192 (
    .a(\u2_Display/n3953 ),
    .b(\u2_Display/n3963 [7]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3988 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1193 (
    .a(\u2_Display/n3952 ),
    .b(\u2_Display/n3963 [8]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3987 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1194 (
    .a(\u2_Display/n3951 ),
    .b(\u2_Display/n3963 [9]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3986 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1195 (
    .a(\u2_Display/n3950 ),
    .b(\u2_Display/n3963 [10]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3985 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1196 (
    .a(\u2_Display/n3949 ),
    .b(\u2_Display/n3963 [11]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3984 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1197 (
    .a(\u2_Display/n3948 ),
    .b(\u2_Display/n3963 [12]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3983 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1198 (
    .a(\u2_Display/n3947 ),
    .b(\u2_Display/n3963 [13]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3982 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1199 (
    .a(\u2_Display/n3946 ),
    .b(\u2_Display/n3963 [14]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3981 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1200 (
    .a(\u2_Display/n3945 ),
    .b(\u2_Display/n3963 [15]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3980 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1201 (
    .a(\u2_Display/n3944 ),
    .b(\u2_Display/n3963 [16]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3979 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1202 (
    .a(\u2_Display/n3943 ),
    .b(\u2_Display/n3963 [17]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3978 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1203 (
    .a(\u2_Display/n3942 ),
    .b(\u2_Display/n3963 [18]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3977 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1204 (
    .a(\u2_Display/n3941 ),
    .b(\u2_Display/n3963 [19]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3976 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1205 (
    .a(\u2_Display/n3940 ),
    .b(\u2_Display/n3963 [20]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3975 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1206 (
    .a(\u2_Display/n3939 ),
    .b(\u2_Display/n3963 [21]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3974 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1207 (
    .a(\u2_Display/n3938 ),
    .b(\u2_Display/n3963 [22]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3973 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1208 (
    .a(\u2_Display/n3937 ),
    .b(\u2_Display/n3963 [23]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3972 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1209 (
    .a(\u2_Display/n3936 ),
    .b(\u2_Display/n3963 [24]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3971 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1210 (
    .a(\u2_Display/n3935 ),
    .b(\u2_Display/n3963 [25]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3970 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1211 (
    .a(\u2_Display/n3934 ),
    .b(\u2_Display/n3963 [26]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3969 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1212 (
    .a(\u2_Display/n3933 ),
    .b(\u2_Display/n3963 [27]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3968 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1213 (
    .a(\u2_Display/n3932 ),
    .b(\u2_Display/n3963 [28]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3967 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1214 (
    .a(\u2_Display/n3931 ),
    .b(\u2_Display/n3963 [29]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3966 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1215 (
    .a(\u2_Display/n3930 ),
    .b(\u2_Display/n3963 [30]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3965 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1216 (
    .a(\u2_Display/n3929 ),
    .b(\u2_Display/n3963 [31]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3964 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1217 (
    .a(\u2_Display/n6241 ),
    .b(\u2_Display/n5086 [0]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6276 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1218 (
    .a(\u2_Display/n6240 ),
    .b(\u2_Display/n5086 [1]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6275 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1219 (
    .a(\u2_Display/n6239 ),
    .b(\u2_Display/n5086 [2]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6274 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1220 (
    .a(\u2_Display/n6238 ),
    .b(\u2_Display/n5086 [3]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6273 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1221 (
    .a(\u2_Display/n6237 ),
    .b(\u2_Display/n5086 [4]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6272 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1222 (
    .a(\u2_Display/n6236 ),
    .b(\u2_Display/n5086 [5]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6271 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1223 (
    .a(\u2_Display/n6235 ),
    .b(\u2_Display/n5086 [6]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6270 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1224 (
    .a(\u2_Display/n6234 ),
    .b(\u2_Display/n5086 [7]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6269 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1225 (
    .a(\u2_Display/n6233 ),
    .b(\u2_Display/n5086 [8]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6268 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1226 (
    .a(\u2_Display/n6232 ),
    .b(\u2_Display/n5086 [9]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6267 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1227 (
    .a(\u2_Display/n6231 ),
    .b(\u2_Display/n5086 [10]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6266 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1228 (
    .a(\u2_Display/n6230 ),
    .b(\u2_Display/n5086 [11]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6265 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1229 (
    .a(\u2_Display/n6229 ),
    .b(\u2_Display/n5086 [12]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6264 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1230 (
    .a(\u2_Display/n6228 ),
    .b(\u2_Display/n5086 [13]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6263 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1231 (
    .a(\u2_Display/n6227 ),
    .b(\u2_Display/n5086 [14]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6262 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1232 (
    .a(\u2_Display/n6226 ),
    .b(\u2_Display/n5086 [15]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6261 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1233 (
    .a(\u2_Display/n6225 ),
    .b(\u2_Display/n5086 [16]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6260 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1234 (
    .a(\u2_Display/n6224 ),
    .b(\u2_Display/n5086 [17]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6259 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1235 (
    .a(\u2_Display/n6223 ),
    .b(\u2_Display/n5086 [18]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6258 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1236 (
    .a(\u2_Display/n6222 ),
    .b(\u2_Display/n5086 [19]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6257 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1237 (
    .a(\u2_Display/n6221 ),
    .b(\u2_Display/n5086 [20]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6256 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1238 (
    .a(\u2_Display/n6220 ),
    .b(\u2_Display/n5086 [21]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6255 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1239 (
    .a(\u2_Display/n6219 ),
    .b(\u2_Display/n5086 [22]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6254 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1240 (
    .a(\u2_Display/n6218 ),
    .b(\u2_Display/n5086 [23]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6253 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1241 (
    .a(\u2_Display/n6217 ),
    .b(\u2_Display/n5086 [24]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6252 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1242 (
    .a(\u2_Display/n6216 ),
    .b(\u2_Display/n5086 [25]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6251 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1243 (
    .a(\u2_Display/n6215 ),
    .b(\u2_Display/n5086 [26]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6250 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1244 (
    .a(\u2_Display/n6214 ),
    .b(\u2_Display/n5086 [27]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6249 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1245 (
    .a(\u2_Display/n6213 ),
    .b(\u2_Display/n5086 [28]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6248 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1246 (
    .a(\u2_Display/n6212 ),
    .b(\u2_Display/n5086 [29]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6247 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1247 (
    .a(\u2_Display/n6211 ),
    .b(\u2_Display/n5086 [30]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6246 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1248 (
    .a(\u2_Display/n6210 ),
    .b(\u2_Display/n5086 [31]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6245 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1249 (
    .a(\u2_Display/n591 ),
    .b(\u2_Display/n594 [0]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n626 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1250 (
    .a(\u2_Display/n590 ),
    .b(\u2_Display/n594 [1]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n625 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1251 (
    .a(\u2_Display/n589 ),
    .b(\u2_Display/n594 [2]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n624 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1252 (
    .a(\u2_Display/n588 ),
    .b(\u2_Display/n594 [3]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n623 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1253 (
    .a(\u2_Display/n587 ),
    .b(\u2_Display/n594 [4]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n622 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1254 (
    .a(\u2_Display/n586 ),
    .b(\u2_Display/n594 [5]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n621 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1255 (
    .a(\u2_Display/n585 ),
    .b(\u2_Display/n594 [6]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n620 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1256 (
    .a(\u2_Display/n584 ),
    .b(\u2_Display/n594 [7]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n619 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1257 (
    .a(\u2_Display/n583 ),
    .b(\u2_Display/n594 [8]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n618 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1258 (
    .a(\u2_Display/n582 ),
    .b(\u2_Display/n594 [9]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n617 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1259 (
    .a(\u2_Display/n581 ),
    .b(\u2_Display/n594 [10]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n616 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1260 (
    .a(\u2_Display/n580 ),
    .b(\u2_Display/n594 [11]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n615 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1261 (
    .a(\u2_Display/n579 ),
    .b(\u2_Display/n594 [12]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n614 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1262 (
    .a(\u2_Display/n578 ),
    .b(\u2_Display/n594 [13]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n613 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1263 (
    .a(\u2_Display/n577 ),
    .b(\u2_Display/n594 [14]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n612 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1264 (
    .a(\u2_Display/n576 ),
    .b(\u2_Display/n594 [15]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n611 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1265 (
    .a(\u2_Display/n575 ),
    .b(\u2_Display/n594 [16]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n610 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1266 (
    .a(\u2_Display/n574 ),
    .b(\u2_Display/n594 [17]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n609 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1267 (
    .a(\u2_Display/n573 ),
    .b(\u2_Display/n594 [18]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n608 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1268 (
    .a(\u2_Display/n572 ),
    .b(\u2_Display/n594 [19]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n607 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1269 (
    .a(\u2_Display/n571 ),
    .b(\u2_Display/n594 [20]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n606 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1270 (
    .a(\u2_Display/n570 ),
    .b(\u2_Display/n594 [21]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n605 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1271 (
    .a(\u2_Display/n569 ),
    .b(\u2_Display/n594 [22]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n604 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1272 (
    .a(\u2_Display/n568 ),
    .b(\u2_Display/n594 [23]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n603 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1273 (
    .a(\u2_Display/n567 ),
    .b(\u2_Display/n594 [24]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n602 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1274 (
    .a(\u2_Display/n566 ),
    .b(\u2_Display/n594 [25]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n601 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1275 (
    .a(\u2_Display/n565 ),
    .b(\u2_Display/n594 [26]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n600 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1276 (
    .a(\u2_Display/n564 ),
    .b(\u2_Display/n594 [27]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n599 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1277 (
    .a(\u2_Display/n563 ),
    .b(\u2_Display/n594 [28]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n598 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1278 (
    .a(\u2_Display/n562 ),
    .b(\u2_Display/n594 [29]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n597 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1279 (
    .a(\u2_Display/n561 ),
    .b(\u2_Display/n594 [30]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n596 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1280 (
    .a(\u2_Display/n560 ),
    .b(\u2_Display/n594 [31]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n595 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1281 (
    .a(\u2_Display/n1714 ),
    .b(\u2_Display/n1717 [0]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1749 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1282 (
    .a(\u2_Display/n1713 ),
    .b(\u2_Display/n1717 [1]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1748 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1283 (
    .a(\u2_Display/n1712 ),
    .b(\u2_Display/n1717 [2]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1747 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1284 (
    .a(\u2_Display/n1711 ),
    .b(\u2_Display/n1717 [3]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1746 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1285 (
    .a(\u2_Display/n1710 ),
    .b(\u2_Display/n1717 [4]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1745 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1286 (
    .a(\u2_Display/n1709 ),
    .b(\u2_Display/n1717 [5]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1744 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1287 (
    .a(\u2_Display/n1708 ),
    .b(\u2_Display/n1717 [6]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1743 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1288 (
    .a(\u2_Display/n1707 ),
    .b(\u2_Display/n1717 [7]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1742 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1289 (
    .a(\u2_Display/n1706 ),
    .b(\u2_Display/n1717 [8]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1741 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1290 (
    .a(\u2_Display/n1705 ),
    .b(\u2_Display/n1717 [9]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1740 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1291 (
    .a(\u2_Display/n1704 ),
    .b(\u2_Display/n1717 [10]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1739 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1292 (
    .a(\u2_Display/n1703 ),
    .b(\u2_Display/n1717 [11]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1738 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1293 (
    .a(\u2_Display/n1702 ),
    .b(\u2_Display/n1717 [12]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1737 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1294 (
    .a(\u2_Display/n1701 ),
    .b(\u2_Display/n1717 [13]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1736 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1295 (
    .a(\u2_Display/n1700 ),
    .b(\u2_Display/n1717 [14]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1735 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1296 (
    .a(\u2_Display/n1699 ),
    .b(\u2_Display/n1717 [15]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1734 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1297 (
    .a(\u2_Display/n1698 ),
    .b(\u2_Display/n1717 [16]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1733 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1298 (
    .a(\u2_Display/n1697 ),
    .b(\u2_Display/n1717 [17]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1732 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1299 (
    .a(\u2_Display/n1696 ),
    .b(\u2_Display/n1717 [18]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1731 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1300 (
    .a(\u2_Display/n1695 ),
    .b(\u2_Display/n1717 [19]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1730 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1301 (
    .a(\u2_Display/n1694 ),
    .b(\u2_Display/n1717 [20]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1729 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1302 (
    .a(\u2_Display/n1693 ),
    .b(\u2_Display/n1717 [21]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1728 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1303 (
    .a(\u2_Display/n1692 ),
    .b(\u2_Display/n1717 [22]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1727 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1304 (
    .a(\u2_Display/n1691 ),
    .b(\u2_Display/n1717 [23]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1726 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1305 (
    .a(\u2_Display/n1690 ),
    .b(\u2_Display/n1717 [24]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1725 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1306 (
    .a(\u2_Display/n1689 ),
    .b(\u2_Display/n1717 [25]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1724 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1307 (
    .a(\u2_Display/n1688 ),
    .b(\u2_Display/n1717 [26]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1723 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1308 (
    .a(\u2_Display/n1687 ),
    .b(\u2_Display/n1717 [27]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1722 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1309 (
    .a(\u2_Display/n1686 ),
    .b(\u2_Display/n1717 [28]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1721 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1310 (
    .a(\u2_Display/n1685 ),
    .b(\u2_Display/n1717 [29]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1720 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1311 (
    .a(\u2_Display/n1684 ),
    .b(\u2_Display/n1717 [30]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1719 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1312 (
    .a(\u2_Display/n1683 ),
    .b(\u2_Display/n1717 [31]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1718 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1313 (
    .a(\u2_Display/n2837 ),
    .b(\u2_Display/n2840 [0]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2872 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1314 (
    .a(\u2_Display/n2836 ),
    .b(\u2_Display/n2840 [1]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2871 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1315 (
    .a(\u2_Display/n2835 ),
    .b(\u2_Display/n2840 [2]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2870 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1316 (
    .a(\u2_Display/n2834 ),
    .b(\u2_Display/n2840 [3]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2869 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1317 (
    .a(\u2_Display/n2833 ),
    .b(\u2_Display/n2840 [4]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2868 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1318 (
    .a(\u2_Display/n2832 ),
    .b(\u2_Display/n2840 [5]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2867 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1319 (
    .a(\u2_Display/n2831 ),
    .b(\u2_Display/n2840 [6]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2866 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1320 (
    .a(\u2_Display/n2830 ),
    .b(\u2_Display/n2840 [7]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2865 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1321 (
    .a(\u2_Display/n2829 ),
    .b(\u2_Display/n2840 [8]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2864 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1322 (
    .a(\u2_Display/n2828 ),
    .b(\u2_Display/n2840 [9]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2863 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1323 (
    .a(\u2_Display/n2827 ),
    .b(\u2_Display/n2840 [10]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2862 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1324 (
    .a(\u2_Display/n2826 ),
    .b(\u2_Display/n2840 [11]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2861 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1325 (
    .a(\u2_Display/n2825 ),
    .b(\u2_Display/n2840 [12]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2860 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1326 (
    .a(\u2_Display/n2824 ),
    .b(\u2_Display/n2840 [13]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2859 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1327 (
    .a(\u2_Display/n2823 ),
    .b(\u2_Display/n2840 [14]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2858 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1328 (
    .a(\u2_Display/n2822 ),
    .b(\u2_Display/n2840 [15]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2857 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1329 (
    .a(\u2_Display/n2821 ),
    .b(\u2_Display/n2840 [16]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2856 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1330 (
    .a(\u2_Display/n2820 ),
    .b(\u2_Display/n2840 [17]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2855 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1331 (
    .a(\u2_Display/n2819 ),
    .b(\u2_Display/n2840 [18]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2854 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1332 (
    .a(\u2_Display/n2818 ),
    .b(\u2_Display/n2840 [19]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2853 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1333 (
    .a(\u2_Display/n2817 ),
    .b(\u2_Display/n2840 [20]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2852 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1334 (
    .a(\u2_Display/n2816 ),
    .b(\u2_Display/n2840 [21]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2851 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1335 (
    .a(\u2_Display/n2815 ),
    .b(\u2_Display/n2840 [22]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2850 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1336 (
    .a(\u2_Display/n2814 ),
    .b(\u2_Display/n2840 [23]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2849 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1337 (
    .a(\u2_Display/n2813 ),
    .b(\u2_Display/n2840 [24]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2848 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1338 (
    .a(\u2_Display/n2812 ),
    .b(\u2_Display/n2840 [25]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2847 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1339 (
    .a(\u2_Display/n2811 ),
    .b(\u2_Display/n2840 [26]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2846 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1340 (
    .a(\u2_Display/n2810 ),
    .b(\u2_Display/n2840 [27]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2845 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1341 (
    .a(\u2_Display/n2809 ),
    .b(\u2_Display/n2840 [28]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2844 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1342 (
    .a(\u2_Display/n2808 ),
    .b(\u2_Display/n2840 [29]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2843 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1343 (
    .a(\u2_Display/n2807 ),
    .b(\u2_Display/n2840 [30]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2842 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1344 (
    .a(\u2_Display/n2806 ),
    .b(\u2_Display/n2840 [31]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2841 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1345 (
    .a(\u2_Display/n [27]),
    .b(\u2_Display/n [28]),
    .c(\u2_Display/n [29]),
    .d(\u2_Display/n [3]),
    .o(_al_u1345_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1346 (
    .a(\u2_Display/n [23]),
    .b(\u2_Display/n [24]),
    .c(\u2_Display/n [25]),
    .d(\u2_Display/n [26]),
    .o(_al_u1346_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u1347 (
    .a(\u2_Display/n [30]),
    .b(\u2_Display/n [4]),
    .c(\u2_Display/n [5]),
    .d(\u2_Display/n [6]),
    .o(_al_u1347_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u1348 (
    .a(_al_u1347_o),
    .b(\u2_Display/n [7]),
    .c(\u2_Display/n [8]),
    .d(\u2_Display/n [9]),
    .o(_al_u1348_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u1349 (
    .a(\u2_Display/n [12]),
    .b(\u2_Display/n [13]),
    .c(\u2_Display/n [14]),
    .d(\u2_Display/n [15]),
    .o(_al_u1349_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u1350 (
    .a(\u2_Display/n [0]),
    .b(\u2_Display/n [1]),
    .c(\u2_Display/n [10]),
    .d(\u2_Display/n [11]),
    .o(_al_u1350_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1351 (
    .a(\u2_Display/n [2]),
    .b(\u2_Display/n [20]),
    .c(\u2_Display/n [21]),
    .d(\u2_Display/n [22]),
    .o(_al_u1351_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1352 (
    .a(\u2_Display/n [16]),
    .b(\u2_Display/n [17]),
    .c(\u2_Display/n [18]),
    .d(\u2_Display/n [19]),
    .o(_al_u1352_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1353 (
    .a(_al_u1349_o),
    .b(_al_u1350_o),
    .c(_al_u1351_o),
    .d(_al_u1352_o),
    .o(_al_u1353_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1354 (
    .a(_al_u1353_o),
    .b(_al_u1348_o),
    .c(_al_u1345_o),
    .d(_al_u1346_o),
    .o(\u2_Display/n35 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1355 (
    .a(\u2_Display/n3995 ),
    .b(\u2_Display/n3998 [0]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4030 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1356 (
    .a(\u2_Display/n3994 ),
    .b(\u2_Display/n3998 [1]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4029 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1357 (
    .a(\u2_Display/n3993 ),
    .b(\u2_Display/n3998 [2]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4028 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1358 (
    .a(\u2_Display/n3992 ),
    .b(\u2_Display/n3998 [3]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4027 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1359 (
    .a(\u2_Display/n3991 ),
    .b(\u2_Display/n3998 [4]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4026 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1360 (
    .a(\u2_Display/n3990 ),
    .b(\u2_Display/n3998 [5]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4025 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1361 (
    .a(\u2_Display/n3989 ),
    .b(\u2_Display/n3998 [6]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4024 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1362 (
    .a(\u2_Display/n3988 ),
    .b(\u2_Display/n3998 [7]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4023 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1363 (
    .a(\u2_Display/n3987 ),
    .b(\u2_Display/n3998 [8]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4022 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1364 (
    .a(\u2_Display/n3986 ),
    .b(\u2_Display/n3998 [9]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4021 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1365 (
    .a(\u2_Display/n3985 ),
    .b(\u2_Display/n3998 [10]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4020 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1366 (
    .a(\u2_Display/n3984 ),
    .b(\u2_Display/n3998 [11]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4019 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1367 (
    .a(\u2_Display/n3983 ),
    .b(\u2_Display/n3998 [12]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4018 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1368 (
    .a(\u2_Display/n3982 ),
    .b(\u2_Display/n3998 [13]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4017 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1369 (
    .a(\u2_Display/n3981 ),
    .b(\u2_Display/n3998 [14]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4016 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1370 (
    .a(\u2_Display/n3980 ),
    .b(\u2_Display/n3998 [15]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4015 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1371 (
    .a(\u2_Display/n3979 ),
    .b(\u2_Display/n3998 [16]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4014 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1372 (
    .a(\u2_Display/n3978 ),
    .b(\u2_Display/n3998 [17]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4013 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1373 (
    .a(\u2_Display/n3977 ),
    .b(\u2_Display/n3998 [18]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4012 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1374 (
    .a(\u2_Display/n3976 ),
    .b(\u2_Display/n3998 [19]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4011 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1375 (
    .a(\u2_Display/n3975 ),
    .b(\u2_Display/n3998 [20]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4010 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1376 (
    .a(\u2_Display/n3974 ),
    .b(\u2_Display/n3998 [21]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4009 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1377 (
    .a(\u2_Display/n3973 ),
    .b(\u2_Display/n3998 [22]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4008 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1378 (
    .a(\u2_Display/n3972 ),
    .b(\u2_Display/n3998 [23]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4007 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1379 (
    .a(\u2_Display/n3971 ),
    .b(\u2_Display/n3998 [24]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4006 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1380 (
    .a(\u2_Display/n3970 ),
    .b(\u2_Display/n3998 [25]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4005 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1381 (
    .a(\u2_Display/n3969 ),
    .b(\u2_Display/n3998 [26]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4004 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1382 (
    .a(\u2_Display/n3968 ),
    .b(\u2_Display/n3998 [27]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4003 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1383 (
    .a(\u2_Display/n3967 ),
    .b(\u2_Display/n3998 [28]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4002 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1384 (
    .a(\u2_Display/n3966 ),
    .b(\u2_Display/n3998 [29]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4001 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1385 (
    .a(\u2_Display/n3965 ),
    .b(\u2_Display/n3998 [30]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4000 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1386 (
    .a(\u2_Display/n3964 ),
    .b(\u2_Display/n3998 [31]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n3999 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1387 (
    .a(\u2_Display/n6276 ),
    .b(\u2_Display/n5121 [0]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6311 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1388 (
    .a(\u2_Display/n6275 ),
    .b(\u2_Display/n5121 [1]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6310 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1389 (
    .a(\u2_Display/n6274 ),
    .b(\u2_Display/n5121 [2]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6309 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1390 (
    .a(\u2_Display/n6273 ),
    .b(\u2_Display/n5121 [3]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6308 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1391 (
    .a(\u2_Display/n6272 ),
    .b(\u2_Display/n5121 [4]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6307 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1392 (
    .a(\u2_Display/n6271 ),
    .b(\u2_Display/n5121 [5]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6306 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1393 (
    .a(\u2_Display/n6270 ),
    .b(\u2_Display/n5121 [6]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6305 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1394 (
    .a(\u2_Display/n6269 ),
    .b(\u2_Display/n5121 [7]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6304 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1395 (
    .a(\u2_Display/n6268 ),
    .b(\u2_Display/n5121 [8]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6303 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1396 (
    .a(\u2_Display/n6267 ),
    .b(\u2_Display/n5121 [9]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6302 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1397 (
    .a(\u2_Display/n6266 ),
    .b(\u2_Display/n5121 [10]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6301 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1398 (
    .a(\u2_Display/n6265 ),
    .b(\u2_Display/n5121 [11]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6300 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1399 (
    .a(\u2_Display/n6264 ),
    .b(\u2_Display/n5121 [12]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6299 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1400 (
    .a(\u2_Display/n6263 ),
    .b(\u2_Display/n5121 [13]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6298 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1401 (
    .a(\u2_Display/n6262 ),
    .b(\u2_Display/n5121 [14]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6297 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1402 (
    .a(\u2_Display/n6261 ),
    .b(\u2_Display/n5121 [15]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6296 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1403 (
    .a(\u2_Display/n6260 ),
    .b(\u2_Display/n5121 [16]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6295 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1404 (
    .a(\u2_Display/n6259 ),
    .b(\u2_Display/n5121 [17]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6294 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1405 (
    .a(\u2_Display/n6258 ),
    .b(\u2_Display/n5121 [18]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6293 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1406 (
    .a(\u2_Display/n6257 ),
    .b(\u2_Display/n5121 [19]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6292 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1407 (
    .a(\u2_Display/n6256 ),
    .b(\u2_Display/n5121 [20]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6291 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1408 (
    .a(\u2_Display/n6255 ),
    .b(\u2_Display/n5121 [21]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6290 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1409 (
    .a(\u2_Display/n6254 ),
    .b(\u2_Display/n5121 [22]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6289 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1410 (
    .a(\u2_Display/n6253 ),
    .b(\u2_Display/n5121 [23]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6288 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1411 (
    .a(\u2_Display/n6252 ),
    .b(\u2_Display/n5121 [24]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6287 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1412 (
    .a(\u2_Display/n6251 ),
    .b(\u2_Display/n5121 [25]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6286 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1413 (
    .a(\u2_Display/n6250 ),
    .b(\u2_Display/n5121 [26]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6285 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1414 (
    .a(\u2_Display/n6249 ),
    .b(\u2_Display/n5121 [27]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6284 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1415 (
    .a(\u2_Display/n6248 ),
    .b(\u2_Display/n5121 [28]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6283 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1416 (
    .a(\u2_Display/n6247 ),
    .b(\u2_Display/n5121 [29]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6282 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1417 (
    .a(\u2_Display/n6246 ),
    .b(\u2_Display/n5121 [30]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6281 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1418 (
    .a(\u2_Display/n6245 ),
    .b(\u2_Display/n5121 [31]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6280 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1419 (
    .a(\u2_Display/n626 ),
    .b(\u2_Display/n629 [0]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n661 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1420 (
    .a(\u2_Display/n625 ),
    .b(\u2_Display/n629 [1]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n660 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1421 (
    .a(\u2_Display/n624 ),
    .b(\u2_Display/n629 [2]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n659 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1422 (
    .a(\u2_Display/n623 ),
    .b(\u2_Display/n629 [3]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n658 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1423 (
    .a(\u2_Display/n622 ),
    .b(\u2_Display/n629 [4]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n657 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1424 (
    .a(\u2_Display/n621 ),
    .b(\u2_Display/n629 [5]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n656 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1425 (
    .a(\u2_Display/n620 ),
    .b(\u2_Display/n629 [6]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n655 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1426 (
    .a(\u2_Display/n619 ),
    .b(\u2_Display/n629 [7]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n654 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1427 (
    .a(\u2_Display/n618 ),
    .b(\u2_Display/n629 [8]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n653 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1428 (
    .a(\u2_Display/n617 ),
    .b(\u2_Display/n629 [9]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n652 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1429 (
    .a(\u2_Display/n616 ),
    .b(\u2_Display/n629 [10]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n651 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1430 (
    .a(\u2_Display/n615 ),
    .b(\u2_Display/n629 [11]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n650 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1431 (
    .a(\u2_Display/n614 ),
    .b(\u2_Display/n629 [12]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n649 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1432 (
    .a(\u2_Display/n613 ),
    .b(\u2_Display/n629 [13]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n648 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1433 (
    .a(\u2_Display/n612 ),
    .b(\u2_Display/n629 [14]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n647 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1434 (
    .a(\u2_Display/n611 ),
    .b(\u2_Display/n629 [15]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n646 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1435 (
    .a(\u2_Display/n610 ),
    .b(\u2_Display/n629 [16]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n645 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1436 (
    .a(\u2_Display/n609 ),
    .b(\u2_Display/n629 [17]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n644 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1437 (
    .a(\u2_Display/n608 ),
    .b(\u2_Display/n629 [18]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n643 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1438 (
    .a(\u2_Display/n607 ),
    .b(\u2_Display/n629 [19]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n642 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1439 (
    .a(\u2_Display/n606 ),
    .b(\u2_Display/n629 [20]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n641 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1440 (
    .a(\u2_Display/n605 ),
    .b(\u2_Display/n629 [21]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n640 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1441 (
    .a(\u2_Display/n604 ),
    .b(\u2_Display/n629 [22]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n639 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1442 (
    .a(\u2_Display/n603 ),
    .b(\u2_Display/n629 [23]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n638 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1443 (
    .a(\u2_Display/n602 ),
    .b(\u2_Display/n629 [24]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n637 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1444 (
    .a(\u2_Display/n601 ),
    .b(\u2_Display/n629 [25]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n636 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1445 (
    .a(\u2_Display/n600 ),
    .b(\u2_Display/n629 [26]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n635 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1446 (
    .a(\u2_Display/n599 ),
    .b(\u2_Display/n629 [27]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n634 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1447 (
    .a(\u2_Display/n598 ),
    .b(\u2_Display/n629 [28]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n633 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1448 (
    .a(\u2_Display/n597 ),
    .b(\u2_Display/n629 [29]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n632 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1449 (
    .a(\u2_Display/n596 ),
    .b(\u2_Display/n629 [30]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n631 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1450 (
    .a(\u2_Display/n595 ),
    .b(\u2_Display/n629 [31]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n630 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1451 (
    .a(\u2_Display/n1749 ),
    .b(\u2_Display/n1752 [0]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1784 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1452 (
    .a(\u2_Display/n1748 ),
    .b(\u2_Display/n1752 [1]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1783 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1453 (
    .a(\u2_Display/n1747 ),
    .b(\u2_Display/n1752 [2]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1782 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1454 (
    .a(\u2_Display/n1746 ),
    .b(\u2_Display/n1752 [3]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1781 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1455 (
    .a(\u2_Display/n1745 ),
    .b(\u2_Display/n1752 [4]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1780 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1456 (
    .a(\u2_Display/n1744 ),
    .b(\u2_Display/n1752 [5]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1779 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1457 (
    .a(\u2_Display/n1743 ),
    .b(\u2_Display/n1752 [6]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1778 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1458 (
    .a(\u2_Display/n1742 ),
    .b(\u2_Display/n1752 [7]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1777 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1459 (
    .a(\u2_Display/n1741 ),
    .b(\u2_Display/n1752 [8]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1776 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1460 (
    .a(\u2_Display/n1740 ),
    .b(\u2_Display/n1752 [9]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1775 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1461 (
    .a(\u2_Display/n1739 ),
    .b(\u2_Display/n1752 [10]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1774 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1462 (
    .a(\u2_Display/n1738 ),
    .b(\u2_Display/n1752 [11]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1773 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1463 (
    .a(\u2_Display/n1737 ),
    .b(\u2_Display/n1752 [12]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1772 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1464 (
    .a(\u2_Display/n1736 ),
    .b(\u2_Display/n1752 [13]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1771 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1465 (
    .a(\u2_Display/n1735 ),
    .b(\u2_Display/n1752 [14]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1770 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1466 (
    .a(\u2_Display/n1734 ),
    .b(\u2_Display/n1752 [15]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1769 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1467 (
    .a(\u2_Display/n1733 ),
    .b(\u2_Display/n1752 [16]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1768 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1468 (
    .a(\u2_Display/n1732 ),
    .b(\u2_Display/n1752 [17]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1767 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1469 (
    .a(\u2_Display/n1731 ),
    .b(\u2_Display/n1752 [18]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1766 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1470 (
    .a(\u2_Display/n1730 ),
    .b(\u2_Display/n1752 [19]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1765 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1471 (
    .a(\u2_Display/n1729 ),
    .b(\u2_Display/n1752 [20]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1764 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1472 (
    .a(\u2_Display/n1728 ),
    .b(\u2_Display/n1752 [21]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1763 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1473 (
    .a(\u2_Display/n1727 ),
    .b(\u2_Display/n1752 [22]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1762 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1474 (
    .a(\u2_Display/n1726 ),
    .b(\u2_Display/n1752 [23]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1761 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1475 (
    .a(\u2_Display/n1725 ),
    .b(\u2_Display/n1752 [24]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1760 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1476 (
    .a(\u2_Display/n1724 ),
    .b(\u2_Display/n1752 [25]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1759 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1477 (
    .a(\u2_Display/n1723 ),
    .b(\u2_Display/n1752 [26]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1758 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1478 (
    .a(\u2_Display/n1722 ),
    .b(\u2_Display/n1752 [27]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1757 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1479 (
    .a(\u2_Display/n1721 ),
    .b(\u2_Display/n1752 [28]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1756 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1480 (
    .a(\u2_Display/n1720 ),
    .b(\u2_Display/n1752 [29]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1755 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1481 (
    .a(\u2_Display/n1719 ),
    .b(\u2_Display/n1752 [30]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1754 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1482 (
    .a(\u2_Display/n1718 ),
    .b(\u2_Display/n1752 [31]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1753 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1483 (
    .a(\u2_Display/n2872 ),
    .b(\u2_Display/n2875 [0]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2907 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1484 (
    .a(\u2_Display/n2871 ),
    .b(\u2_Display/n2875 [1]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2906 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1485 (
    .a(\u2_Display/n2870 ),
    .b(\u2_Display/n2875 [2]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2905 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1486 (
    .a(\u2_Display/n2869 ),
    .b(\u2_Display/n2875 [3]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2904 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1487 (
    .a(\u2_Display/n2868 ),
    .b(\u2_Display/n2875 [4]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2903 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1488 (
    .a(\u2_Display/n2867 ),
    .b(\u2_Display/n2875 [5]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2902 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1489 (
    .a(\u2_Display/n2866 ),
    .b(\u2_Display/n2875 [6]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2901 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1490 (
    .a(\u2_Display/n2865 ),
    .b(\u2_Display/n2875 [7]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2900 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1491 (
    .a(\u2_Display/n2864 ),
    .b(\u2_Display/n2875 [8]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2899 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1492 (
    .a(\u2_Display/n2863 ),
    .b(\u2_Display/n2875 [9]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2898 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1493 (
    .a(\u2_Display/n2862 ),
    .b(\u2_Display/n2875 [10]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2897 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1494 (
    .a(\u2_Display/n2861 ),
    .b(\u2_Display/n2875 [11]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2896 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1495 (
    .a(\u2_Display/n2860 ),
    .b(\u2_Display/n2875 [12]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2895 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1496 (
    .a(\u2_Display/n2859 ),
    .b(\u2_Display/n2875 [13]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2894 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1497 (
    .a(\u2_Display/n2858 ),
    .b(\u2_Display/n2875 [14]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2893 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1498 (
    .a(\u2_Display/n2857 ),
    .b(\u2_Display/n2875 [15]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2892 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1499 (
    .a(\u2_Display/n2856 ),
    .b(\u2_Display/n2875 [16]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2891 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1500 (
    .a(\u2_Display/n2855 ),
    .b(\u2_Display/n2875 [17]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2890 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1501 (
    .a(\u2_Display/n2854 ),
    .b(\u2_Display/n2875 [18]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2889 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1502 (
    .a(\u2_Display/n2853 ),
    .b(\u2_Display/n2875 [19]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2888 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1503 (
    .a(\u2_Display/n2852 ),
    .b(\u2_Display/n2875 [20]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2887 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1504 (
    .a(\u2_Display/n2851 ),
    .b(\u2_Display/n2875 [21]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2886 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1505 (
    .a(\u2_Display/n2850 ),
    .b(\u2_Display/n2875 [22]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2885 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1506 (
    .a(\u2_Display/n2849 ),
    .b(\u2_Display/n2875 [23]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2884 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1507 (
    .a(\u2_Display/n2848 ),
    .b(\u2_Display/n2875 [24]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2883 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1508 (
    .a(\u2_Display/n2847 ),
    .b(\u2_Display/n2875 [25]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2882 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1509 (
    .a(\u2_Display/n2846 ),
    .b(\u2_Display/n2875 [26]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2881 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1510 (
    .a(\u2_Display/n2845 ),
    .b(\u2_Display/n2875 [27]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2880 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1511 (
    .a(\u2_Display/n2844 ),
    .b(\u2_Display/n2875 [28]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2879 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1512 (
    .a(\u2_Display/n2843 ),
    .b(\u2_Display/n2875 [29]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2878 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1513 (
    .a(\u2_Display/n2842 ),
    .b(\u2_Display/n2875 [30]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2877 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1514 (
    .a(\u2_Display/n2841 ),
    .b(\u2_Display/n2875 [31]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2876 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1515 (
    .a(\u2_Display/n4030 ),
    .b(\u2_Display/n4033 [0]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4065 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1516 (
    .a(\u2_Display/n4029 ),
    .b(\u2_Display/n4033 [1]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4064 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1517 (
    .a(\u2_Display/n4028 ),
    .b(\u2_Display/n4033 [2]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4063 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1518 (
    .a(\u2_Display/n4027 ),
    .b(\u2_Display/n4033 [3]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4062 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1519 (
    .a(\u2_Display/n4026 ),
    .b(\u2_Display/n4033 [4]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4061 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1520 (
    .a(\u2_Display/n4025 ),
    .b(\u2_Display/n4033 [5]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4060 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1521 (
    .a(\u2_Display/n4024 ),
    .b(\u2_Display/n4033 [6]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4059 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1522 (
    .a(\u2_Display/n4023 ),
    .b(\u2_Display/n4033 [7]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4058 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1523 (
    .a(\u2_Display/n4022 ),
    .b(\u2_Display/n4033 [8]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4057 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1524 (
    .a(\u2_Display/n4021 ),
    .b(\u2_Display/n4033 [9]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4056 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1525 (
    .a(\u2_Display/n4020 ),
    .b(\u2_Display/n4033 [10]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4055 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1526 (
    .a(\u2_Display/n4019 ),
    .b(\u2_Display/n4033 [11]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4054 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1527 (
    .a(\u2_Display/n4018 ),
    .b(\u2_Display/n4033 [12]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4053 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1528 (
    .a(\u2_Display/n4017 ),
    .b(\u2_Display/n4033 [13]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4052 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1529 (
    .a(\u2_Display/n4016 ),
    .b(\u2_Display/n4033 [14]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4051 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1530 (
    .a(\u2_Display/n4015 ),
    .b(\u2_Display/n4033 [15]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4050 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1531 (
    .a(\u2_Display/n4014 ),
    .b(\u2_Display/n4033 [16]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4049 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1532 (
    .a(\u2_Display/n4013 ),
    .b(\u2_Display/n4033 [17]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4048 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1533 (
    .a(\u2_Display/n4012 ),
    .b(\u2_Display/n4033 [18]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4047 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1534 (
    .a(\u2_Display/n4011 ),
    .b(\u2_Display/n4033 [19]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4046 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1535 (
    .a(\u2_Display/n4010 ),
    .b(\u2_Display/n4033 [20]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4045 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1536 (
    .a(\u2_Display/n4009 ),
    .b(\u2_Display/n4033 [21]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4044 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1537 (
    .a(\u2_Display/n4008 ),
    .b(\u2_Display/n4033 [22]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4043 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1538 (
    .a(\u2_Display/n4007 ),
    .b(\u2_Display/n4033 [23]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4042 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1539 (
    .a(\u2_Display/n4006 ),
    .b(\u2_Display/n4033 [24]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4041 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1540 (
    .a(\u2_Display/n4005 ),
    .b(\u2_Display/n4033 [25]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4040 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1541 (
    .a(\u2_Display/n4004 ),
    .b(\u2_Display/n4033 [26]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4039 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1542 (
    .a(\u2_Display/n4003 ),
    .b(\u2_Display/n4033 [27]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4038 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1543 (
    .a(\u2_Display/n4002 ),
    .b(\u2_Display/n4033 [28]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4037 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1544 (
    .a(\u2_Display/n4001 ),
    .b(\u2_Display/n4033 [29]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4036 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1545 (
    .a(\u2_Display/n4000 ),
    .b(\u2_Display/n4033 [30]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4035 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1546 (
    .a(\u2_Display/n3999 ),
    .b(\u2_Display/n4033 [31]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4034 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1547 (
    .a(\u2_Display/n6311 ),
    .b(\u2_Display/n5156 [0]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6346 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1548 (
    .a(\u2_Display/n6310 ),
    .b(\u2_Display/n5156 [1]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6345 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1549 (
    .a(\u2_Display/n6309 ),
    .b(\u2_Display/n5156 [2]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6344 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1550 (
    .a(\u2_Display/n6308 ),
    .b(\u2_Display/n5156 [3]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6343 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1551 (
    .a(\u2_Display/n6307 ),
    .b(\u2_Display/n5156 [4]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6342 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1552 (
    .a(\u2_Display/n6306 ),
    .b(\u2_Display/n5156 [5]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6341 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1553 (
    .a(\u2_Display/n6305 ),
    .b(\u2_Display/n5156 [6]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6340 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1554 (
    .a(\u2_Display/n6304 ),
    .b(\u2_Display/n5156 [7]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6339 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1555 (
    .a(\u2_Display/n6303 ),
    .b(\u2_Display/n5156 [8]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6338 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1556 (
    .a(\u2_Display/n6302 ),
    .b(\u2_Display/n5156 [9]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6337 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1557 (
    .a(\u2_Display/n6301 ),
    .b(\u2_Display/n5156 [10]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6336 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1558 (
    .a(\u2_Display/n6300 ),
    .b(\u2_Display/n5156 [11]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6335 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1559 (
    .a(\u2_Display/n6299 ),
    .b(\u2_Display/n5156 [12]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6334 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1560 (
    .a(\u2_Display/n6298 ),
    .b(\u2_Display/n5156 [13]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6333 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1561 (
    .a(\u2_Display/n6297 ),
    .b(\u2_Display/n5156 [14]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6332 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1562 (
    .a(\u2_Display/n6296 ),
    .b(\u2_Display/n5156 [15]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6331 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1563 (
    .a(\u2_Display/n6295 ),
    .b(\u2_Display/n5156 [16]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6330 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1564 (
    .a(\u2_Display/n6294 ),
    .b(\u2_Display/n5156 [17]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6329 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1565 (
    .a(\u2_Display/n6293 ),
    .b(\u2_Display/n5156 [18]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6328 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1566 (
    .a(\u2_Display/n6292 ),
    .b(\u2_Display/n5156 [19]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6327 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1567 (
    .a(\u2_Display/n6291 ),
    .b(\u2_Display/n5156 [20]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6326 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1568 (
    .a(\u2_Display/n6290 ),
    .b(\u2_Display/n5156 [21]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6325 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1569 (
    .a(\u2_Display/n6289 ),
    .b(\u2_Display/n5156 [22]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6324 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1570 (
    .a(\u2_Display/n6288 ),
    .b(\u2_Display/n5156 [23]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6323 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1571 (
    .a(\u2_Display/n6287 ),
    .b(\u2_Display/n5156 [24]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6322 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1572 (
    .a(\u2_Display/n6286 ),
    .b(\u2_Display/n5156 [25]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6321 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1573 (
    .a(\u2_Display/n6285 ),
    .b(\u2_Display/n5156 [26]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6320 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1574 (
    .a(\u2_Display/n6284 ),
    .b(\u2_Display/n5156 [27]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6319 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1575 (
    .a(\u2_Display/n6283 ),
    .b(\u2_Display/n5156 [28]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6318 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1576 (
    .a(\u2_Display/n6282 ),
    .b(\u2_Display/n5156 [29]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6317 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1577 (
    .a(\u2_Display/n6281 ),
    .b(\u2_Display/n5156 [30]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6316 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1578 (
    .a(\u2_Display/n6280 ),
    .b(\u2_Display/n5156 [31]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6315 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1579 (
    .a(\u2_Display/n661 ),
    .b(\u2_Display/n664 [0]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n696 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1580 (
    .a(\u2_Display/n660 ),
    .b(\u2_Display/n664 [1]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n695 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1581 (
    .a(\u2_Display/n659 ),
    .b(\u2_Display/n664 [2]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n694 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1582 (
    .a(\u2_Display/n658 ),
    .b(\u2_Display/n664 [3]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n693 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1583 (
    .a(\u2_Display/n657 ),
    .b(\u2_Display/n664 [4]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n692 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1584 (
    .a(\u2_Display/n656 ),
    .b(\u2_Display/n664 [5]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n691 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1585 (
    .a(\u2_Display/n655 ),
    .b(\u2_Display/n664 [6]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n690 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1586 (
    .a(\u2_Display/n654 ),
    .b(\u2_Display/n664 [7]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n689 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1587 (
    .a(\u2_Display/n653 ),
    .b(\u2_Display/n664 [8]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n688 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1588 (
    .a(\u2_Display/n652 ),
    .b(\u2_Display/n664 [9]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n687 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1589 (
    .a(\u2_Display/n651 ),
    .b(\u2_Display/n664 [10]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n686 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1590 (
    .a(\u2_Display/n650 ),
    .b(\u2_Display/n664 [11]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n685 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1591 (
    .a(\u2_Display/n649 ),
    .b(\u2_Display/n664 [12]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n684 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1592 (
    .a(\u2_Display/n648 ),
    .b(\u2_Display/n664 [13]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n683 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1593 (
    .a(\u2_Display/n647 ),
    .b(\u2_Display/n664 [14]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n682 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1594 (
    .a(\u2_Display/n646 ),
    .b(\u2_Display/n664 [15]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n681 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1595 (
    .a(\u2_Display/n645 ),
    .b(\u2_Display/n664 [16]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n680 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1596 (
    .a(\u2_Display/n644 ),
    .b(\u2_Display/n664 [17]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n679 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1597 (
    .a(\u2_Display/n643 ),
    .b(\u2_Display/n664 [18]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n678 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1598 (
    .a(\u2_Display/n642 ),
    .b(\u2_Display/n664 [19]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n677 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1599 (
    .a(\u2_Display/n641 ),
    .b(\u2_Display/n664 [20]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n676 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1600 (
    .a(\u2_Display/n640 ),
    .b(\u2_Display/n664 [21]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n675 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1601 (
    .a(\u2_Display/n639 ),
    .b(\u2_Display/n664 [22]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n674 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1602 (
    .a(\u2_Display/n638 ),
    .b(\u2_Display/n664 [23]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n673 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1603 (
    .a(\u2_Display/n637 ),
    .b(\u2_Display/n664 [24]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n672 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1604 (
    .a(\u2_Display/n636 ),
    .b(\u2_Display/n664 [25]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n671 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1605 (
    .a(\u2_Display/n635 ),
    .b(\u2_Display/n664 [26]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n670 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1606 (
    .a(\u2_Display/n634 ),
    .b(\u2_Display/n664 [27]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n669 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1607 (
    .a(\u2_Display/n633 ),
    .b(\u2_Display/n664 [28]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n668 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1608 (
    .a(\u2_Display/n632 ),
    .b(\u2_Display/n664 [29]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n667 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1609 (
    .a(\u2_Display/n631 ),
    .b(\u2_Display/n664 [30]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n666 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1610 (
    .a(\u2_Display/n630 ),
    .b(\u2_Display/n664 [31]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n665 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1611 (
    .a(\u2_Display/n1784 ),
    .b(\u2_Display/n1787 [0]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1819 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1612 (
    .a(\u2_Display/n1783 ),
    .b(\u2_Display/n1787 [1]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1818 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1613 (
    .a(\u2_Display/n1782 ),
    .b(\u2_Display/n1787 [2]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1817 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1614 (
    .a(\u2_Display/n1781 ),
    .b(\u2_Display/n1787 [3]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1816 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1615 (
    .a(\u2_Display/n1780 ),
    .b(\u2_Display/n1787 [4]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1815 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1616 (
    .a(\u2_Display/n1779 ),
    .b(\u2_Display/n1787 [5]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1814 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1617 (
    .a(\u2_Display/n1778 ),
    .b(\u2_Display/n1787 [6]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1813 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1618 (
    .a(\u2_Display/n1777 ),
    .b(\u2_Display/n1787 [7]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1812 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1619 (
    .a(\u2_Display/n1776 ),
    .b(\u2_Display/n1787 [8]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1811 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1620 (
    .a(\u2_Display/n1775 ),
    .b(\u2_Display/n1787 [9]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1810 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1621 (
    .a(\u2_Display/n1774 ),
    .b(\u2_Display/n1787 [10]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1809 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1622 (
    .a(\u2_Display/n1773 ),
    .b(\u2_Display/n1787 [11]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1808 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1623 (
    .a(\u2_Display/n1772 ),
    .b(\u2_Display/n1787 [12]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1807 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1624 (
    .a(\u2_Display/n1771 ),
    .b(\u2_Display/n1787 [13]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1806 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1625 (
    .a(\u2_Display/n1770 ),
    .b(\u2_Display/n1787 [14]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1805 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1626 (
    .a(\u2_Display/n1769 ),
    .b(\u2_Display/n1787 [15]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1804 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1627 (
    .a(\u2_Display/n1768 ),
    .b(\u2_Display/n1787 [16]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1803 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1628 (
    .a(\u2_Display/n1767 ),
    .b(\u2_Display/n1787 [17]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1802 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1629 (
    .a(\u2_Display/n1766 ),
    .b(\u2_Display/n1787 [18]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1801 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1630 (
    .a(\u2_Display/n1765 ),
    .b(\u2_Display/n1787 [19]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1800 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1631 (
    .a(\u2_Display/n1764 ),
    .b(\u2_Display/n1787 [20]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1799 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1632 (
    .a(\u2_Display/n1763 ),
    .b(\u2_Display/n1787 [21]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1798 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1633 (
    .a(\u2_Display/n1762 ),
    .b(\u2_Display/n1787 [22]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1797 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1634 (
    .a(\u2_Display/n1761 ),
    .b(\u2_Display/n1787 [23]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1796 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1635 (
    .a(\u2_Display/n1760 ),
    .b(\u2_Display/n1787 [24]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1795 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1636 (
    .a(\u2_Display/n1759 ),
    .b(\u2_Display/n1787 [25]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1794 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1637 (
    .a(\u2_Display/n1758 ),
    .b(\u2_Display/n1787 [26]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1793 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1638 (
    .a(\u2_Display/n1757 ),
    .b(\u2_Display/n1787 [27]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1792 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1639 (
    .a(\u2_Display/n1756 ),
    .b(\u2_Display/n1787 [28]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1791 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1640 (
    .a(\u2_Display/n1755 ),
    .b(\u2_Display/n1787 [29]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1790 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1641 (
    .a(\u2_Display/n1754 ),
    .b(\u2_Display/n1787 [30]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1789 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1642 (
    .a(\u2_Display/n1753 ),
    .b(\u2_Display/n1787 [31]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1788 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1643 (
    .a(\u2_Display/n2907 ),
    .b(\u2_Display/n2910 [0]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2942 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1644 (
    .a(\u2_Display/n2906 ),
    .b(\u2_Display/n2910 [1]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2941 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1645 (
    .a(\u2_Display/n2905 ),
    .b(\u2_Display/n2910 [2]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2940 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1646 (
    .a(\u2_Display/n2904 ),
    .b(\u2_Display/n2910 [3]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2939 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1647 (
    .a(\u2_Display/n2903 ),
    .b(\u2_Display/n2910 [4]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2938 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1648 (
    .a(\u2_Display/n2902 ),
    .b(\u2_Display/n2910 [5]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2937 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1649 (
    .a(\u2_Display/n2901 ),
    .b(\u2_Display/n2910 [6]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2936 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1650 (
    .a(\u2_Display/n2900 ),
    .b(\u2_Display/n2910 [7]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2935 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1651 (
    .a(\u2_Display/n2899 ),
    .b(\u2_Display/n2910 [8]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2934 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1652 (
    .a(\u2_Display/n2898 ),
    .b(\u2_Display/n2910 [9]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2933 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1653 (
    .a(\u2_Display/n2897 ),
    .b(\u2_Display/n2910 [10]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2932 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1654 (
    .a(\u2_Display/n2896 ),
    .b(\u2_Display/n2910 [11]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2931 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1655 (
    .a(\u2_Display/n2895 ),
    .b(\u2_Display/n2910 [12]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2930 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1656 (
    .a(\u2_Display/n2894 ),
    .b(\u2_Display/n2910 [13]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2929 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1657 (
    .a(\u2_Display/n2893 ),
    .b(\u2_Display/n2910 [14]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2928 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1658 (
    .a(\u2_Display/n2892 ),
    .b(\u2_Display/n2910 [15]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2927 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1659 (
    .a(\u2_Display/n2891 ),
    .b(\u2_Display/n2910 [16]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2926 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1660 (
    .a(\u2_Display/n2890 ),
    .b(\u2_Display/n2910 [17]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2925 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1661 (
    .a(\u2_Display/n2889 ),
    .b(\u2_Display/n2910 [18]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2924 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1662 (
    .a(\u2_Display/n2888 ),
    .b(\u2_Display/n2910 [19]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2923 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1663 (
    .a(\u2_Display/n2887 ),
    .b(\u2_Display/n2910 [20]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2922 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1664 (
    .a(\u2_Display/n2886 ),
    .b(\u2_Display/n2910 [21]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2921 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1665 (
    .a(\u2_Display/n2885 ),
    .b(\u2_Display/n2910 [22]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2920 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1666 (
    .a(\u2_Display/n2884 ),
    .b(\u2_Display/n2910 [23]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2919 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1667 (
    .a(\u2_Display/n2883 ),
    .b(\u2_Display/n2910 [24]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2918 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1668 (
    .a(\u2_Display/n2882 ),
    .b(\u2_Display/n2910 [25]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2917 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1669 (
    .a(\u2_Display/n2881 ),
    .b(\u2_Display/n2910 [26]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2916 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1670 (
    .a(\u2_Display/n2880 ),
    .b(\u2_Display/n2910 [27]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2915 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1671 (
    .a(\u2_Display/n2879 ),
    .b(\u2_Display/n2910 [28]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2914 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1672 (
    .a(\u2_Display/n2878 ),
    .b(\u2_Display/n2910 [29]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2913 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1673 (
    .a(\u2_Display/n2877 ),
    .b(\u2_Display/n2910 [30]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2912 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1674 (
    .a(\u2_Display/n2876 ),
    .b(\u2_Display/n2910 [31]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2911 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1675 (
    .a(\u2_Display/n4065 ),
    .b(\u2_Display/n4068 [0]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4100 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1676 (
    .a(\u2_Display/n4064 ),
    .b(\u2_Display/n4068 [1]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4099 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1677 (
    .a(\u2_Display/n4063 ),
    .b(\u2_Display/n4068 [2]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4098 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1678 (
    .a(\u2_Display/n4062 ),
    .b(\u2_Display/n4068 [3]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4097 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1679 (
    .a(\u2_Display/n4061 ),
    .b(\u2_Display/n4068 [4]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4096 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1680 (
    .a(\u2_Display/n4060 ),
    .b(\u2_Display/n4068 [5]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4095 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1681 (
    .a(\u2_Display/n4059 ),
    .b(\u2_Display/n4068 [6]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4094 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1682 (
    .a(\u2_Display/n4058 ),
    .b(\u2_Display/n4068 [7]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4093 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1683 (
    .a(\u2_Display/n4057 ),
    .b(\u2_Display/n4068 [8]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4092 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1684 (
    .a(\u2_Display/n4056 ),
    .b(\u2_Display/n4068 [9]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4091 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1685 (
    .a(\u2_Display/n4055 ),
    .b(\u2_Display/n4068 [10]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4090 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1686 (
    .a(\u2_Display/n4054 ),
    .b(\u2_Display/n4068 [11]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4089 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1687 (
    .a(\u2_Display/n4053 ),
    .b(\u2_Display/n4068 [12]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4088 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1688 (
    .a(\u2_Display/n4052 ),
    .b(\u2_Display/n4068 [13]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4087 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1689 (
    .a(\u2_Display/n4051 ),
    .b(\u2_Display/n4068 [14]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4086 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1690 (
    .a(\u2_Display/n4050 ),
    .b(\u2_Display/n4068 [15]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4085 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1691 (
    .a(\u2_Display/n4049 ),
    .b(\u2_Display/n4068 [16]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4084 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1692 (
    .a(\u2_Display/n4048 ),
    .b(\u2_Display/n4068 [17]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4083 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1693 (
    .a(\u2_Display/n4047 ),
    .b(\u2_Display/n4068 [18]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4082 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1694 (
    .a(\u2_Display/n4046 ),
    .b(\u2_Display/n4068 [19]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4081 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1695 (
    .a(\u2_Display/n4045 ),
    .b(\u2_Display/n4068 [20]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4080 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1696 (
    .a(\u2_Display/n4044 ),
    .b(\u2_Display/n4068 [21]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4079 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1697 (
    .a(\u2_Display/n4043 ),
    .b(\u2_Display/n4068 [22]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4078 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1698 (
    .a(\u2_Display/n4042 ),
    .b(\u2_Display/n4068 [23]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4077 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1699 (
    .a(\u2_Display/n4041 ),
    .b(\u2_Display/n4068 [24]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4076 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1700 (
    .a(\u2_Display/n4040 ),
    .b(\u2_Display/n4068 [25]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4075 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1701 (
    .a(\u2_Display/n4039 ),
    .b(\u2_Display/n4068 [26]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4074 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1702 (
    .a(\u2_Display/n4038 ),
    .b(\u2_Display/n4068 [27]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4073 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1703 (
    .a(\u2_Display/n4037 ),
    .b(\u2_Display/n4068 [28]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4072 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1704 (
    .a(\u2_Display/n4036 ),
    .b(\u2_Display/n4068 [29]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4071 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1705 (
    .a(\u2_Display/n4035 ),
    .b(\u2_Display/n4068 [30]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4070 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1706 (
    .a(\u2_Display/n4034 ),
    .b(\u2_Display/n4068 [31]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4069 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1707 (
    .a(\u2_Display/n6346 ),
    .b(\u2_Display/n5191 [0]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5223 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1708 (
    .a(\u2_Display/n6345 ),
    .b(\u2_Display/n5191 [1]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5222 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1709 (
    .a(\u2_Display/n6344 ),
    .b(\u2_Display/n5191 [2]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5221 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1710 (
    .a(\u2_Display/n6343 ),
    .b(\u2_Display/n5191 [3]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5220 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1711 (
    .a(\u2_Display/n6342 ),
    .b(\u2_Display/n5191 [4]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5219 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1712 (
    .a(\u2_Display/n6341 ),
    .b(\u2_Display/n5191 [5]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5218 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1713 (
    .a(\u2_Display/n6340 ),
    .b(\u2_Display/n5191 [6]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5217 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1714 (
    .a(\u2_Display/n6339 ),
    .b(\u2_Display/n5191 [7]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5216 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1715 (
    .a(\u2_Display/n6338 ),
    .b(\u2_Display/n5191 [8]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5215 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1716 (
    .a(\u2_Display/n6337 ),
    .b(\u2_Display/n5191 [9]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5214 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1717 (
    .a(\u2_Display/n6336 ),
    .b(\u2_Display/n5191 [10]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5213 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1718 (
    .a(\u2_Display/n6335 ),
    .b(\u2_Display/n5191 [11]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5212 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1719 (
    .a(\u2_Display/n6334 ),
    .b(\u2_Display/n5191 [12]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5211 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1720 (
    .a(\u2_Display/n6333 ),
    .b(\u2_Display/n5191 [13]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5210 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1721 (
    .a(\u2_Display/n6332 ),
    .b(\u2_Display/n5191 [14]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5209 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1722 (
    .a(\u2_Display/n6331 ),
    .b(\u2_Display/n5191 [15]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5208 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1723 (
    .a(\u2_Display/n6330 ),
    .b(\u2_Display/n5191 [16]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5207 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1724 (
    .a(\u2_Display/n6329 ),
    .b(\u2_Display/n5191 [17]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5206 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1725 (
    .a(\u2_Display/n6328 ),
    .b(\u2_Display/n5191 [18]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5205 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1726 (
    .a(\u2_Display/n6327 ),
    .b(\u2_Display/n5191 [19]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5204 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1727 (
    .a(\u2_Display/n6326 ),
    .b(\u2_Display/n5191 [20]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5203 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1728 (
    .a(\u2_Display/n6325 ),
    .b(\u2_Display/n5191 [21]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5202 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1729 (
    .a(\u2_Display/n6324 ),
    .b(\u2_Display/n5191 [22]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5201 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1730 (
    .a(\u2_Display/n6323 ),
    .b(\u2_Display/n5191 [23]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5200 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1731 (
    .a(\u2_Display/n6322 ),
    .b(\u2_Display/n5191 [24]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5199 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1732 (
    .a(\u2_Display/n6321 ),
    .b(\u2_Display/n5191 [25]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5198 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1733 (
    .a(\u2_Display/n6320 ),
    .b(\u2_Display/n5191 [26]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5197 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1734 (
    .a(\u2_Display/n6319 ),
    .b(\u2_Display/n5191 [27]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5196 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1735 (
    .a(\u2_Display/n6318 ),
    .b(\u2_Display/n5191 [28]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n6353 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1736 (
    .a(\u2_Display/n6317 ),
    .b(\u2_Display/n5191 [29]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n6352 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1737 (
    .a(\u2_Display/n6316 ),
    .b(\u2_Display/n5191 [30]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n6351 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1738 (
    .a(\u2_Display/n6315 ),
    .b(\u2_Display/n5191 [31]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n6350 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1739 (
    .a(\u2_Display/n696 ),
    .b(\u2_Display/n699 [0]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n731 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1740 (
    .a(\u2_Display/n695 ),
    .b(\u2_Display/n699 [1]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n730 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1741 (
    .a(\u2_Display/n694 ),
    .b(\u2_Display/n699 [2]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n729 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1742 (
    .a(\u2_Display/n693 ),
    .b(\u2_Display/n699 [3]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n728 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1743 (
    .a(\u2_Display/n692 ),
    .b(\u2_Display/n699 [4]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n727 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1744 (
    .a(\u2_Display/n691 ),
    .b(\u2_Display/n699 [5]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n726 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1745 (
    .a(\u2_Display/n690 ),
    .b(\u2_Display/n699 [6]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n725 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1746 (
    .a(\u2_Display/n689 ),
    .b(\u2_Display/n699 [7]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n724 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1747 (
    .a(\u2_Display/n688 ),
    .b(\u2_Display/n699 [8]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n723 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1748 (
    .a(\u2_Display/n687 ),
    .b(\u2_Display/n699 [9]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n722 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1749 (
    .a(\u2_Display/n686 ),
    .b(\u2_Display/n699 [10]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n721 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1750 (
    .a(\u2_Display/n685 ),
    .b(\u2_Display/n699 [11]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n720 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1751 (
    .a(\u2_Display/n684 ),
    .b(\u2_Display/n699 [12]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n719 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1752 (
    .a(\u2_Display/n683 ),
    .b(\u2_Display/n699 [13]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n718 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1753 (
    .a(\u2_Display/n682 ),
    .b(\u2_Display/n699 [14]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n717 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1754 (
    .a(\u2_Display/n681 ),
    .b(\u2_Display/n699 [15]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n716 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1755 (
    .a(\u2_Display/n680 ),
    .b(\u2_Display/n699 [16]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n715 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1756 (
    .a(\u2_Display/n679 ),
    .b(\u2_Display/n699 [17]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n714 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1757 (
    .a(\u2_Display/n678 ),
    .b(\u2_Display/n699 [18]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n713 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1758 (
    .a(\u2_Display/n677 ),
    .b(\u2_Display/n699 [19]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n712 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1759 (
    .a(\u2_Display/n676 ),
    .b(\u2_Display/n699 [20]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n711 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1760 (
    .a(\u2_Display/n675 ),
    .b(\u2_Display/n699 [21]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n710 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1761 (
    .a(\u2_Display/n674 ),
    .b(\u2_Display/n699 [22]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n709 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1762 (
    .a(\u2_Display/n673 ),
    .b(\u2_Display/n699 [23]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n708 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1763 (
    .a(\u2_Display/n672 ),
    .b(\u2_Display/n699 [24]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n707 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1764 (
    .a(\u2_Display/n671 ),
    .b(\u2_Display/n699 [25]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n706 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1765 (
    .a(\u2_Display/n670 ),
    .b(\u2_Display/n699 [26]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n705 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1766 (
    .a(\u2_Display/n669 ),
    .b(\u2_Display/n699 [27]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n704 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1767 (
    .a(\u2_Display/n668 ),
    .b(\u2_Display/n699 [28]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n703 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1768 (
    .a(\u2_Display/n667 ),
    .b(\u2_Display/n699 [29]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n702 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1769 (
    .a(\u2_Display/n666 ),
    .b(\u2_Display/n699 [30]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n701 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1770 (
    .a(\u2_Display/n665 ),
    .b(\u2_Display/n699 [31]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n700 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1771 (
    .a(\u2_Display/n1819 ),
    .b(\u2_Display/n1822 [0]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1854 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1772 (
    .a(\u2_Display/n1818 ),
    .b(\u2_Display/n1822 [1]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1853 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1773 (
    .a(\u2_Display/n1817 ),
    .b(\u2_Display/n1822 [2]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1852 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1774 (
    .a(\u2_Display/n1816 ),
    .b(\u2_Display/n1822 [3]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1851 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1775 (
    .a(\u2_Display/n1815 ),
    .b(\u2_Display/n1822 [4]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1850 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1776 (
    .a(\u2_Display/n1814 ),
    .b(\u2_Display/n1822 [5]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1849 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1777 (
    .a(\u2_Display/n1813 ),
    .b(\u2_Display/n1822 [6]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1848 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1778 (
    .a(\u2_Display/n1812 ),
    .b(\u2_Display/n1822 [7]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1847 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1779 (
    .a(\u2_Display/n1811 ),
    .b(\u2_Display/n1822 [8]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1846 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1780 (
    .a(\u2_Display/n1810 ),
    .b(\u2_Display/n1822 [9]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1845 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1781 (
    .a(\u2_Display/n1809 ),
    .b(\u2_Display/n1822 [10]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1844 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1782 (
    .a(\u2_Display/n1808 ),
    .b(\u2_Display/n1822 [11]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1843 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1783 (
    .a(\u2_Display/n1807 ),
    .b(\u2_Display/n1822 [12]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1842 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1784 (
    .a(\u2_Display/n1806 ),
    .b(\u2_Display/n1822 [13]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1841 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1785 (
    .a(\u2_Display/n1805 ),
    .b(\u2_Display/n1822 [14]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1840 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1786 (
    .a(\u2_Display/n1804 ),
    .b(\u2_Display/n1822 [15]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1839 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1787 (
    .a(\u2_Display/n1803 ),
    .b(\u2_Display/n1822 [16]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1838 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1788 (
    .a(\u2_Display/n1802 ),
    .b(\u2_Display/n1822 [17]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1837 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1789 (
    .a(\u2_Display/n1801 ),
    .b(\u2_Display/n1822 [18]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1836 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1790 (
    .a(\u2_Display/n1800 ),
    .b(\u2_Display/n1822 [19]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1835 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1791 (
    .a(\u2_Display/n1799 ),
    .b(\u2_Display/n1822 [20]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1834 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1792 (
    .a(\u2_Display/n1798 ),
    .b(\u2_Display/n1822 [21]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1833 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1793 (
    .a(\u2_Display/n1797 ),
    .b(\u2_Display/n1822 [22]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1832 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1794 (
    .a(\u2_Display/n1796 ),
    .b(\u2_Display/n1822 [23]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1831 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1795 (
    .a(\u2_Display/n1795 ),
    .b(\u2_Display/n1822 [24]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1830 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1796 (
    .a(\u2_Display/n1794 ),
    .b(\u2_Display/n1822 [25]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1829 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1797 (
    .a(\u2_Display/n1793 ),
    .b(\u2_Display/n1822 [26]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1828 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1798 (
    .a(\u2_Display/n1792 ),
    .b(\u2_Display/n1822 [27]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1827 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1799 (
    .a(\u2_Display/n1791 ),
    .b(\u2_Display/n1822 [28]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1826 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1800 (
    .a(\u2_Display/n1790 ),
    .b(\u2_Display/n1822 [29]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1825 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1801 (
    .a(\u2_Display/n1789 ),
    .b(\u2_Display/n1822 [30]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1824 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1802 (
    .a(\u2_Display/n1788 ),
    .b(\u2_Display/n1822 [31]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1823 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1803 (
    .a(\u2_Display/n2942 ),
    .b(\u2_Display/n2945 [0]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2977 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1804 (
    .a(\u2_Display/n2941 ),
    .b(\u2_Display/n2945 [1]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2976 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1805 (
    .a(\u2_Display/n2940 ),
    .b(\u2_Display/n2945 [2]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2975 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1806 (
    .a(\u2_Display/n2939 ),
    .b(\u2_Display/n2945 [3]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2974 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1807 (
    .a(\u2_Display/n2938 ),
    .b(\u2_Display/n2945 [4]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2973 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1808 (
    .a(\u2_Display/n2937 ),
    .b(\u2_Display/n2945 [5]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2972 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1809 (
    .a(\u2_Display/n2936 ),
    .b(\u2_Display/n2945 [6]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2971 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1810 (
    .a(\u2_Display/n2935 ),
    .b(\u2_Display/n2945 [7]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2970 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1811 (
    .a(\u2_Display/n2934 ),
    .b(\u2_Display/n2945 [8]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2969 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1812 (
    .a(\u2_Display/n2933 ),
    .b(\u2_Display/n2945 [9]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2968 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1813 (
    .a(\u2_Display/n2932 ),
    .b(\u2_Display/n2945 [10]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2967 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1814 (
    .a(\u2_Display/n2931 ),
    .b(\u2_Display/n2945 [11]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2966 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1815 (
    .a(\u2_Display/n2930 ),
    .b(\u2_Display/n2945 [12]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2965 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1816 (
    .a(\u2_Display/n2929 ),
    .b(\u2_Display/n2945 [13]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2964 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1817 (
    .a(\u2_Display/n2928 ),
    .b(\u2_Display/n2945 [14]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2963 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1818 (
    .a(\u2_Display/n2927 ),
    .b(\u2_Display/n2945 [15]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2962 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1819 (
    .a(\u2_Display/n2926 ),
    .b(\u2_Display/n2945 [16]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2961 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1820 (
    .a(\u2_Display/n2925 ),
    .b(\u2_Display/n2945 [17]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2960 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1821 (
    .a(\u2_Display/n2924 ),
    .b(\u2_Display/n2945 [18]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2959 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1822 (
    .a(\u2_Display/n2923 ),
    .b(\u2_Display/n2945 [19]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2958 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1823 (
    .a(\u2_Display/n2922 ),
    .b(\u2_Display/n2945 [20]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2957 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1824 (
    .a(\u2_Display/n2921 ),
    .b(\u2_Display/n2945 [21]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2956 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1825 (
    .a(\u2_Display/n2920 ),
    .b(\u2_Display/n2945 [22]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2955 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1826 (
    .a(\u2_Display/n2919 ),
    .b(\u2_Display/n2945 [23]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2954 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1827 (
    .a(\u2_Display/n2918 ),
    .b(\u2_Display/n2945 [24]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2953 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1828 (
    .a(\u2_Display/n2917 ),
    .b(\u2_Display/n2945 [25]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2952 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1829 (
    .a(\u2_Display/n2916 ),
    .b(\u2_Display/n2945 [26]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2951 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1830 (
    .a(\u2_Display/n2915 ),
    .b(\u2_Display/n2945 [27]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2950 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1831 (
    .a(\u2_Display/n2914 ),
    .b(\u2_Display/n2945 [28]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2949 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1832 (
    .a(\u2_Display/n2913 ),
    .b(\u2_Display/n2945 [29]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2948 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1833 (
    .a(\u2_Display/n2912 ),
    .b(\u2_Display/n2945 [30]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2947 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1834 (
    .a(\u2_Display/n2911 ),
    .b(\u2_Display/n2945 [31]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2946 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1835 (
    .a(\u2_Display/n4100 ),
    .b(\u2_Display/n4103 [0]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4135 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1836 (
    .a(\u2_Display/n4099 ),
    .b(\u2_Display/n4103 [1]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4134 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1837 (
    .a(\u2_Display/n4098 ),
    .b(\u2_Display/n4103 [2]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4133 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1838 (
    .a(\u2_Display/n4097 ),
    .b(\u2_Display/n4103 [3]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4132 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1839 (
    .a(\u2_Display/n4096 ),
    .b(\u2_Display/n4103 [4]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4131 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1840 (
    .a(\u2_Display/n4095 ),
    .b(\u2_Display/n4103 [5]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4130 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1841 (
    .a(\u2_Display/n4094 ),
    .b(\u2_Display/n4103 [6]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4129 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1842 (
    .a(\u2_Display/n4093 ),
    .b(\u2_Display/n4103 [7]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4128 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1843 (
    .a(\u2_Display/n4092 ),
    .b(\u2_Display/n4103 [8]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4127 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1844 (
    .a(\u2_Display/n4091 ),
    .b(\u2_Display/n4103 [9]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4126 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1845 (
    .a(\u2_Display/n4090 ),
    .b(\u2_Display/n4103 [10]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4125 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1846 (
    .a(\u2_Display/n4089 ),
    .b(\u2_Display/n4103 [11]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4124 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1847 (
    .a(\u2_Display/n4088 ),
    .b(\u2_Display/n4103 [12]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4123 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1848 (
    .a(\u2_Display/n4087 ),
    .b(\u2_Display/n4103 [13]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4122 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1849 (
    .a(\u2_Display/n4086 ),
    .b(\u2_Display/n4103 [14]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4121 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1850 (
    .a(\u2_Display/n4085 ),
    .b(\u2_Display/n4103 [15]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4120 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1851 (
    .a(\u2_Display/n4084 ),
    .b(\u2_Display/n4103 [16]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4119 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1852 (
    .a(\u2_Display/n4083 ),
    .b(\u2_Display/n4103 [17]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4118 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1853 (
    .a(\u2_Display/n4082 ),
    .b(\u2_Display/n4103 [18]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4117 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1854 (
    .a(\u2_Display/n4081 ),
    .b(\u2_Display/n4103 [19]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4116 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1855 (
    .a(\u2_Display/n4080 ),
    .b(\u2_Display/n4103 [20]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4115 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1856 (
    .a(\u2_Display/n4079 ),
    .b(\u2_Display/n4103 [21]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4114 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1857 (
    .a(\u2_Display/n4078 ),
    .b(\u2_Display/n4103 [22]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4113 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1858 (
    .a(\u2_Display/n4077 ),
    .b(\u2_Display/n4103 [23]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4112 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1859 (
    .a(\u2_Display/n4076 ),
    .b(\u2_Display/n4103 [24]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4111 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1860 (
    .a(\u2_Display/n4075 ),
    .b(\u2_Display/n4103 [25]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4110 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1861 (
    .a(\u2_Display/n4074 ),
    .b(\u2_Display/n4103 [26]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4109 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1862 (
    .a(\u2_Display/n4073 ),
    .b(\u2_Display/n4103 [27]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4108 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1863 (
    .a(\u2_Display/n4072 ),
    .b(\u2_Display/n4103 [28]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4107 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1864 (
    .a(\u2_Display/n4071 ),
    .b(\u2_Display/n4103 [29]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4106 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1865 (
    .a(\u2_Display/n4070 ),
    .b(\u2_Display/n4103 [30]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4105 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1866 (
    .a(\u2_Display/n4069 ),
    .b(\u2_Display/n4103 [31]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4104 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1867 (
    .a(\u2_Display/n5223 ),
    .b(\u2_Display/n5226 [0]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5258 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1868 (
    .a(\u2_Display/n5222 ),
    .b(\u2_Display/n5226 [1]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5257 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1869 (
    .a(\u2_Display/n5221 ),
    .b(\u2_Display/n5226 [2]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5256 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1870 (
    .a(\u2_Display/n5220 ),
    .b(\u2_Display/n5226 [3]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5255 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1871 (
    .a(\u2_Display/n5219 ),
    .b(\u2_Display/n5226 [4]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5254 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1872 (
    .a(\u2_Display/n5218 ),
    .b(\u2_Display/n5226 [5]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5253 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1873 (
    .a(\u2_Display/n5217 ),
    .b(\u2_Display/n5226 [6]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5252 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1874 (
    .a(\u2_Display/n5216 ),
    .b(\u2_Display/n5226 [7]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5251 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1875 (
    .a(\u2_Display/n5215 ),
    .b(\u2_Display/n5226 [8]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5250 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1876 (
    .a(\u2_Display/n5214 ),
    .b(\u2_Display/n5226 [9]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5249 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1877 (
    .a(\u2_Display/n5213 ),
    .b(\u2_Display/n5226 [10]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5248 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1878 (
    .a(\u2_Display/n5212 ),
    .b(\u2_Display/n5226 [11]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5247 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1879 (
    .a(\u2_Display/n5211 ),
    .b(\u2_Display/n5226 [12]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5246 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1880 (
    .a(\u2_Display/n5210 ),
    .b(\u2_Display/n5226 [13]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5245 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1881 (
    .a(\u2_Display/n5209 ),
    .b(\u2_Display/n5226 [14]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5244 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1882 (
    .a(\u2_Display/n5208 ),
    .b(\u2_Display/n5226 [15]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5243 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1883 (
    .a(\u2_Display/n5207 ),
    .b(\u2_Display/n5226 [16]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5242 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1884 (
    .a(\u2_Display/n5206 ),
    .b(\u2_Display/n5226 [17]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5241 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1885 (
    .a(\u2_Display/n5205 ),
    .b(\u2_Display/n5226 [18]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5240 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1886 (
    .a(\u2_Display/n5204 ),
    .b(\u2_Display/n5226 [19]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5239 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1887 (
    .a(\u2_Display/n5203 ),
    .b(\u2_Display/n5226 [20]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5238 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1888 (
    .a(\u2_Display/n5202 ),
    .b(\u2_Display/n5226 [21]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5237 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1889 (
    .a(\u2_Display/n5201 ),
    .b(\u2_Display/n5226 [22]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5236 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1890 (
    .a(\u2_Display/n5200 ),
    .b(\u2_Display/n5226 [23]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5235 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1891 (
    .a(\u2_Display/n5199 ),
    .b(\u2_Display/n5226 [24]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5234 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1892 (
    .a(\u2_Display/n5198 ),
    .b(\u2_Display/n5226 [25]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5233 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1893 (
    .a(\u2_Display/n5197 ),
    .b(\u2_Display/n5226 [26]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5232 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1894 (
    .a(\u2_Display/n5196 ),
    .b(\u2_Display/n5226 [27]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5231 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1895 (
    .a(\u2_Display/n6353 ),
    .b(\u2_Display/n5226 [28]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5230 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1896 (
    .a(\u2_Display/n6352 ),
    .b(\u2_Display/n5226 [29]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5229 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1897 (
    .a(\u2_Display/n6351 ),
    .b(\u2_Display/n5226 [30]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5228 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1898 (
    .a(\u2_Display/n6350 ),
    .b(\u2_Display/n5226 [31]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5227 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1899 (
    .a(\u2_Display/n731 ),
    .b(\u2_Display/n734 [0]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n766 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1900 (
    .a(\u2_Display/n730 ),
    .b(\u2_Display/n734 [1]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n765 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1901 (
    .a(\u2_Display/n729 ),
    .b(\u2_Display/n734 [2]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n764 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1902 (
    .a(\u2_Display/n728 ),
    .b(\u2_Display/n734 [3]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n763 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1903 (
    .a(\u2_Display/n727 ),
    .b(\u2_Display/n734 [4]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n762 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1904 (
    .a(\u2_Display/n726 ),
    .b(\u2_Display/n734 [5]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n761 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1905 (
    .a(\u2_Display/n725 ),
    .b(\u2_Display/n734 [6]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n760 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1906 (
    .a(\u2_Display/n724 ),
    .b(\u2_Display/n734 [7]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n759 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1907 (
    .a(\u2_Display/n723 ),
    .b(\u2_Display/n734 [8]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n758 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1908 (
    .a(\u2_Display/n722 ),
    .b(\u2_Display/n734 [9]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n757 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1909 (
    .a(\u2_Display/n721 ),
    .b(\u2_Display/n734 [10]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n756 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1910 (
    .a(\u2_Display/n720 ),
    .b(\u2_Display/n734 [11]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n755 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1911 (
    .a(\u2_Display/n719 ),
    .b(\u2_Display/n734 [12]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n754 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1912 (
    .a(\u2_Display/n718 ),
    .b(\u2_Display/n734 [13]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n753 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1913 (
    .a(\u2_Display/n717 ),
    .b(\u2_Display/n734 [14]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n752 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1914 (
    .a(\u2_Display/n716 ),
    .b(\u2_Display/n734 [15]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n751 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1915 (
    .a(\u2_Display/n715 ),
    .b(\u2_Display/n734 [16]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n750 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1916 (
    .a(\u2_Display/n714 ),
    .b(\u2_Display/n734 [17]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n749 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1917 (
    .a(\u2_Display/n713 ),
    .b(\u2_Display/n734 [18]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n748 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1918 (
    .a(\u2_Display/n712 ),
    .b(\u2_Display/n734 [19]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n747 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1919 (
    .a(\u2_Display/n711 ),
    .b(\u2_Display/n734 [20]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n746 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1920 (
    .a(\u2_Display/n710 ),
    .b(\u2_Display/n734 [21]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n745 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1921 (
    .a(\u2_Display/n709 ),
    .b(\u2_Display/n734 [22]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n744 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1922 (
    .a(\u2_Display/n708 ),
    .b(\u2_Display/n734 [23]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n743 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1923 (
    .a(\u2_Display/n707 ),
    .b(\u2_Display/n734 [24]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n742 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1924 (
    .a(\u2_Display/n706 ),
    .b(\u2_Display/n734 [25]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n741 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1925 (
    .a(\u2_Display/n705 ),
    .b(\u2_Display/n734 [26]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n740 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1926 (
    .a(\u2_Display/n704 ),
    .b(\u2_Display/n734 [27]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n739 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1927 (
    .a(\u2_Display/n703 ),
    .b(\u2_Display/n734 [28]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n738 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1928 (
    .a(\u2_Display/n702 ),
    .b(\u2_Display/n734 [29]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n737 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1929 (
    .a(\u2_Display/n701 ),
    .b(\u2_Display/n734 [30]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n736 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1930 (
    .a(\u2_Display/n700 ),
    .b(\u2_Display/n734 [31]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n735 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1931 (
    .a(\u2_Display/n1854 ),
    .b(\u2_Display/n1857 [0]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1889 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1932 (
    .a(\u2_Display/n1853 ),
    .b(\u2_Display/n1857 [1]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1888 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1933 (
    .a(\u2_Display/n1852 ),
    .b(\u2_Display/n1857 [2]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1887 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1934 (
    .a(\u2_Display/n1851 ),
    .b(\u2_Display/n1857 [3]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1886 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1935 (
    .a(\u2_Display/n1850 ),
    .b(\u2_Display/n1857 [4]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1885 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1936 (
    .a(\u2_Display/n1849 ),
    .b(\u2_Display/n1857 [5]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1884 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1937 (
    .a(\u2_Display/n1848 ),
    .b(\u2_Display/n1857 [6]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1883 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1938 (
    .a(\u2_Display/n1847 ),
    .b(\u2_Display/n1857 [7]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1882 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1939 (
    .a(\u2_Display/n1846 ),
    .b(\u2_Display/n1857 [8]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1881 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1940 (
    .a(\u2_Display/n1845 ),
    .b(\u2_Display/n1857 [9]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1880 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1941 (
    .a(\u2_Display/n1844 ),
    .b(\u2_Display/n1857 [10]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1879 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1942 (
    .a(\u2_Display/n1843 ),
    .b(\u2_Display/n1857 [11]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1878 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1943 (
    .a(\u2_Display/n1842 ),
    .b(\u2_Display/n1857 [12]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1877 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1944 (
    .a(\u2_Display/n1841 ),
    .b(\u2_Display/n1857 [13]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1876 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1945 (
    .a(\u2_Display/n1840 ),
    .b(\u2_Display/n1857 [14]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1875 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1946 (
    .a(\u2_Display/n1839 ),
    .b(\u2_Display/n1857 [15]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1874 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1947 (
    .a(\u2_Display/n1838 ),
    .b(\u2_Display/n1857 [16]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1873 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1948 (
    .a(\u2_Display/n1837 ),
    .b(\u2_Display/n1857 [17]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1872 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1949 (
    .a(\u2_Display/n1836 ),
    .b(\u2_Display/n1857 [18]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1871 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1950 (
    .a(\u2_Display/n1835 ),
    .b(\u2_Display/n1857 [19]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1870 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1951 (
    .a(\u2_Display/n1834 ),
    .b(\u2_Display/n1857 [20]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1869 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1952 (
    .a(\u2_Display/n1833 ),
    .b(\u2_Display/n1857 [21]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1868 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1953 (
    .a(\u2_Display/n1832 ),
    .b(\u2_Display/n1857 [22]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1867 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1954 (
    .a(\u2_Display/n1831 ),
    .b(\u2_Display/n1857 [23]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1866 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1955 (
    .a(\u2_Display/n1830 ),
    .b(\u2_Display/n1857 [24]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1865 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1956 (
    .a(\u2_Display/n1829 ),
    .b(\u2_Display/n1857 [25]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1864 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1957 (
    .a(\u2_Display/n1828 ),
    .b(\u2_Display/n1857 [26]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1863 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1958 (
    .a(\u2_Display/n1827 ),
    .b(\u2_Display/n1857 [27]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1862 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1959 (
    .a(\u2_Display/n1826 ),
    .b(\u2_Display/n1857 [28]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1861 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1960 (
    .a(\u2_Display/n1825 ),
    .b(\u2_Display/n1857 [29]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1860 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1961 (
    .a(\u2_Display/n1824 ),
    .b(\u2_Display/n1857 [30]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1859 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1962 (
    .a(\u2_Display/n1823 ),
    .b(\u2_Display/n1857 [31]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1858 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1963 (
    .a(\u2_Display/n2977 ),
    .b(\u2_Display/n2980 [0]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3012 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1964 (
    .a(\u2_Display/n2976 ),
    .b(\u2_Display/n2980 [1]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3011 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1965 (
    .a(\u2_Display/n2975 ),
    .b(\u2_Display/n2980 [2]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3010 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1966 (
    .a(\u2_Display/n2974 ),
    .b(\u2_Display/n2980 [3]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3009 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1967 (
    .a(\u2_Display/n2973 ),
    .b(\u2_Display/n2980 [4]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3008 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1968 (
    .a(\u2_Display/n2972 ),
    .b(\u2_Display/n2980 [5]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3007 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1969 (
    .a(\u2_Display/n2971 ),
    .b(\u2_Display/n2980 [6]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3006 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1970 (
    .a(\u2_Display/n2970 ),
    .b(\u2_Display/n2980 [7]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3005 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1971 (
    .a(\u2_Display/n2969 ),
    .b(\u2_Display/n2980 [8]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3004 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1972 (
    .a(\u2_Display/n2968 ),
    .b(\u2_Display/n2980 [9]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3003 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1973 (
    .a(\u2_Display/n2967 ),
    .b(\u2_Display/n2980 [10]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3002 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1974 (
    .a(\u2_Display/n2966 ),
    .b(\u2_Display/n2980 [11]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3001 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1975 (
    .a(\u2_Display/n2965 ),
    .b(\u2_Display/n2980 [12]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3000 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1976 (
    .a(\u2_Display/n2964 ),
    .b(\u2_Display/n2980 [13]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2999 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1977 (
    .a(\u2_Display/n2963 ),
    .b(\u2_Display/n2980 [14]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2998 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1978 (
    .a(\u2_Display/n2962 ),
    .b(\u2_Display/n2980 [15]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2997 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1979 (
    .a(\u2_Display/n2961 ),
    .b(\u2_Display/n2980 [16]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2996 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1980 (
    .a(\u2_Display/n2960 ),
    .b(\u2_Display/n2980 [17]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2995 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1981 (
    .a(\u2_Display/n2959 ),
    .b(\u2_Display/n2980 [18]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2994 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1982 (
    .a(\u2_Display/n2958 ),
    .b(\u2_Display/n2980 [19]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2993 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1983 (
    .a(\u2_Display/n2957 ),
    .b(\u2_Display/n2980 [20]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2992 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1984 (
    .a(\u2_Display/n2956 ),
    .b(\u2_Display/n2980 [21]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2991 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1985 (
    .a(\u2_Display/n2955 ),
    .b(\u2_Display/n2980 [22]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2990 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1986 (
    .a(\u2_Display/n2954 ),
    .b(\u2_Display/n2980 [23]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2989 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1987 (
    .a(\u2_Display/n2953 ),
    .b(\u2_Display/n2980 [24]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2988 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1988 (
    .a(\u2_Display/n2952 ),
    .b(\u2_Display/n2980 [25]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2987 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1989 (
    .a(\u2_Display/n2951 ),
    .b(\u2_Display/n2980 [26]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2986 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1990 (
    .a(\u2_Display/n2950 ),
    .b(\u2_Display/n2980 [27]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2985 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1991 (
    .a(\u2_Display/n2949 ),
    .b(\u2_Display/n2980 [28]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2984 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1992 (
    .a(\u2_Display/n2948 ),
    .b(\u2_Display/n2980 [29]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2983 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1993 (
    .a(\u2_Display/n2947 ),
    .b(\u2_Display/n2980 [30]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2982 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1994 (
    .a(\u2_Display/n2946 ),
    .b(\u2_Display/n2980 [31]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2981 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1995 (
    .a(\u2_Display/n4135 ),
    .b(\u2_Display/n4138 [0]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4170 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1996 (
    .a(\u2_Display/n4134 ),
    .b(\u2_Display/n4138 [1]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4169 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1997 (
    .a(\u2_Display/n4133 ),
    .b(\u2_Display/n4138 [2]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4168 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1998 (
    .a(\u2_Display/n4132 ),
    .b(\u2_Display/n4138 [3]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4167 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1999 (
    .a(\u2_Display/n4131 ),
    .b(\u2_Display/n4138 [4]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4166 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2000 (
    .a(\u2_Display/n4130 ),
    .b(\u2_Display/n4138 [5]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4165 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2001 (
    .a(\u2_Display/n4129 ),
    .b(\u2_Display/n4138 [6]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4164 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2002 (
    .a(\u2_Display/n4128 ),
    .b(\u2_Display/n4138 [7]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4163 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2003 (
    .a(\u2_Display/n4127 ),
    .b(\u2_Display/n4138 [8]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4162 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2004 (
    .a(\u2_Display/n4126 ),
    .b(\u2_Display/n4138 [9]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4161 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2005 (
    .a(\u2_Display/n4125 ),
    .b(\u2_Display/n4138 [10]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4160 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2006 (
    .a(\u2_Display/n4124 ),
    .b(\u2_Display/n4138 [11]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4159 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2007 (
    .a(\u2_Display/n4123 ),
    .b(\u2_Display/n4138 [12]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4158 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2008 (
    .a(\u2_Display/n4122 ),
    .b(\u2_Display/n4138 [13]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4157 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2009 (
    .a(\u2_Display/n4121 ),
    .b(\u2_Display/n4138 [14]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4156 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2010 (
    .a(\u2_Display/n4120 ),
    .b(\u2_Display/n4138 [15]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4155 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2011 (
    .a(\u2_Display/n4119 ),
    .b(\u2_Display/n4138 [16]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4154 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2012 (
    .a(\u2_Display/n4118 ),
    .b(\u2_Display/n4138 [17]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4153 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2013 (
    .a(\u2_Display/n4117 ),
    .b(\u2_Display/n4138 [18]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4152 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2014 (
    .a(\u2_Display/n4116 ),
    .b(\u2_Display/n4138 [19]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4151 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2015 (
    .a(\u2_Display/n4115 ),
    .b(\u2_Display/n4138 [20]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4150 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2016 (
    .a(\u2_Display/n4114 ),
    .b(\u2_Display/n4138 [21]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4149 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2017 (
    .a(\u2_Display/n4113 ),
    .b(\u2_Display/n4138 [22]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4148 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2018 (
    .a(\u2_Display/n4112 ),
    .b(\u2_Display/n4138 [23]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4147 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2019 (
    .a(\u2_Display/n4111 ),
    .b(\u2_Display/n4138 [24]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4146 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2020 (
    .a(\u2_Display/n4110 ),
    .b(\u2_Display/n4138 [25]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4145 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2021 (
    .a(\u2_Display/n4109 ),
    .b(\u2_Display/n4138 [26]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4144 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2022 (
    .a(\u2_Display/n4108 ),
    .b(\u2_Display/n4138 [27]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4143 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2023 (
    .a(\u2_Display/n4107 ),
    .b(\u2_Display/n4138 [28]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4142 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2024 (
    .a(\u2_Display/n4106 ),
    .b(\u2_Display/n4138 [29]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4141 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2025 (
    .a(\u2_Display/n4105 ),
    .b(\u2_Display/n4138 [30]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4140 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2026 (
    .a(\u2_Display/n4104 ),
    .b(\u2_Display/n4138 [31]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4139 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2027 (
    .a(\u2_Display/n5258 ),
    .b(\u2_Display/n5261 [0]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5293 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2028 (
    .a(\u2_Display/n5257 ),
    .b(\u2_Display/n5261 [1]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5292 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2029 (
    .a(\u2_Display/n5256 ),
    .b(\u2_Display/n5261 [2]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5291 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2030 (
    .a(\u2_Display/n5255 ),
    .b(\u2_Display/n5261 [3]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5290 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2031 (
    .a(\u2_Display/n5254 ),
    .b(\u2_Display/n5261 [4]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5289 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2032 (
    .a(\u2_Display/n5253 ),
    .b(\u2_Display/n5261 [5]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5288 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2033 (
    .a(\u2_Display/n5252 ),
    .b(\u2_Display/n5261 [6]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5287 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2034 (
    .a(\u2_Display/n5251 ),
    .b(\u2_Display/n5261 [7]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5286 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2035 (
    .a(\u2_Display/n5250 ),
    .b(\u2_Display/n5261 [8]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5285 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2036 (
    .a(\u2_Display/n5249 ),
    .b(\u2_Display/n5261 [9]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5284 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2037 (
    .a(\u2_Display/n5248 ),
    .b(\u2_Display/n5261 [10]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5283 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2038 (
    .a(\u2_Display/n5247 ),
    .b(\u2_Display/n5261 [11]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5282 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2039 (
    .a(\u2_Display/n5246 ),
    .b(\u2_Display/n5261 [12]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5281 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2040 (
    .a(\u2_Display/n5245 ),
    .b(\u2_Display/n5261 [13]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5280 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2041 (
    .a(\u2_Display/n5244 ),
    .b(\u2_Display/n5261 [14]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5279 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2042 (
    .a(\u2_Display/n5243 ),
    .b(\u2_Display/n5261 [15]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5278 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2043 (
    .a(\u2_Display/n5242 ),
    .b(\u2_Display/n5261 [16]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5277 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2044 (
    .a(\u2_Display/n5241 ),
    .b(\u2_Display/n5261 [17]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5276 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2045 (
    .a(\u2_Display/n5240 ),
    .b(\u2_Display/n5261 [18]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5275 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2046 (
    .a(\u2_Display/n5239 ),
    .b(\u2_Display/n5261 [19]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5274 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2047 (
    .a(\u2_Display/n5238 ),
    .b(\u2_Display/n5261 [20]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5273 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2048 (
    .a(\u2_Display/n5237 ),
    .b(\u2_Display/n5261 [21]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5272 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2049 (
    .a(\u2_Display/n5236 ),
    .b(\u2_Display/n5261 [22]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5271 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2050 (
    .a(\u2_Display/n5235 ),
    .b(\u2_Display/n5261 [23]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5270 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2051 (
    .a(\u2_Display/n5234 ),
    .b(\u2_Display/n5261 [24]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5269 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2052 (
    .a(\u2_Display/n5233 ),
    .b(\u2_Display/n5261 [25]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5268 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2053 (
    .a(\u2_Display/n5232 ),
    .b(\u2_Display/n5261 [26]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5267 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2054 (
    .a(\u2_Display/n5231 ),
    .b(\u2_Display/n5261 [27]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5266 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2055 (
    .a(\u2_Display/n5230 ),
    .b(\u2_Display/n5261 [28]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5265 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2056 (
    .a(\u2_Display/n5229 ),
    .b(\u2_Display/n5261 [29]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5264 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2057 (
    .a(\u2_Display/n5228 ),
    .b(\u2_Display/n5261 [30]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5263 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2058 (
    .a(\u2_Display/n5227 ),
    .b(\u2_Display/n5261 [31]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5262 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2059 (
    .a(\u2_Display/n766 ),
    .b(\u2_Display/n769 [0]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n801 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2060 (
    .a(\u2_Display/n765 ),
    .b(\u2_Display/n769 [1]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n800 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2061 (
    .a(\u2_Display/n764 ),
    .b(\u2_Display/n769 [2]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n799 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2062 (
    .a(\u2_Display/n763 ),
    .b(\u2_Display/n769 [3]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n798 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2063 (
    .a(\u2_Display/n762 ),
    .b(\u2_Display/n769 [4]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n797 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2064 (
    .a(\u2_Display/n761 ),
    .b(\u2_Display/n769 [5]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n796 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2065 (
    .a(\u2_Display/n760 ),
    .b(\u2_Display/n769 [6]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n795 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2066 (
    .a(\u2_Display/n759 ),
    .b(\u2_Display/n769 [7]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n794 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2067 (
    .a(\u2_Display/n758 ),
    .b(\u2_Display/n769 [8]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n793 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2068 (
    .a(\u2_Display/n757 ),
    .b(\u2_Display/n769 [9]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n792 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2069 (
    .a(\u2_Display/n756 ),
    .b(\u2_Display/n769 [10]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n791 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2070 (
    .a(\u2_Display/n755 ),
    .b(\u2_Display/n769 [11]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n790 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2071 (
    .a(\u2_Display/n754 ),
    .b(\u2_Display/n769 [12]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n789 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2072 (
    .a(\u2_Display/n753 ),
    .b(\u2_Display/n769 [13]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n788 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2073 (
    .a(\u2_Display/n752 ),
    .b(\u2_Display/n769 [14]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n787 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2074 (
    .a(\u2_Display/n751 ),
    .b(\u2_Display/n769 [15]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n786 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2075 (
    .a(\u2_Display/n750 ),
    .b(\u2_Display/n769 [16]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n785 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2076 (
    .a(\u2_Display/n749 ),
    .b(\u2_Display/n769 [17]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n784 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2077 (
    .a(\u2_Display/n748 ),
    .b(\u2_Display/n769 [18]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n783 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2078 (
    .a(\u2_Display/n747 ),
    .b(\u2_Display/n769 [19]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n782 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2079 (
    .a(\u2_Display/n746 ),
    .b(\u2_Display/n769 [20]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n781 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2080 (
    .a(\u2_Display/n745 ),
    .b(\u2_Display/n769 [21]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n780 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2081 (
    .a(\u2_Display/n744 ),
    .b(\u2_Display/n769 [22]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n779 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2082 (
    .a(\u2_Display/n743 ),
    .b(\u2_Display/n769 [23]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n778 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2083 (
    .a(\u2_Display/n742 ),
    .b(\u2_Display/n769 [24]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n777 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2084 (
    .a(\u2_Display/n741 ),
    .b(\u2_Display/n769 [25]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n776 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2085 (
    .a(\u2_Display/n740 ),
    .b(\u2_Display/n769 [26]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n775 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2086 (
    .a(\u2_Display/n739 ),
    .b(\u2_Display/n769 [27]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n774 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2087 (
    .a(\u2_Display/n738 ),
    .b(\u2_Display/n769 [28]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n773 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2088 (
    .a(\u2_Display/n737 ),
    .b(\u2_Display/n769 [29]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n772 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2089 (
    .a(\u2_Display/n736 ),
    .b(\u2_Display/n769 [30]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n771 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2090 (
    .a(\u2_Display/n735 ),
    .b(\u2_Display/n769 [31]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n770 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2091 (
    .a(\u2_Display/n1889 ),
    .b(\u2_Display/n1892 [0]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1924 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2092 (
    .a(\u2_Display/n1888 ),
    .b(\u2_Display/n1892 [1]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1923 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2093 (
    .a(\u2_Display/n1887 ),
    .b(\u2_Display/n1892 [2]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1922 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2094 (
    .a(\u2_Display/n1886 ),
    .b(\u2_Display/n1892 [3]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1921 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2095 (
    .a(\u2_Display/n1885 ),
    .b(\u2_Display/n1892 [4]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1920 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2096 (
    .a(\u2_Display/n1884 ),
    .b(\u2_Display/n1892 [5]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1919 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2097 (
    .a(\u2_Display/n1883 ),
    .b(\u2_Display/n1892 [6]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1918 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2098 (
    .a(\u2_Display/n1882 ),
    .b(\u2_Display/n1892 [7]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1917 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2099 (
    .a(\u2_Display/n1881 ),
    .b(\u2_Display/n1892 [8]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1916 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2100 (
    .a(\u2_Display/n1880 ),
    .b(\u2_Display/n1892 [9]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1915 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2101 (
    .a(\u2_Display/n1879 ),
    .b(\u2_Display/n1892 [10]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1914 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2102 (
    .a(\u2_Display/n1878 ),
    .b(\u2_Display/n1892 [11]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1913 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2103 (
    .a(\u2_Display/n1877 ),
    .b(\u2_Display/n1892 [12]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1912 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2104 (
    .a(\u2_Display/n1876 ),
    .b(\u2_Display/n1892 [13]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1911 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2105 (
    .a(\u2_Display/n1875 ),
    .b(\u2_Display/n1892 [14]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1910 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2106 (
    .a(\u2_Display/n1874 ),
    .b(\u2_Display/n1892 [15]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1909 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2107 (
    .a(\u2_Display/n1873 ),
    .b(\u2_Display/n1892 [16]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1908 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2108 (
    .a(\u2_Display/n1872 ),
    .b(\u2_Display/n1892 [17]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1907 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2109 (
    .a(\u2_Display/n1871 ),
    .b(\u2_Display/n1892 [18]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1906 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2110 (
    .a(\u2_Display/n1870 ),
    .b(\u2_Display/n1892 [19]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1905 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2111 (
    .a(\u2_Display/n1869 ),
    .b(\u2_Display/n1892 [20]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1904 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2112 (
    .a(\u2_Display/n1868 ),
    .b(\u2_Display/n1892 [21]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1903 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2113 (
    .a(\u2_Display/n1867 ),
    .b(\u2_Display/n1892 [22]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1902 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2114 (
    .a(\u2_Display/n1866 ),
    .b(\u2_Display/n1892 [23]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1901 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2115 (
    .a(\u2_Display/n1865 ),
    .b(\u2_Display/n1892 [24]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1900 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2116 (
    .a(\u2_Display/n1864 ),
    .b(\u2_Display/n1892 [25]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1899 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2117 (
    .a(\u2_Display/n1863 ),
    .b(\u2_Display/n1892 [26]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1898 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2118 (
    .a(\u2_Display/n1862 ),
    .b(\u2_Display/n1892 [27]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1897 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2119 (
    .a(\u2_Display/n1861 ),
    .b(\u2_Display/n1892 [28]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1896 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2120 (
    .a(\u2_Display/n1860 ),
    .b(\u2_Display/n1892 [29]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1895 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2121 (
    .a(\u2_Display/n1859 ),
    .b(\u2_Display/n1892 [30]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1894 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2122 (
    .a(\u2_Display/n1858 ),
    .b(\u2_Display/n1892 [31]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1893 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2123 (
    .a(\u2_Display/n3012 ),
    .b(\u2_Display/n3015 [0]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3047 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2124 (
    .a(\u2_Display/n3011 ),
    .b(\u2_Display/n3015 [1]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3046 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2125 (
    .a(\u2_Display/n3010 ),
    .b(\u2_Display/n3015 [2]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3045 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2126 (
    .a(\u2_Display/n3009 ),
    .b(\u2_Display/n3015 [3]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3044 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2127 (
    .a(\u2_Display/n3008 ),
    .b(\u2_Display/n3015 [4]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3043 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2128 (
    .a(\u2_Display/n3007 ),
    .b(\u2_Display/n3015 [5]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3042 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2129 (
    .a(\u2_Display/n3006 ),
    .b(\u2_Display/n3015 [6]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3041 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2130 (
    .a(\u2_Display/n3005 ),
    .b(\u2_Display/n3015 [7]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3040 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2131 (
    .a(\u2_Display/n3004 ),
    .b(\u2_Display/n3015 [8]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3039 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2132 (
    .a(\u2_Display/n3003 ),
    .b(\u2_Display/n3015 [9]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3038 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2133 (
    .a(\u2_Display/n3002 ),
    .b(\u2_Display/n3015 [10]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3037 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2134 (
    .a(\u2_Display/n3001 ),
    .b(\u2_Display/n3015 [11]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3036 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2135 (
    .a(\u2_Display/n3000 ),
    .b(\u2_Display/n3015 [12]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3035 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2136 (
    .a(\u2_Display/n2999 ),
    .b(\u2_Display/n3015 [13]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3034 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2137 (
    .a(\u2_Display/n2998 ),
    .b(\u2_Display/n3015 [14]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3033 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2138 (
    .a(\u2_Display/n2997 ),
    .b(\u2_Display/n3015 [15]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3032 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2139 (
    .a(\u2_Display/n2996 ),
    .b(\u2_Display/n3015 [16]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3031 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2140 (
    .a(\u2_Display/n2995 ),
    .b(\u2_Display/n3015 [17]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3030 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2141 (
    .a(\u2_Display/n2994 ),
    .b(\u2_Display/n3015 [18]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3029 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2142 (
    .a(\u2_Display/n2993 ),
    .b(\u2_Display/n3015 [19]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3028 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2143 (
    .a(\u2_Display/n2992 ),
    .b(\u2_Display/n3015 [20]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3027 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2144 (
    .a(\u2_Display/n2991 ),
    .b(\u2_Display/n3015 [21]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3026 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2145 (
    .a(\u2_Display/n2990 ),
    .b(\u2_Display/n3015 [22]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3025 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2146 (
    .a(\u2_Display/n2989 ),
    .b(\u2_Display/n3015 [23]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3024 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2147 (
    .a(\u2_Display/n2988 ),
    .b(\u2_Display/n3015 [24]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3023 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2148 (
    .a(\u2_Display/n2987 ),
    .b(\u2_Display/n3015 [25]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3022 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2149 (
    .a(\u2_Display/n2986 ),
    .b(\u2_Display/n3015 [26]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3021 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2150 (
    .a(\u2_Display/n2985 ),
    .b(\u2_Display/n3015 [27]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3020 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2151 (
    .a(\u2_Display/n2984 ),
    .b(\u2_Display/n3015 [28]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3019 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2152 (
    .a(\u2_Display/n2983 ),
    .b(\u2_Display/n3015 [29]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3018 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2153 (
    .a(\u2_Display/n2982 ),
    .b(\u2_Display/n3015 [30]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3017 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2154 (
    .a(\u2_Display/n2981 ),
    .b(\u2_Display/n3015 [31]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3016 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2155 (
    .a(\u2_Display/n4170 ),
    .b(\u2_Display/n4173 [0]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4205 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2156 (
    .a(\u2_Display/n4169 ),
    .b(\u2_Display/n4173 [1]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4204 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2157 (
    .a(\u2_Display/n4168 ),
    .b(\u2_Display/n4173 [2]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4203 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2158 (
    .a(\u2_Display/n4167 ),
    .b(\u2_Display/n4173 [3]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4202 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2159 (
    .a(\u2_Display/n4166 ),
    .b(\u2_Display/n4173 [4]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4201 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2160 (
    .a(\u2_Display/n4165 ),
    .b(\u2_Display/n4173 [5]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4200 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2161 (
    .a(\u2_Display/n4164 ),
    .b(\u2_Display/n4173 [6]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4199 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2162 (
    .a(\u2_Display/n4163 ),
    .b(\u2_Display/n4173 [7]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4198 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2163 (
    .a(\u2_Display/n4162 ),
    .b(\u2_Display/n4173 [8]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4197 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2164 (
    .a(\u2_Display/n4161 ),
    .b(\u2_Display/n4173 [9]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4196 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2165 (
    .a(\u2_Display/n4160 ),
    .b(\u2_Display/n4173 [10]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4195 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2166 (
    .a(\u2_Display/n4159 ),
    .b(\u2_Display/n4173 [11]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4194 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2167 (
    .a(\u2_Display/n4158 ),
    .b(\u2_Display/n4173 [12]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4193 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2168 (
    .a(\u2_Display/n4157 ),
    .b(\u2_Display/n4173 [13]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4192 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2169 (
    .a(\u2_Display/n4156 ),
    .b(\u2_Display/n4173 [14]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4191 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2170 (
    .a(\u2_Display/n4155 ),
    .b(\u2_Display/n4173 [15]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4190 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2171 (
    .a(\u2_Display/n4154 ),
    .b(\u2_Display/n4173 [16]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4189 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2172 (
    .a(\u2_Display/n4153 ),
    .b(\u2_Display/n4173 [17]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4188 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2173 (
    .a(\u2_Display/n4152 ),
    .b(\u2_Display/n4173 [18]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4187 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2174 (
    .a(\u2_Display/n4151 ),
    .b(\u2_Display/n4173 [19]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4186 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2175 (
    .a(\u2_Display/n4150 ),
    .b(\u2_Display/n4173 [20]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4185 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2176 (
    .a(\u2_Display/n4149 ),
    .b(\u2_Display/n4173 [21]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4184 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2177 (
    .a(\u2_Display/n4148 ),
    .b(\u2_Display/n4173 [22]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4183 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2178 (
    .a(\u2_Display/n4147 ),
    .b(\u2_Display/n4173 [23]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4182 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2179 (
    .a(\u2_Display/n4146 ),
    .b(\u2_Display/n4173 [24]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4181 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2180 (
    .a(\u2_Display/n4145 ),
    .b(\u2_Display/n4173 [25]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4180 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2181 (
    .a(\u2_Display/n4144 ),
    .b(\u2_Display/n4173 [26]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4179 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2182 (
    .a(\u2_Display/n4143 ),
    .b(\u2_Display/n4173 [27]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4178 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2183 (
    .a(\u2_Display/n4142 ),
    .b(\u2_Display/n4173 [28]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4177 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2184 (
    .a(\u2_Display/n4141 ),
    .b(\u2_Display/n4173 [29]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4176 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2185 (
    .a(\u2_Display/n4140 ),
    .b(\u2_Display/n4173 [30]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4175 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2186 (
    .a(\u2_Display/n4139 ),
    .b(\u2_Display/n4173 [31]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4174 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2187 (
    .a(\u2_Display/n5293 ),
    .b(\u2_Display/n5296 [0]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5328 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2188 (
    .a(\u2_Display/n5292 ),
    .b(\u2_Display/n5296 [1]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5327 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2189 (
    .a(\u2_Display/n5291 ),
    .b(\u2_Display/n5296 [2]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5326 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2190 (
    .a(\u2_Display/n5290 ),
    .b(\u2_Display/n5296 [3]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5325 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2191 (
    .a(\u2_Display/n5289 ),
    .b(\u2_Display/n5296 [4]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5324 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2192 (
    .a(\u2_Display/n5288 ),
    .b(\u2_Display/n5296 [5]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5323 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2193 (
    .a(\u2_Display/n5287 ),
    .b(\u2_Display/n5296 [6]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5322 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2194 (
    .a(\u2_Display/n5286 ),
    .b(\u2_Display/n5296 [7]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5321 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2195 (
    .a(\u2_Display/n5285 ),
    .b(\u2_Display/n5296 [8]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5320 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2196 (
    .a(\u2_Display/n5284 ),
    .b(\u2_Display/n5296 [9]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5319 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2197 (
    .a(\u2_Display/n5283 ),
    .b(\u2_Display/n5296 [10]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5318 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2198 (
    .a(\u2_Display/n5282 ),
    .b(\u2_Display/n5296 [11]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5317 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2199 (
    .a(\u2_Display/n5281 ),
    .b(\u2_Display/n5296 [12]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5316 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2200 (
    .a(\u2_Display/n5280 ),
    .b(\u2_Display/n5296 [13]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5315 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2201 (
    .a(\u2_Display/n5279 ),
    .b(\u2_Display/n5296 [14]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5314 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2202 (
    .a(\u2_Display/n5278 ),
    .b(\u2_Display/n5296 [15]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5313 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2203 (
    .a(\u2_Display/n5277 ),
    .b(\u2_Display/n5296 [16]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5312 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2204 (
    .a(\u2_Display/n5276 ),
    .b(\u2_Display/n5296 [17]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5311 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2205 (
    .a(\u2_Display/n5275 ),
    .b(\u2_Display/n5296 [18]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5310 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2206 (
    .a(\u2_Display/n5274 ),
    .b(\u2_Display/n5296 [19]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5309 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2207 (
    .a(\u2_Display/n5273 ),
    .b(\u2_Display/n5296 [20]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5308 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2208 (
    .a(\u2_Display/n5272 ),
    .b(\u2_Display/n5296 [21]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5307 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2209 (
    .a(\u2_Display/n5271 ),
    .b(\u2_Display/n5296 [22]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5306 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2210 (
    .a(\u2_Display/n5270 ),
    .b(\u2_Display/n5296 [23]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5305 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2211 (
    .a(\u2_Display/n5269 ),
    .b(\u2_Display/n5296 [24]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5304 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2212 (
    .a(\u2_Display/n5268 ),
    .b(\u2_Display/n5296 [25]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5303 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2213 (
    .a(\u2_Display/n5267 ),
    .b(\u2_Display/n5296 [26]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5302 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2214 (
    .a(\u2_Display/n5266 ),
    .b(\u2_Display/n5296 [27]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5301 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2215 (
    .a(\u2_Display/n5265 ),
    .b(\u2_Display/n5296 [28]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5300 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2216 (
    .a(\u2_Display/n5264 ),
    .b(\u2_Display/n5296 [29]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5299 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2217 (
    .a(\u2_Display/n5263 ),
    .b(\u2_Display/n5296 [30]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5298 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2218 (
    .a(\u2_Display/n5262 ),
    .b(\u2_Display/n5296 [31]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5297 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2219 (
    .a(\u2_Display/n801 ),
    .b(\u2_Display/n804 [0]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n836 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2220 (
    .a(\u2_Display/n800 ),
    .b(\u2_Display/n804 [1]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n835 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2221 (
    .a(\u2_Display/n799 ),
    .b(\u2_Display/n804 [2]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n834 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2222 (
    .a(\u2_Display/n798 ),
    .b(\u2_Display/n804 [3]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n833 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2223 (
    .a(\u2_Display/n797 ),
    .b(\u2_Display/n804 [4]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n832 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2224 (
    .a(\u2_Display/n796 ),
    .b(\u2_Display/n804 [5]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n831 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2225 (
    .a(\u2_Display/n795 ),
    .b(\u2_Display/n804 [6]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n830 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2226 (
    .a(\u2_Display/n794 ),
    .b(\u2_Display/n804 [7]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n829 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2227 (
    .a(\u2_Display/n793 ),
    .b(\u2_Display/n804 [8]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n828 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2228 (
    .a(\u2_Display/n792 ),
    .b(\u2_Display/n804 [9]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n827 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2229 (
    .a(\u2_Display/n791 ),
    .b(\u2_Display/n804 [10]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n826 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2230 (
    .a(\u2_Display/n790 ),
    .b(\u2_Display/n804 [11]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n825 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2231 (
    .a(\u2_Display/n789 ),
    .b(\u2_Display/n804 [12]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n824 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2232 (
    .a(\u2_Display/n788 ),
    .b(\u2_Display/n804 [13]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n823 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2233 (
    .a(\u2_Display/n787 ),
    .b(\u2_Display/n804 [14]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n822 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2234 (
    .a(\u2_Display/n786 ),
    .b(\u2_Display/n804 [15]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n821 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2235 (
    .a(\u2_Display/n785 ),
    .b(\u2_Display/n804 [16]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n820 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2236 (
    .a(\u2_Display/n784 ),
    .b(\u2_Display/n804 [17]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n819 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2237 (
    .a(\u2_Display/n783 ),
    .b(\u2_Display/n804 [18]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n818 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2238 (
    .a(\u2_Display/n782 ),
    .b(\u2_Display/n804 [19]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n817 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2239 (
    .a(\u2_Display/n781 ),
    .b(\u2_Display/n804 [20]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n816 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2240 (
    .a(\u2_Display/n780 ),
    .b(\u2_Display/n804 [21]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n815 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2241 (
    .a(\u2_Display/n779 ),
    .b(\u2_Display/n804 [22]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n814 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2242 (
    .a(\u2_Display/n778 ),
    .b(\u2_Display/n804 [23]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n813 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2243 (
    .a(\u2_Display/n777 ),
    .b(\u2_Display/n804 [24]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n812 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2244 (
    .a(\u2_Display/n776 ),
    .b(\u2_Display/n804 [25]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n811 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2245 (
    .a(\u2_Display/n775 ),
    .b(\u2_Display/n804 [26]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n810 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2246 (
    .a(\u2_Display/n774 ),
    .b(\u2_Display/n804 [27]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n809 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2247 (
    .a(\u2_Display/n773 ),
    .b(\u2_Display/n804 [28]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n808 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2248 (
    .a(\u2_Display/n772 ),
    .b(\u2_Display/n804 [29]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n807 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2249 (
    .a(\u2_Display/n771 ),
    .b(\u2_Display/n804 [30]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n806 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2250 (
    .a(\u2_Display/n770 ),
    .b(\u2_Display/n804 [31]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n805 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2251 (
    .a(\u2_Display/n1924 ),
    .b(\u2_Display/n1927 [0]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1959 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2252 (
    .a(\u2_Display/n1923 ),
    .b(\u2_Display/n1927 [1]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1958 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2253 (
    .a(\u2_Display/n1922 ),
    .b(\u2_Display/n1927 [2]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1957 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2254 (
    .a(\u2_Display/n1921 ),
    .b(\u2_Display/n1927 [3]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1956 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2255 (
    .a(\u2_Display/n1920 ),
    .b(\u2_Display/n1927 [4]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1955 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2256 (
    .a(\u2_Display/n1919 ),
    .b(\u2_Display/n1927 [5]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1954 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2257 (
    .a(\u2_Display/n1918 ),
    .b(\u2_Display/n1927 [6]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1953 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2258 (
    .a(\u2_Display/n1917 ),
    .b(\u2_Display/n1927 [7]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1952 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2259 (
    .a(\u2_Display/n1916 ),
    .b(\u2_Display/n1927 [8]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1951 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2260 (
    .a(\u2_Display/n1915 ),
    .b(\u2_Display/n1927 [9]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1950 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2261 (
    .a(\u2_Display/n1914 ),
    .b(\u2_Display/n1927 [10]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1949 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2262 (
    .a(\u2_Display/n1913 ),
    .b(\u2_Display/n1927 [11]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1948 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2263 (
    .a(\u2_Display/n1912 ),
    .b(\u2_Display/n1927 [12]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1947 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2264 (
    .a(\u2_Display/n1911 ),
    .b(\u2_Display/n1927 [13]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1946 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2265 (
    .a(\u2_Display/n1910 ),
    .b(\u2_Display/n1927 [14]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1945 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2266 (
    .a(\u2_Display/n1909 ),
    .b(\u2_Display/n1927 [15]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1944 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2267 (
    .a(\u2_Display/n1908 ),
    .b(\u2_Display/n1927 [16]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1943 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2268 (
    .a(\u2_Display/n1907 ),
    .b(\u2_Display/n1927 [17]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1942 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2269 (
    .a(\u2_Display/n1906 ),
    .b(\u2_Display/n1927 [18]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1941 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2270 (
    .a(\u2_Display/n1905 ),
    .b(\u2_Display/n1927 [19]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1940 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2271 (
    .a(\u2_Display/n1904 ),
    .b(\u2_Display/n1927 [20]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1939 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2272 (
    .a(\u2_Display/n1903 ),
    .b(\u2_Display/n1927 [21]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1938 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2273 (
    .a(\u2_Display/n1902 ),
    .b(\u2_Display/n1927 [22]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1937 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2274 (
    .a(\u2_Display/n1901 ),
    .b(\u2_Display/n1927 [23]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1936 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2275 (
    .a(\u2_Display/n1900 ),
    .b(\u2_Display/n1927 [24]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1935 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2276 (
    .a(\u2_Display/n1899 ),
    .b(\u2_Display/n1927 [25]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1934 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2277 (
    .a(\u2_Display/n1898 ),
    .b(\u2_Display/n1927 [26]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1933 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2278 (
    .a(\u2_Display/n1897 ),
    .b(\u2_Display/n1927 [27]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1932 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2279 (
    .a(\u2_Display/n1896 ),
    .b(\u2_Display/n1927 [28]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1931 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2280 (
    .a(\u2_Display/n1895 ),
    .b(\u2_Display/n1927 [29]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1930 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2281 (
    .a(\u2_Display/n1894 ),
    .b(\u2_Display/n1927 [30]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1929 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2282 (
    .a(\u2_Display/n1893 ),
    .b(\u2_Display/n1927 [31]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1928 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2283 (
    .a(\u2_Display/n3047 ),
    .b(\u2_Display/n3050 [0]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3082 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2284 (
    .a(\u2_Display/n3046 ),
    .b(\u2_Display/n3050 [1]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3081 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2285 (
    .a(\u2_Display/n3045 ),
    .b(\u2_Display/n3050 [2]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3080 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2286 (
    .a(\u2_Display/n3044 ),
    .b(\u2_Display/n3050 [3]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3079 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2287 (
    .a(\u2_Display/n3043 ),
    .b(\u2_Display/n3050 [4]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3078 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2288 (
    .a(\u2_Display/n3042 ),
    .b(\u2_Display/n3050 [5]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3077 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2289 (
    .a(\u2_Display/n3041 ),
    .b(\u2_Display/n3050 [6]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3076 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2290 (
    .a(\u2_Display/n3040 ),
    .b(\u2_Display/n3050 [7]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3075 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2291 (
    .a(\u2_Display/n3039 ),
    .b(\u2_Display/n3050 [8]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3074 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2292 (
    .a(\u2_Display/n3038 ),
    .b(\u2_Display/n3050 [9]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3073 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2293 (
    .a(\u2_Display/n3037 ),
    .b(\u2_Display/n3050 [10]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3072 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2294 (
    .a(\u2_Display/n3036 ),
    .b(\u2_Display/n3050 [11]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3071 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2295 (
    .a(\u2_Display/n3035 ),
    .b(\u2_Display/n3050 [12]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3070 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2296 (
    .a(\u2_Display/n3034 ),
    .b(\u2_Display/n3050 [13]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3069 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2297 (
    .a(\u2_Display/n3033 ),
    .b(\u2_Display/n3050 [14]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3068 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2298 (
    .a(\u2_Display/n3032 ),
    .b(\u2_Display/n3050 [15]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3067 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2299 (
    .a(\u2_Display/n3031 ),
    .b(\u2_Display/n3050 [16]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3066 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2300 (
    .a(\u2_Display/n3030 ),
    .b(\u2_Display/n3050 [17]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3065 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2301 (
    .a(\u2_Display/n3029 ),
    .b(\u2_Display/n3050 [18]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3064 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2302 (
    .a(\u2_Display/n3028 ),
    .b(\u2_Display/n3050 [19]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3063 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2303 (
    .a(\u2_Display/n3027 ),
    .b(\u2_Display/n3050 [20]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3062 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2304 (
    .a(\u2_Display/n3026 ),
    .b(\u2_Display/n3050 [21]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3061 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2305 (
    .a(\u2_Display/n3025 ),
    .b(\u2_Display/n3050 [22]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3060 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2306 (
    .a(\u2_Display/n3024 ),
    .b(\u2_Display/n3050 [23]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3059 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2307 (
    .a(\u2_Display/n3023 ),
    .b(\u2_Display/n3050 [24]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3058 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2308 (
    .a(\u2_Display/n3022 ),
    .b(\u2_Display/n3050 [25]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3057 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2309 (
    .a(\u2_Display/n3021 ),
    .b(\u2_Display/n3050 [26]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3056 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2310 (
    .a(\u2_Display/n3020 ),
    .b(\u2_Display/n3050 [27]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3055 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2311 (
    .a(\u2_Display/n3019 ),
    .b(\u2_Display/n3050 [28]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3054 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2312 (
    .a(\u2_Display/n3018 ),
    .b(\u2_Display/n3050 [29]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3053 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2313 (
    .a(\u2_Display/n3017 ),
    .b(\u2_Display/n3050 [30]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3052 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2314 (
    .a(\u2_Display/n3016 ),
    .b(\u2_Display/n3050 [31]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3051 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2315 (
    .a(\u2_Display/n4205 ),
    .b(\u2_Display/n4208 [0]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4240 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2316 (
    .a(\u2_Display/n4204 ),
    .b(\u2_Display/n4208 [1]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4239 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2317 (
    .a(\u2_Display/n4203 ),
    .b(\u2_Display/n4208 [2]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4238 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2318 (
    .a(\u2_Display/n4202 ),
    .b(\u2_Display/n4208 [3]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4237 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2319 (
    .a(\u2_Display/n4201 ),
    .b(\u2_Display/n4208 [4]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4236 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2320 (
    .a(\u2_Display/n4200 ),
    .b(\u2_Display/n4208 [5]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4235 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2321 (
    .a(\u2_Display/n4199 ),
    .b(\u2_Display/n4208 [6]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4234 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2322 (
    .a(\u2_Display/n4198 ),
    .b(\u2_Display/n4208 [7]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4233 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2323 (
    .a(\u2_Display/n4197 ),
    .b(\u2_Display/n4208 [8]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4232 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2324 (
    .a(\u2_Display/n4196 ),
    .b(\u2_Display/n4208 [9]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4231 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2325 (
    .a(\u2_Display/n4195 ),
    .b(\u2_Display/n4208 [10]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4230 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2326 (
    .a(\u2_Display/n4194 ),
    .b(\u2_Display/n4208 [11]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4229 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2327 (
    .a(\u2_Display/n4193 ),
    .b(\u2_Display/n4208 [12]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4228 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2328 (
    .a(\u2_Display/n4192 ),
    .b(\u2_Display/n4208 [13]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4227 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2329 (
    .a(\u2_Display/n4191 ),
    .b(\u2_Display/n4208 [14]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4226 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2330 (
    .a(\u2_Display/n4190 ),
    .b(\u2_Display/n4208 [15]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4225 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2331 (
    .a(\u2_Display/n4189 ),
    .b(\u2_Display/n4208 [16]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4224 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2332 (
    .a(\u2_Display/n4188 ),
    .b(\u2_Display/n4208 [17]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4223 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2333 (
    .a(\u2_Display/n4187 ),
    .b(\u2_Display/n4208 [18]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4222 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2334 (
    .a(\u2_Display/n4186 ),
    .b(\u2_Display/n4208 [19]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4221 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2335 (
    .a(\u2_Display/n4185 ),
    .b(\u2_Display/n4208 [20]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4220 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2336 (
    .a(\u2_Display/n4184 ),
    .b(\u2_Display/n4208 [21]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4219 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2337 (
    .a(\u2_Display/n4183 ),
    .b(\u2_Display/n4208 [22]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4218 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2338 (
    .a(\u2_Display/n4182 ),
    .b(\u2_Display/n4208 [23]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4217 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2339 (
    .a(\u2_Display/n4181 ),
    .b(\u2_Display/n4208 [24]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4216 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2340 (
    .a(\u2_Display/n4180 ),
    .b(\u2_Display/n4208 [25]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4215 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2341 (
    .a(\u2_Display/n4179 ),
    .b(\u2_Display/n4208 [26]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4214 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2342 (
    .a(\u2_Display/n4178 ),
    .b(\u2_Display/n4208 [27]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4213 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2343 (
    .a(\u2_Display/n4177 ),
    .b(\u2_Display/n4208 [28]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4212 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2344 (
    .a(\u2_Display/n4176 ),
    .b(\u2_Display/n4208 [29]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4211 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2345 (
    .a(\u2_Display/n4175 ),
    .b(\u2_Display/n4208 [30]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4210 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2346 (
    .a(\u2_Display/n4174 ),
    .b(\u2_Display/n4208 [31]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4209 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2347 (
    .a(\u2_Display/n5328 ),
    .b(\u2_Display/n5331 [0]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5363 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2348 (
    .a(\u2_Display/n5327 ),
    .b(\u2_Display/n5331 [1]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5362 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2349 (
    .a(\u2_Display/n5326 ),
    .b(\u2_Display/n5331 [2]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5361 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2350 (
    .a(\u2_Display/n5325 ),
    .b(\u2_Display/n5331 [3]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5360 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2351 (
    .a(\u2_Display/n5324 ),
    .b(\u2_Display/n5331 [4]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5359 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2352 (
    .a(\u2_Display/n5323 ),
    .b(\u2_Display/n5331 [5]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5358 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2353 (
    .a(\u2_Display/n5322 ),
    .b(\u2_Display/n5331 [6]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5357 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2354 (
    .a(\u2_Display/n5321 ),
    .b(\u2_Display/n5331 [7]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5356 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2355 (
    .a(\u2_Display/n5320 ),
    .b(\u2_Display/n5331 [8]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5355 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2356 (
    .a(\u2_Display/n5319 ),
    .b(\u2_Display/n5331 [9]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5354 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2357 (
    .a(\u2_Display/n5318 ),
    .b(\u2_Display/n5331 [10]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5353 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2358 (
    .a(\u2_Display/n5317 ),
    .b(\u2_Display/n5331 [11]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5352 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2359 (
    .a(\u2_Display/n5316 ),
    .b(\u2_Display/n5331 [12]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5351 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2360 (
    .a(\u2_Display/n5315 ),
    .b(\u2_Display/n5331 [13]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5350 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2361 (
    .a(\u2_Display/n5314 ),
    .b(\u2_Display/n5331 [14]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5349 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2362 (
    .a(\u2_Display/n5313 ),
    .b(\u2_Display/n5331 [15]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5348 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2363 (
    .a(\u2_Display/n5312 ),
    .b(\u2_Display/n5331 [16]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5347 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2364 (
    .a(\u2_Display/n5311 ),
    .b(\u2_Display/n5331 [17]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5346 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2365 (
    .a(\u2_Display/n5310 ),
    .b(\u2_Display/n5331 [18]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5345 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2366 (
    .a(\u2_Display/n5309 ),
    .b(\u2_Display/n5331 [19]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5344 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2367 (
    .a(\u2_Display/n5308 ),
    .b(\u2_Display/n5331 [20]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5343 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2368 (
    .a(\u2_Display/n5307 ),
    .b(\u2_Display/n5331 [21]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5342 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2369 (
    .a(\u2_Display/n5306 ),
    .b(\u2_Display/n5331 [22]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5341 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2370 (
    .a(\u2_Display/n5305 ),
    .b(\u2_Display/n5331 [23]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5340 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2371 (
    .a(\u2_Display/n5304 ),
    .b(\u2_Display/n5331 [24]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5339 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2372 (
    .a(\u2_Display/n5303 ),
    .b(\u2_Display/n5331 [25]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5338 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2373 (
    .a(\u2_Display/n5302 ),
    .b(\u2_Display/n5331 [26]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5337 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2374 (
    .a(\u2_Display/n5301 ),
    .b(\u2_Display/n5331 [27]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5336 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2375 (
    .a(\u2_Display/n5300 ),
    .b(\u2_Display/n5331 [28]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5335 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2376 (
    .a(\u2_Display/n5299 ),
    .b(\u2_Display/n5331 [29]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5334 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2377 (
    .a(\u2_Display/n5298 ),
    .b(\u2_Display/n5331 [30]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5333 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2378 (
    .a(\u2_Display/n5297 ),
    .b(\u2_Display/n5331 [31]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5332 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2379 (
    .a(\u2_Display/n836 ),
    .b(\u2_Display/n839 [0]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n871 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2380 (
    .a(\u2_Display/n835 ),
    .b(\u2_Display/n839 [1]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n870 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2381 (
    .a(\u2_Display/n834 ),
    .b(\u2_Display/n839 [2]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n869 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2382 (
    .a(\u2_Display/n833 ),
    .b(\u2_Display/n839 [3]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n868 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2383 (
    .a(\u2_Display/n832 ),
    .b(\u2_Display/n839 [4]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n867 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2384 (
    .a(\u2_Display/n831 ),
    .b(\u2_Display/n839 [5]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n866 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2385 (
    .a(\u2_Display/n830 ),
    .b(\u2_Display/n839 [6]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n865 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2386 (
    .a(\u2_Display/n829 ),
    .b(\u2_Display/n839 [7]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n864 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2387 (
    .a(\u2_Display/n828 ),
    .b(\u2_Display/n839 [8]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n863 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2388 (
    .a(\u2_Display/n827 ),
    .b(\u2_Display/n839 [9]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n862 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2389 (
    .a(\u2_Display/n826 ),
    .b(\u2_Display/n839 [10]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n861 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2390 (
    .a(\u2_Display/n825 ),
    .b(\u2_Display/n839 [11]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n860 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2391 (
    .a(\u2_Display/n824 ),
    .b(\u2_Display/n839 [12]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n859 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2392 (
    .a(\u2_Display/n823 ),
    .b(\u2_Display/n839 [13]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n858 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2393 (
    .a(\u2_Display/n822 ),
    .b(\u2_Display/n839 [14]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n857 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2394 (
    .a(\u2_Display/n821 ),
    .b(\u2_Display/n839 [15]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n856 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2395 (
    .a(\u2_Display/n820 ),
    .b(\u2_Display/n839 [16]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n855 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2396 (
    .a(\u2_Display/n819 ),
    .b(\u2_Display/n839 [17]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n854 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2397 (
    .a(\u2_Display/n818 ),
    .b(\u2_Display/n839 [18]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n853 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2398 (
    .a(\u2_Display/n817 ),
    .b(\u2_Display/n839 [19]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n852 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2399 (
    .a(\u2_Display/n816 ),
    .b(\u2_Display/n839 [20]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n851 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2400 (
    .a(\u2_Display/n815 ),
    .b(\u2_Display/n839 [21]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n850 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2401 (
    .a(\u2_Display/n814 ),
    .b(\u2_Display/n839 [22]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n849 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2402 (
    .a(\u2_Display/n813 ),
    .b(\u2_Display/n839 [23]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n848 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2403 (
    .a(\u2_Display/n812 ),
    .b(\u2_Display/n839 [24]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n847 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2404 (
    .a(\u2_Display/n811 ),
    .b(\u2_Display/n839 [25]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n846 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2405 (
    .a(\u2_Display/n810 ),
    .b(\u2_Display/n839 [26]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n845 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2406 (
    .a(\u2_Display/n809 ),
    .b(\u2_Display/n839 [27]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n844 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2407 (
    .a(\u2_Display/n808 ),
    .b(\u2_Display/n839 [28]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n843 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2408 (
    .a(\u2_Display/n807 ),
    .b(\u2_Display/n839 [29]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n842 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2409 (
    .a(\u2_Display/n806 ),
    .b(\u2_Display/n839 [30]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n841 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2410 (
    .a(\u2_Display/n805 ),
    .b(\u2_Display/n839 [31]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n840 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2411 (
    .a(\u2_Display/n1959 ),
    .b(\u2_Display/n1962 [0]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1994 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2412 (
    .a(\u2_Display/n1958 ),
    .b(\u2_Display/n1962 [1]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1993 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2413 (
    .a(\u2_Display/n1957 ),
    .b(\u2_Display/n1962 [2]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1992 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2414 (
    .a(\u2_Display/n1956 ),
    .b(\u2_Display/n1962 [3]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1991 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2415 (
    .a(\u2_Display/n1955 ),
    .b(\u2_Display/n1962 [4]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1990 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2416 (
    .a(\u2_Display/n1954 ),
    .b(\u2_Display/n1962 [5]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1989 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2417 (
    .a(\u2_Display/n1953 ),
    .b(\u2_Display/n1962 [6]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1988 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2418 (
    .a(\u2_Display/n1952 ),
    .b(\u2_Display/n1962 [7]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1987 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2419 (
    .a(\u2_Display/n1951 ),
    .b(\u2_Display/n1962 [8]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1986 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2420 (
    .a(\u2_Display/n1950 ),
    .b(\u2_Display/n1962 [9]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1985 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2421 (
    .a(\u2_Display/n1949 ),
    .b(\u2_Display/n1962 [10]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1984 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2422 (
    .a(\u2_Display/n1948 ),
    .b(\u2_Display/n1962 [11]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1983 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2423 (
    .a(\u2_Display/n1947 ),
    .b(\u2_Display/n1962 [12]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1982 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2424 (
    .a(\u2_Display/n1946 ),
    .b(\u2_Display/n1962 [13]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1981 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2425 (
    .a(\u2_Display/n1945 ),
    .b(\u2_Display/n1962 [14]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1980 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2426 (
    .a(\u2_Display/n1944 ),
    .b(\u2_Display/n1962 [15]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1979 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2427 (
    .a(\u2_Display/n1943 ),
    .b(\u2_Display/n1962 [16]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1978 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2428 (
    .a(\u2_Display/n1942 ),
    .b(\u2_Display/n1962 [17]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1977 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2429 (
    .a(\u2_Display/n1941 ),
    .b(\u2_Display/n1962 [18]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1976 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2430 (
    .a(\u2_Display/n1940 ),
    .b(\u2_Display/n1962 [19]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1975 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2431 (
    .a(\u2_Display/n1939 ),
    .b(\u2_Display/n1962 [20]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1974 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2432 (
    .a(\u2_Display/n1938 ),
    .b(\u2_Display/n1962 [21]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1973 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2433 (
    .a(\u2_Display/n1937 ),
    .b(\u2_Display/n1962 [22]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1972 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2434 (
    .a(\u2_Display/n1936 ),
    .b(\u2_Display/n1962 [23]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1971 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2435 (
    .a(\u2_Display/n1935 ),
    .b(\u2_Display/n1962 [24]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1970 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2436 (
    .a(\u2_Display/n1934 ),
    .b(\u2_Display/n1962 [25]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1969 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2437 (
    .a(\u2_Display/n1933 ),
    .b(\u2_Display/n1962 [26]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1968 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2438 (
    .a(\u2_Display/n1932 ),
    .b(\u2_Display/n1962 [27]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1967 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2439 (
    .a(\u2_Display/n1931 ),
    .b(\u2_Display/n1962 [28]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1966 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2440 (
    .a(\u2_Display/n1930 ),
    .b(\u2_Display/n1962 [29]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1965 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2441 (
    .a(\u2_Display/n1929 ),
    .b(\u2_Display/n1962 [30]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1964 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2442 (
    .a(\u2_Display/n1928 ),
    .b(\u2_Display/n1962 [31]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1963 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2443 (
    .a(\u2_Display/n3082 ),
    .b(\u2_Display/n3085 [0]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3117 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2444 (
    .a(\u2_Display/n3081 ),
    .b(\u2_Display/n3085 [1]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3116 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2445 (
    .a(\u2_Display/n3080 ),
    .b(\u2_Display/n3085 [2]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3115 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2446 (
    .a(\u2_Display/n3079 ),
    .b(\u2_Display/n3085 [3]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3114 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2447 (
    .a(\u2_Display/n3078 ),
    .b(\u2_Display/n3085 [4]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3113 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2448 (
    .a(\u2_Display/n3077 ),
    .b(\u2_Display/n3085 [5]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3112 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2449 (
    .a(\u2_Display/n3076 ),
    .b(\u2_Display/n3085 [6]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3111 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2450 (
    .a(\u2_Display/n3075 ),
    .b(\u2_Display/n3085 [7]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3110 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2451 (
    .a(\u2_Display/n3074 ),
    .b(\u2_Display/n3085 [8]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3109 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2452 (
    .a(\u2_Display/n3073 ),
    .b(\u2_Display/n3085 [9]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3108 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2453 (
    .a(\u2_Display/n3072 ),
    .b(\u2_Display/n3085 [10]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3107 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2454 (
    .a(\u2_Display/n3071 ),
    .b(\u2_Display/n3085 [11]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3106 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2455 (
    .a(\u2_Display/n3070 ),
    .b(\u2_Display/n3085 [12]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3105 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2456 (
    .a(\u2_Display/n3069 ),
    .b(\u2_Display/n3085 [13]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3104 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2457 (
    .a(\u2_Display/n3068 ),
    .b(\u2_Display/n3085 [14]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3103 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2458 (
    .a(\u2_Display/n3067 ),
    .b(\u2_Display/n3085 [15]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3102 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2459 (
    .a(\u2_Display/n3066 ),
    .b(\u2_Display/n3085 [16]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3101 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2460 (
    .a(\u2_Display/n3065 ),
    .b(\u2_Display/n3085 [17]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3100 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2461 (
    .a(\u2_Display/n3064 ),
    .b(\u2_Display/n3085 [18]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3099 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2462 (
    .a(\u2_Display/n3063 ),
    .b(\u2_Display/n3085 [19]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3098 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2463 (
    .a(\u2_Display/n3062 ),
    .b(\u2_Display/n3085 [20]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3097 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2464 (
    .a(\u2_Display/n3061 ),
    .b(\u2_Display/n3085 [21]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3096 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2465 (
    .a(\u2_Display/n3060 ),
    .b(\u2_Display/n3085 [22]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3095 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2466 (
    .a(\u2_Display/n3059 ),
    .b(\u2_Display/n3085 [23]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3094 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2467 (
    .a(\u2_Display/n3058 ),
    .b(\u2_Display/n3085 [24]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3093 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2468 (
    .a(\u2_Display/n3057 ),
    .b(\u2_Display/n3085 [25]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3092 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2469 (
    .a(\u2_Display/n3056 ),
    .b(\u2_Display/n3085 [26]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3091 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2470 (
    .a(\u2_Display/n3055 ),
    .b(\u2_Display/n3085 [27]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3090 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2471 (
    .a(\u2_Display/n3054 ),
    .b(\u2_Display/n3085 [28]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3089 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2472 (
    .a(\u2_Display/n3053 ),
    .b(\u2_Display/n3085 [29]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3088 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2473 (
    .a(\u2_Display/n3052 ),
    .b(\u2_Display/n3085 [30]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3087 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2474 (
    .a(\u2_Display/n3051 ),
    .b(\u2_Display/n3085 [31]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3086 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2475 (
    .a(\u2_Display/n4240 ),
    .b(\u2_Display/n4243 [0]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4275 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2476 (
    .a(\u2_Display/n4239 ),
    .b(\u2_Display/n4243 [1]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4274 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2477 (
    .a(\u2_Display/n4238 ),
    .b(\u2_Display/n4243 [2]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4273 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2478 (
    .a(\u2_Display/n4237 ),
    .b(\u2_Display/n4243 [3]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4272 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2479 (
    .a(\u2_Display/n4236 ),
    .b(\u2_Display/n4243 [4]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4271 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2480 (
    .a(\u2_Display/n4235 ),
    .b(\u2_Display/n4243 [5]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4270 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2481 (
    .a(\u2_Display/n4234 ),
    .b(\u2_Display/n4243 [6]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4269 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2482 (
    .a(\u2_Display/n4233 ),
    .b(\u2_Display/n4243 [7]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4268 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2483 (
    .a(\u2_Display/n4232 ),
    .b(\u2_Display/n4243 [8]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4267 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2484 (
    .a(\u2_Display/n4231 ),
    .b(\u2_Display/n4243 [9]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4266 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2485 (
    .a(\u2_Display/n4230 ),
    .b(\u2_Display/n4243 [10]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4265 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2486 (
    .a(\u2_Display/n4229 ),
    .b(\u2_Display/n4243 [11]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4264 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2487 (
    .a(\u2_Display/n4228 ),
    .b(\u2_Display/n4243 [12]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4263 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2488 (
    .a(\u2_Display/n4227 ),
    .b(\u2_Display/n4243 [13]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4262 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2489 (
    .a(\u2_Display/n4226 ),
    .b(\u2_Display/n4243 [14]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4261 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2490 (
    .a(\u2_Display/n4225 ),
    .b(\u2_Display/n4243 [15]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4260 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2491 (
    .a(\u2_Display/n4224 ),
    .b(\u2_Display/n4243 [16]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4259 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2492 (
    .a(\u2_Display/n4223 ),
    .b(\u2_Display/n4243 [17]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4258 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2493 (
    .a(\u2_Display/n4222 ),
    .b(\u2_Display/n4243 [18]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4257 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2494 (
    .a(\u2_Display/n4221 ),
    .b(\u2_Display/n4243 [19]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4256 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2495 (
    .a(\u2_Display/n4220 ),
    .b(\u2_Display/n4243 [20]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4255 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2496 (
    .a(\u2_Display/n4219 ),
    .b(\u2_Display/n4243 [21]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4254 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2497 (
    .a(\u2_Display/n4218 ),
    .b(\u2_Display/n4243 [22]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4253 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2498 (
    .a(\u2_Display/n4217 ),
    .b(\u2_Display/n4243 [23]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4252 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2499 (
    .a(\u2_Display/n4216 ),
    .b(\u2_Display/n4243 [24]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4251 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2500 (
    .a(\u2_Display/n4215 ),
    .b(\u2_Display/n4243 [25]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4250 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2501 (
    .a(\u2_Display/n4214 ),
    .b(\u2_Display/n4243 [26]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4249 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2502 (
    .a(\u2_Display/n4213 ),
    .b(\u2_Display/n4243 [27]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4248 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2503 (
    .a(\u2_Display/n4212 ),
    .b(\u2_Display/n4243 [28]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4247 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2504 (
    .a(\u2_Display/n4211 ),
    .b(\u2_Display/n4243 [29]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4246 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2505 (
    .a(\u2_Display/n4210 ),
    .b(\u2_Display/n4243 [30]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4245 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2506 (
    .a(\u2_Display/n4209 ),
    .b(\u2_Display/n4243 [31]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4244 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2507 (
    .a(\u2_Display/n5363 ),
    .b(\u2_Display/n5366 [0]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5398 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2508 (
    .a(\u2_Display/n5362 ),
    .b(\u2_Display/n5366 [1]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5397 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2509 (
    .a(\u2_Display/n5361 ),
    .b(\u2_Display/n5366 [2]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5396 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2510 (
    .a(\u2_Display/n5360 ),
    .b(\u2_Display/n5366 [3]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5395 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2511 (
    .a(\u2_Display/n5359 ),
    .b(\u2_Display/n5366 [4]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5394 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2512 (
    .a(\u2_Display/n5358 ),
    .b(\u2_Display/n5366 [5]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5393 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2513 (
    .a(\u2_Display/n5357 ),
    .b(\u2_Display/n5366 [6]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5392 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2514 (
    .a(\u2_Display/n5356 ),
    .b(\u2_Display/n5366 [7]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5391 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2515 (
    .a(\u2_Display/n5355 ),
    .b(\u2_Display/n5366 [8]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5390 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2516 (
    .a(\u2_Display/n5354 ),
    .b(\u2_Display/n5366 [9]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5389 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2517 (
    .a(\u2_Display/n5353 ),
    .b(\u2_Display/n5366 [10]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5388 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2518 (
    .a(\u2_Display/n5352 ),
    .b(\u2_Display/n5366 [11]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5387 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2519 (
    .a(\u2_Display/n5351 ),
    .b(\u2_Display/n5366 [12]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5386 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2520 (
    .a(\u2_Display/n5350 ),
    .b(\u2_Display/n5366 [13]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5385 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2521 (
    .a(\u2_Display/n5349 ),
    .b(\u2_Display/n5366 [14]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5384 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2522 (
    .a(\u2_Display/n5348 ),
    .b(\u2_Display/n5366 [15]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5383 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2523 (
    .a(\u2_Display/n5347 ),
    .b(\u2_Display/n5366 [16]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5382 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2524 (
    .a(\u2_Display/n5346 ),
    .b(\u2_Display/n5366 [17]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5381 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2525 (
    .a(\u2_Display/n5345 ),
    .b(\u2_Display/n5366 [18]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5380 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2526 (
    .a(\u2_Display/n5344 ),
    .b(\u2_Display/n5366 [19]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5379 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2527 (
    .a(\u2_Display/n5343 ),
    .b(\u2_Display/n5366 [20]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5378 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2528 (
    .a(\u2_Display/n5342 ),
    .b(\u2_Display/n5366 [21]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5377 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2529 (
    .a(\u2_Display/n5341 ),
    .b(\u2_Display/n5366 [22]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5376 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2530 (
    .a(\u2_Display/n5340 ),
    .b(\u2_Display/n5366 [23]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5375 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2531 (
    .a(\u2_Display/n5339 ),
    .b(\u2_Display/n5366 [24]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5374 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2532 (
    .a(\u2_Display/n5338 ),
    .b(\u2_Display/n5366 [25]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5373 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2533 (
    .a(\u2_Display/n5337 ),
    .b(\u2_Display/n5366 [26]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5372 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2534 (
    .a(\u2_Display/n5336 ),
    .b(\u2_Display/n5366 [27]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5371 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2535 (
    .a(\u2_Display/n5335 ),
    .b(\u2_Display/n5366 [28]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5370 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2536 (
    .a(\u2_Display/n5334 ),
    .b(\u2_Display/n5366 [29]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5369 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2537 (
    .a(\u2_Display/n5333 ),
    .b(\u2_Display/n5366 [30]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5368 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2538 (
    .a(\u2_Display/n5332 ),
    .b(\u2_Display/n5366 [31]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5367 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2539 (
    .a(\u2_Display/n871 ),
    .b(\u2_Display/n874 [0]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n906 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2540 (
    .a(\u2_Display/n870 ),
    .b(\u2_Display/n874 [1]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n905 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2541 (
    .a(\u2_Display/n869 ),
    .b(\u2_Display/n874 [2]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n904 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2542 (
    .a(\u2_Display/n868 ),
    .b(\u2_Display/n874 [3]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n903 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2543 (
    .a(\u2_Display/n867 ),
    .b(\u2_Display/n874 [4]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n902 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2544 (
    .a(\u2_Display/n866 ),
    .b(\u2_Display/n874 [5]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n901 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2545 (
    .a(\u2_Display/n865 ),
    .b(\u2_Display/n874 [6]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n900 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2546 (
    .a(\u2_Display/n864 ),
    .b(\u2_Display/n874 [7]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n899 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2547 (
    .a(\u2_Display/n863 ),
    .b(\u2_Display/n874 [8]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n898 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2548 (
    .a(\u2_Display/n862 ),
    .b(\u2_Display/n874 [9]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n897 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2549 (
    .a(\u2_Display/n861 ),
    .b(\u2_Display/n874 [10]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n896 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2550 (
    .a(\u2_Display/n860 ),
    .b(\u2_Display/n874 [11]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n895 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2551 (
    .a(\u2_Display/n859 ),
    .b(\u2_Display/n874 [12]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n894 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2552 (
    .a(\u2_Display/n858 ),
    .b(\u2_Display/n874 [13]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n893 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2553 (
    .a(\u2_Display/n857 ),
    .b(\u2_Display/n874 [14]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n892 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2554 (
    .a(\u2_Display/n856 ),
    .b(\u2_Display/n874 [15]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n891 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2555 (
    .a(\u2_Display/n855 ),
    .b(\u2_Display/n874 [16]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n890 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2556 (
    .a(\u2_Display/n854 ),
    .b(\u2_Display/n874 [17]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n889 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2557 (
    .a(\u2_Display/n853 ),
    .b(\u2_Display/n874 [18]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n888 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2558 (
    .a(\u2_Display/n852 ),
    .b(\u2_Display/n874 [19]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n887 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2559 (
    .a(\u2_Display/n851 ),
    .b(\u2_Display/n874 [20]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n886 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2560 (
    .a(\u2_Display/n850 ),
    .b(\u2_Display/n874 [21]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n885 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2561 (
    .a(\u2_Display/n849 ),
    .b(\u2_Display/n874 [22]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n884 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2562 (
    .a(\u2_Display/n848 ),
    .b(\u2_Display/n874 [23]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n883 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2563 (
    .a(\u2_Display/n847 ),
    .b(\u2_Display/n874 [24]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n882 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2564 (
    .a(\u2_Display/n846 ),
    .b(\u2_Display/n874 [25]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n881 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2565 (
    .a(\u2_Display/n845 ),
    .b(\u2_Display/n874 [26]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n880 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2566 (
    .a(\u2_Display/n844 ),
    .b(\u2_Display/n874 [27]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n879 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2567 (
    .a(\u2_Display/n843 ),
    .b(\u2_Display/n874 [28]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n878 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2568 (
    .a(\u2_Display/n842 ),
    .b(\u2_Display/n874 [29]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n877 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2569 (
    .a(\u2_Display/n841 ),
    .b(\u2_Display/n874 [30]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n876 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2570 (
    .a(\u2_Display/n840 ),
    .b(\u2_Display/n874 [31]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n875 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2571 (
    .a(\u2_Display/n1994 ),
    .b(\u2_Display/n1997 [0]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2029 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2572 (
    .a(\u2_Display/n1993 ),
    .b(\u2_Display/n1997 [1]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2028 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2573 (
    .a(\u2_Display/n1992 ),
    .b(\u2_Display/n1997 [2]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2027 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2574 (
    .a(\u2_Display/n1991 ),
    .b(\u2_Display/n1997 [3]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2026 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2575 (
    .a(\u2_Display/n1990 ),
    .b(\u2_Display/n1997 [4]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2025 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2576 (
    .a(\u2_Display/n1989 ),
    .b(\u2_Display/n1997 [5]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2024 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2577 (
    .a(\u2_Display/n1988 ),
    .b(\u2_Display/n1997 [6]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2023 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2578 (
    .a(\u2_Display/n1987 ),
    .b(\u2_Display/n1997 [7]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2022 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2579 (
    .a(\u2_Display/n1986 ),
    .b(\u2_Display/n1997 [8]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2021 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2580 (
    .a(\u2_Display/n1985 ),
    .b(\u2_Display/n1997 [9]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2020 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2581 (
    .a(\u2_Display/n1984 ),
    .b(\u2_Display/n1997 [10]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2019 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2582 (
    .a(\u2_Display/n1983 ),
    .b(\u2_Display/n1997 [11]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2018 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2583 (
    .a(\u2_Display/n1982 ),
    .b(\u2_Display/n1997 [12]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2017 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2584 (
    .a(\u2_Display/n1981 ),
    .b(\u2_Display/n1997 [13]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2016 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2585 (
    .a(\u2_Display/n1980 ),
    .b(\u2_Display/n1997 [14]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2015 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2586 (
    .a(\u2_Display/n1979 ),
    .b(\u2_Display/n1997 [15]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2014 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2587 (
    .a(\u2_Display/n1978 ),
    .b(\u2_Display/n1997 [16]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2013 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2588 (
    .a(\u2_Display/n1977 ),
    .b(\u2_Display/n1997 [17]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2012 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2589 (
    .a(\u2_Display/n1976 ),
    .b(\u2_Display/n1997 [18]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2011 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2590 (
    .a(\u2_Display/n1975 ),
    .b(\u2_Display/n1997 [19]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2010 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2591 (
    .a(\u2_Display/n1974 ),
    .b(\u2_Display/n1997 [20]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2009 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2592 (
    .a(\u2_Display/n1973 ),
    .b(\u2_Display/n1997 [21]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2008 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2593 (
    .a(\u2_Display/n1972 ),
    .b(\u2_Display/n1997 [22]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2007 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2594 (
    .a(\u2_Display/n1971 ),
    .b(\u2_Display/n1997 [23]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2006 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2595 (
    .a(\u2_Display/n1970 ),
    .b(\u2_Display/n1997 [24]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2005 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2596 (
    .a(\u2_Display/n1969 ),
    .b(\u2_Display/n1997 [25]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2004 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2597 (
    .a(\u2_Display/n1968 ),
    .b(\u2_Display/n1997 [26]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2003 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2598 (
    .a(\u2_Display/n1967 ),
    .b(\u2_Display/n1997 [27]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2002 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2599 (
    .a(\u2_Display/n1966 ),
    .b(\u2_Display/n1997 [28]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2001 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2600 (
    .a(\u2_Display/n1965 ),
    .b(\u2_Display/n1997 [29]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2000 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2601 (
    .a(\u2_Display/n1964 ),
    .b(\u2_Display/n1997 [30]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n1999 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2602 (
    .a(\u2_Display/n1963 ),
    .b(\u2_Display/n1997 [31]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n1998 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2603 (
    .a(\u2_Display/n3117 ),
    .b(\u2_Display/n3120 [0]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3152 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2604 (
    .a(\u2_Display/n3116 ),
    .b(\u2_Display/n3120 [1]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3151 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2605 (
    .a(\u2_Display/n3115 ),
    .b(\u2_Display/n3120 [2]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3150 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2606 (
    .a(\u2_Display/n3114 ),
    .b(\u2_Display/n3120 [3]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3149 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2607 (
    .a(\u2_Display/n3113 ),
    .b(\u2_Display/n3120 [4]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3148 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2608 (
    .a(\u2_Display/n3112 ),
    .b(\u2_Display/n3120 [5]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3147 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2609 (
    .a(\u2_Display/n3111 ),
    .b(\u2_Display/n3120 [6]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3146 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2610 (
    .a(\u2_Display/n3110 ),
    .b(\u2_Display/n3120 [7]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3145 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2611 (
    .a(\u2_Display/n3109 ),
    .b(\u2_Display/n3120 [8]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3144 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2612 (
    .a(\u2_Display/n3108 ),
    .b(\u2_Display/n3120 [9]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3143 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2613 (
    .a(\u2_Display/n3107 ),
    .b(\u2_Display/n3120 [10]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3142 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2614 (
    .a(\u2_Display/n3106 ),
    .b(\u2_Display/n3120 [11]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3141 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2615 (
    .a(\u2_Display/n3105 ),
    .b(\u2_Display/n3120 [12]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3140 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2616 (
    .a(\u2_Display/n3104 ),
    .b(\u2_Display/n3120 [13]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3139 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2617 (
    .a(\u2_Display/n3103 ),
    .b(\u2_Display/n3120 [14]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3138 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2618 (
    .a(\u2_Display/n3102 ),
    .b(\u2_Display/n3120 [15]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3137 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2619 (
    .a(\u2_Display/n3101 ),
    .b(\u2_Display/n3120 [16]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3136 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2620 (
    .a(\u2_Display/n3100 ),
    .b(\u2_Display/n3120 [17]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3135 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2621 (
    .a(\u2_Display/n3099 ),
    .b(\u2_Display/n3120 [18]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3134 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2622 (
    .a(\u2_Display/n3098 ),
    .b(\u2_Display/n3120 [19]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3133 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2623 (
    .a(\u2_Display/n3097 ),
    .b(\u2_Display/n3120 [20]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3132 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2624 (
    .a(\u2_Display/n3096 ),
    .b(\u2_Display/n3120 [21]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3131 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2625 (
    .a(\u2_Display/n3095 ),
    .b(\u2_Display/n3120 [22]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3130 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2626 (
    .a(\u2_Display/n3094 ),
    .b(\u2_Display/n3120 [23]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3129 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2627 (
    .a(\u2_Display/n3093 ),
    .b(\u2_Display/n3120 [24]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3128 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2628 (
    .a(\u2_Display/n3092 ),
    .b(\u2_Display/n3120 [25]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3127 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2629 (
    .a(\u2_Display/n3091 ),
    .b(\u2_Display/n3120 [26]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3126 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2630 (
    .a(\u2_Display/n3090 ),
    .b(\u2_Display/n3120 [27]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3125 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2631 (
    .a(\u2_Display/n3089 ),
    .b(\u2_Display/n3120 [28]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3124 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2632 (
    .a(\u2_Display/n3088 ),
    .b(\u2_Display/n3120 [29]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3123 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2633 (
    .a(\u2_Display/n3087 ),
    .b(\u2_Display/n3120 [30]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3122 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2634 (
    .a(\u2_Display/n3086 ),
    .b(\u2_Display/n3120 [31]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3121 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2635 (
    .a(\u2_Display/n4275 ),
    .b(\u2_Display/n4278 [0]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4310 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2636 (
    .a(\u2_Display/n4274 ),
    .b(\u2_Display/n4278 [1]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4309 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2637 (
    .a(\u2_Display/n4273 ),
    .b(\u2_Display/n4278 [2]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4308 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2638 (
    .a(\u2_Display/n4272 ),
    .b(\u2_Display/n4278 [3]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4307 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2639 (
    .a(\u2_Display/n4271 ),
    .b(\u2_Display/n4278 [4]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4306 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2640 (
    .a(\u2_Display/n4270 ),
    .b(\u2_Display/n4278 [5]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4305 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2641 (
    .a(\u2_Display/n4269 ),
    .b(\u2_Display/n4278 [6]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4304 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2642 (
    .a(\u2_Display/n4268 ),
    .b(\u2_Display/n4278 [7]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4303 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2643 (
    .a(\u2_Display/n4267 ),
    .b(\u2_Display/n4278 [8]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4302 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2644 (
    .a(\u2_Display/n4266 ),
    .b(\u2_Display/n4278 [9]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4301 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2645 (
    .a(\u2_Display/n4265 ),
    .b(\u2_Display/n4278 [10]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4300 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2646 (
    .a(\u2_Display/n4264 ),
    .b(\u2_Display/n4278 [11]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4299 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2647 (
    .a(\u2_Display/n4263 ),
    .b(\u2_Display/n4278 [12]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4298 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2648 (
    .a(\u2_Display/n4262 ),
    .b(\u2_Display/n4278 [13]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4297 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2649 (
    .a(\u2_Display/n4261 ),
    .b(\u2_Display/n4278 [14]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4296 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2650 (
    .a(\u2_Display/n4260 ),
    .b(\u2_Display/n4278 [15]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4295 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2651 (
    .a(\u2_Display/n4259 ),
    .b(\u2_Display/n4278 [16]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4294 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2652 (
    .a(\u2_Display/n4258 ),
    .b(\u2_Display/n4278 [17]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4293 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2653 (
    .a(\u2_Display/n4257 ),
    .b(\u2_Display/n4278 [18]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4292 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2654 (
    .a(\u2_Display/n4256 ),
    .b(\u2_Display/n4278 [19]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4291 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2655 (
    .a(\u2_Display/n4255 ),
    .b(\u2_Display/n4278 [20]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4290 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2656 (
    .a(\u2_Display/n4254 ),
    .b(\u2_Display/n4278 [21]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4289 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2657 (
    .a(\u2_Display/n4253 ),
    .b(\u2_Display/n4278 [22]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4288 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2658 (
    .a(\u2_Display/n4252 ),
    .b(\u2_Display/n4278 [23]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4287 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2659 (
    .a(\u2_Display/n4251 ),
    .b(\u2_Display/n4278 [24]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4286 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2660 (
    .a(\u2_Display/n4250 ),
    .b(\u2_Display/n4278 [25]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4285 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2661 (
    .a(\u2_Display/n4249 ),
    .b(\u2_Display/n4278 [26]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4284 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2662 (
    .a(\u2_Display/n4248 ),
    .b(\u2_Display/n4278 [27]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4283 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2663 (
    .a(\u2_Display/n4247 ),
    .b(\u2_Display/n4278 [28]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4282 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2664 (
    .a(\u2_Display/n4246 ),
    .b(\u2_Display/n4278 [29]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4281 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2665 (
    .a(\u2_Display/n4245 ),
    .b(\u2_Display/n4278 [30]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4280 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2666 (
    .a(\u2_Display/n4244 ),
    .b(\u2_Display/n4278 [31]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4279 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2667 (
    .a(\u2_Display/n5398 ),
    .b(\u2_Display/n5401 [0]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5433 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2668 (
    .a(\u2_Display/n5397 ),
    .b(\u2_Display/n5401 [1]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5432 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2669 (
    .a(\u2_Display/n5396 ),
    .b(\u2_Display/n5401 [2]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5431 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2670 (
    .a(\u2_Display/n5395 ),
    .b(\u2_Display/n5401 [3]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5430 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2671 (
    .a(\u2_Display/n5394 ),
    .b(\u2_Display/n5401 [4]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5429 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2672 (
    .a(\u2_Display/n5393 ),
    .b(\u2_Display/n5401 [5]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5428 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2673 (
    .a(\u2_Display/n5392 ),
    .b(\u2_Display/n5401 [6]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5427 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2674 (
    .a(\u2_Display/n5391 ),
    .b(\u2_Display/n5401 [7]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5426 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2675 (
    .a(\u2_Display/n5390 ),
    .b(\u2_Display/n5401 [8]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5425 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2676 (
    .a(\u2_Display/n5389 ),
    .b(\u2_Display/n5401 [9]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5424 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2677 (
    .a(\u2_Display/n5388 ),
    .b(\u2_Display/n5401 [10]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5423 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2678 (
    .a(\u2_Display/n5387 ),
    .b(\u2_Display/n5401 [11]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5422 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2679 (
    .a(\u2_Display/n5386 ),
    .b(\u2_Display/n5401 [12]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5421 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2680 (
    .a(\u2_Display/n5385 ),
    .b(\u2_Display/n5401 [13]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5420 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2681 (
    .a(\u2_Display/n5384 ),
    .b(\u2_Display/n5401 [14]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5419 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2682 (
    .a(\u2_Display/n5383 ),
    .b(\u2_Display/n5401 [15]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5418 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2683 (
    .a(\u2_Display/n5382 ),
    .b(\u2_Display/n5401 [16]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5417 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2684 (
    .a(\u2_Display/n5381 ),
    .b(\u2_Display/n5401 [17]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5416 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2685 (
    .a(\u2_Display/n5380 ),
    .b(\u2_Display/n5401 [18]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5415 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2686 (
    .a(\u2_Display/n5379 ),
    .b(\u2_Display/n5401 [19]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5414 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2687 (
    .a(\u2_Display/n5378 ),
    .b(\u2_Display/n5401 [20]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5413 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2688 (
    .a(\u2_Display/n5377 ),
    .b(\u2_Display/n5401 [21]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5412 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2689 (
    .a(\u2_Display/n5376 ),
    .b(\u2_Display/n5401 [22]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5411 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2690 (
    .a(\u2_Display/n5375 ),
    .b(\u2_Display/n5401 [23]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5410 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2691 (
    .a(\u2_Display/n5374 ),
    .b(\u2_Display/n5401 [24]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5409 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2692 (
    .a(\u2_Display/n5373 ),
    .b(\u2_Display/n5401 [25]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5408 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2693 (
    .a(\u2_Display/n5372 ),
    .b(\u2_Display/n5401 [26]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5407 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2694 (
    .a(\u2_Display/n5371 ),
    .b(\u2_Display/n5401 [27]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5406 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2695 (
    .a(\u2_Display/n5370 ),
    .b(\u2_Display/n5401 [28]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5405 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2696 (
    .a(\u2_Display/n5369 ),
    .b(\u2_Display/n5401 [29]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5404 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2697 (
    .a(\u2_Display/n5368 ),
    .b(\u2_Display/n5401 [30]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5403 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2698 (
    .a(\u2_Display/n5367 ),
    .b(\u2_Display/n5401 [31]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5402 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2699 (
    .a(\u2_Display/n906 ),
    .b(\u2_Display/n909 [0]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n941 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2700 (
    .a(\u2_Display/n905 ),
    .b(\u2_Display/n909 [1]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n940 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2701 (
    .a(\u2_Display/n904 ),
    .b(\u2_Display/n909 [2]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n939 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2702 (
    .a(\u2_Display/n903 ),
    .b(\u2_Display/n909 [3]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n938 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2703 (
    .a(\u2_Display/n902 ),
    .b(\u2_Display/n909 [4]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n937 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2704 (
    .a(\u2_Display/n901 ),
    .b(\u2_Display/n909 [5]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n936 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2705 (
    .a(\u2_Display/n900 ),
    .b(\u2_Display/n909 [6]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n935 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2706 (
    .a(\u2_Display/n899 ),
    .b(\u2_Display/n909 [7]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n934 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2707 (
    .a(\u2_Display/n898 ),
    .b(\u2_Display/n909 [8]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n933 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2708 (
    .a(\u2_Display/n897 ),
    .b(\u2_Display/n909 [9]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n932 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2709 (
    .a(\u2_Display/n896 ),
    .b(\u2_Display/n909 [10]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n931 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2710 (
    .a(\u2_Display/n895 ),
    .b(\u2_Display/n909 [11]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n930 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2711 (
    .a(\u2_Display/n894 ),
    .b(\u2_Display/n909 [12]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n929 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2712 (
    .a(\u2_Display/n893 ),
    .b(\u2_Display/n909 [13]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n928 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2713 (
    .a(\u2_Display/n892 ),
    .b(\u2_Display/n909 [14]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n927 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2714 (
    .a(\u2_Display/n891 ),
    .b(\u2_Display/n909 [15]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n926 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2715 (
    .a(\u2_Display/n890 ),
    .b(\u2_Display/n909 [16]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n925 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2716 (
    .a(\u2_Display/n889 ),
    .b(\u2_Display/n909 [17]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n924 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2717 (
    .a(\u2_Display/n888 ),
    .b(\u2_Display/n909 [18]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n923 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2718 (
    .a(\u2_Display/n887 ),
    .b(\u2_Display/n909 [19]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n922 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2719 (
    .a(\u2_Display/n886 ),
    .b(\u2_Display/n909 [20]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n921 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2720 (
    .a(\u2_Display/n885 ),
    .b(\u2_Display/n909 [21]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n920 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2721 (
    .a(\u2_Display/n884 ),
    .b(\u2_Display/n909 [22]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n919 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2722 (
    .a(\u2_Display/n883 ),
    .b(\u2_Display/n909 [23]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n918 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2723 (
    .a(\u2_Display/n882 ),
    .b(\u2_Display/n909 [24]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n917 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2724 (
    .a(\u2_Display/n881 ),
    .b(\u2_Display/n909 [25]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n916 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2725 (
    .a(\u2_Display/n880 ),
    .b(\u2_Display/n909 [26]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n915 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2726 (
    .a(\u2_Display/n879 ),
    .b(\u2_Display/n909 [27]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n914 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2727 (
    .a(\u2_Display/n878 ),
    .b(\u2_Display/n909 [28]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n913 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2728 (
    .a(\u2_Display/n877 ),
    .b(\u2_Display/n909 [29]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n912 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2729 (
    .a(\u2_Display/n876 ),
    .b(\u2_Display/n909 [30]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n911 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2730 (
    .a(\u2_Display/n875 ),
    .b(\u2_Display/n909 [31]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n910 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2731 (
    .a(\u2_Display/n2029 ),
    .b(\u2_Display/n2032 [0]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2064 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2732 (
    .a(\u2_Display/n2028 ),
    .b(\u2_Display/n2032 [1]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2063 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2733 (
    .a(\u2_Display/n2027 ),
    .b(\u2_Display/n2032 [2]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2062 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2734 (
    .a(\u2_Display/n2026 ),
    .b(\u2_Display/n2032 [3]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2061 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2735 (
    .a(\u2_Display/n2025 ),
    .b(\u2_Display/n2032 [4]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2060 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2736 (
    .a(\u2_Display/n2024 ),
    .b(\u2_Display/n2032 [5]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2059 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2737 (
    .a(\u2_Display/n2023 ),
    .b(\u2_Display/n2032 [6]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2058 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2738 (
    .a(\u2_Display/n2022 ),
    .b(\u2_Display/n2032 [7]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2057 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2739 (
    .a(\u2_Display/n2021 ),
    .b(\u2_Display/n2032 [8]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2056 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2740 (
    .a(\u2_Display/n2020 ),
    .b(\u2_Display/n2032 [9]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2055 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2741 (
    .a(\u2_Display/n2019 ),
    .b(\u2_Display/n2032 [10]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2054 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2742 (
    .a(\u2_Display/n2018 ),
    .b(\u2_Display/n2032 [11]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2053 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2743 (
    .a(\u2_Display/n2017 ),
    .b(\u2_Display/n2032 [12]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2052 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2744 (
    .a(\u2_Display/n2016 ),
    .b(\u2_Display/n2032 [13]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2051 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2745 (
    .a(\u2_Display/n2015 ),
    .b(\u2_Display/n2032 [14]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2050 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2746 (
    .a(\u2_Display/n2014 ),
    .b(\u2_Display/n2032 [15]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2049 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2747 (
    .a(\u2_Display/n2013 ),
    .b(\u2_Display/n2032 [16]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2048 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2748 (
    .a(\u2_Display/n2012 ),
    .b(\u2_Display/n2032 [17]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2047 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2749 (
    .a(\u2_Display/n2011 ),
    .b(\u2_Display/n2032 [18]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2046 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2750 (
    .a(\u2_Display/n2010 ),
    .b(\u2_Display/n2032 [19]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2045 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2751 (
    .a(\u2_Display/n2009 ),
    .b(\u2_Display/n2032 [20]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2044 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2752 (
    .a(\u2_Display/n2008 ),
    .b(\u2_Display/n2032 [21]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2043 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2753 (
    .a(\u2_Display/n2007 ),
    .b(\u2_Display/n2032 [22]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2042 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2754 (
    .a(\u2_Display/n2006 ),
    .b(\u2_Display/n2032 [23]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2041 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2755 (
    .a(\u2_Display/n2005 ),
    .b(\u2_Display/n2032 [24]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2040 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2756 (
    .a(\u2_Display/n2004 ),
    .b(\u2_Display/n2032 [25]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2039 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2757 (
    .a(\u2_Display/n2003 ),
    .b(\u2_Display/n2032 [26]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2038 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2758 (
    .a(\u2_Display/n2002 ),
    .b(\u2_Display/n2032 [27]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2037 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2759 (
    .a(\u2_Display/n2001 ),
    .b(\u2_Display/n2032 [28]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2036 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2760 (
    .a(\u2_Display/n2000 ),
    .b(\u2_Display/n2032 [29]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2035 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2761 (
    .a(\u2_Display/n1999 ),
    .b(\u2_Display/n2032 [30]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2034 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2762 (
    .a(\u2_Display/n1998 ),
    .b(\u2_Display/n2032 [31]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2033 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2763 (
    .a(\u2_Display/n3152 ),
    .b(\u2_Display/n3155 [0]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3187 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2764 (
    .a(\u2_Display/n3151 ),
    .b(\u2_Display/n3155 [1]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3186 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2765 (
    .a(\u2_Display/n3150 ),
    .b(\u2_Display/n3155 [2]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3185 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2766 (
    .a(\u2_Display/n3149 ),
    .b(\u2_Display/n3155 [3]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3184 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2767 (
    .a(\u2_Display/n3148 ),
    .b(\u2_Display/n3155 [4]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3183 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2768 (
    .a(\u2_Display/n3147 ),
    .b(\u2_Display/n3155 [5]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3182 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2769 (
    .a(\u2_Display/n3146 ),
    .b(\u2_Display/n3155 [6]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3181 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2770 (
    .a(\u2_Display/n3145 ),
    .b(\u2_Display/n3155 [7]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3180 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2771 (
    .a(\u2_Display/n3144 ),
    .b(\u2_Display/n3155 [8]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3179 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2772 (
    .a(\u2_Display/n3143 ),
    .b(\u2_Display/n3155 [9]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3178 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2773 (
    .a(\u2_Display/n3142 ),
    .b(\u2_Display/n3155 [10]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3177 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2774 (
    .a(\u2_Display/n3141 ),
    .b(\u2_Display/n3155 [11]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3176 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2775 (
    .a(\u2_Display/n3140 ),
    .b(\u2_Display/n3155 [12]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3175 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2776 (
    .a(\u2_Display/n3139 ),
    .b(\u2_Display/n3155 [13]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3174 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2777 (
    .a(\u2_Display/n3138 ),
    .b(\u2_Display/n3155 [14]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3173 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2778 (
    .a(\u2_Display/n3137 ),
    .b(\u2_Display/n3155 [15]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3172 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2779 (
    .a(\u2_Display/n3136 ),
    .b(\u2_Display/n3155 [16]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3171 ));
  EG_PHY_PAD #(
    //.LOCATION("K14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u278 (
    .ipad(clk_24m),
    .di(clk_24m_pad));  // source/rtl/VGA_Demo.v(4)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2780 (
    .a(\u2_Display/n3135 ),
    .b(\u2_Display/n3155 [17]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3170 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2781 (
    .a(\u2_Display/n3134 ),
    .b(\u2_Display/n3155 [18]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3169 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2782 (
    .a(\u2_Display/n3133 ),
    .b(\u2_Display/n3155 [19]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3168 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2783 (
    .a(\u2_Display/n3132 ),
    .b(\u2_Display/n3155 [20]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3167 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2784 (
    .a(\u2_Display/n3131 ),
    .b(\u2_Display/n3155 [21]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3166 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2785 (
    .a(\u2_Display/n3130 ),
    .b(\u2_Display/n3155 [22]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3165 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2786 (
    .a(\u2_Display/n3129 ),
    .b(\u2_Display/n3155 [23]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3164 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2787 (
    .a(\u2_Display/n3128 ),
    .b(\u2_Display/n3155 [24]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3163 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2788 (
    .a(\u2_Display/n3127 ),
    .b(\u2_Display/n3155 [25]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3162 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2789 (
    .a(\u2_Display/n3126 ),
    .b(\u2_Display/n3155 [26]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3161 ));
  EG_PHY_PAD #(
    //.LOCATION("P8"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u279 (
    .ipad(on_off[7]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2790 (
    .a(\u2_Display/n3125 ),
    .b(\u2_Display/n3155 [27]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3160 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2791 (
    .a(\u2_Display/n3124 ),
    .b(\u2_Display/n3155 [28]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3159 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2792 (
    .a(\u2_Display/n3123 ),
    .b(\u2_Display/n3155 [29]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3158 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2793 (
    .a(\u2_Display/n3122 ),
    .b(\u2_Display/n3155 [30]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3157 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2794 (
    .a(\u2_Display/n3121 ),
    .b(\u2_Display/n3155 [31]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3156 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2795 (
    .a(\u2_Display/n4310 ),
    .b(\u2_Display/n4313 [0]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4345 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2796 (
    .a(\u2_Display/n4309 ),
    .b(\u2_Display/n4313 [1]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4344 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2797 (
    .a(\u2_Display/n4308 ),
    .b(\u2_Display/n4313 [2]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4343 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2798 (
    .a(\u2_Display/n4307 ),
    .b(\u2_Display/n4313 [3]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4342 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2799 (
    .a(\u2_Display/n4306 ),
    .b(\u2_Display/n4313 [4]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4341 ));
  EG_PHY_PAD #(
    //.LOCATION("N6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u280 (
    .ipad(on_off[6]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2800 (
    .a(\u2_Display/n4305 ),
    .b(\u2_Display/n4313 [5]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4340 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2801 (
    .a(\u2_Display/n4304 ),
    .b(\u2_Display/n4313 [6]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4339 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2802 (
    .a(\u2_Display/n4303 ),
    .b(\u2_Display/n4313 [7]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4338 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2803 (
    .a(\u2_Display/n4302 ),
    .b(\u2_Display/n4313 [8]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4337 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2804 (
    .a(\u2_Display/n4301 ),
    .b(\u2_Display/n4313 [9]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4336 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2805 (
    .a(\u2_Display/n4300 ),
    .b(\u2_Display/n4313 [10]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4335 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2806 (
    .a(\u2_Display/n4299 ),
    .b(\u2_Display/n4313 [11]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4334 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2807 (
    .a(\u2_Display/n4298 ),
    .b(\u2_Display/n4313 [12]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4333 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2808 (
    .a(\u2_Display/n4297 ),
    .b(\u2_Display/n4313 [13]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4332 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2809 (
    .a(\u2_Display/n4296 ),
    .b(\u2_Display/n4313 [14]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4331 ));
  EG_PHY_PAD #(
    //.LOCATION("P6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u281 (
    .ipad(on_off[5]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2810 (
    .a(\u2_Display/n4295 ),
    .b(\u2_Display/n4313 [15]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4330 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2811 (
    .a(\u2_Display/n4294 ),
    .b(\u2_Display/n4313 [16]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4329 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2812 (
    .a(\u2_Display/n4293 ),
    .b(\u2_Display/n4313 [17]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4328 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2813 (
    .a(\u2_Display/n4292 ),
    .b(\u2_Display/n4313 [18]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4327 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2814 (
    .a(\u2_Display/n4291 ),
    .b(\u2_Display/n4313 [19]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4326 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2815 (
    .a(\u2_Display/n4290 ),
    .b(\u2_Display/n4313 [20]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4325 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2816 (
    .a(\u2_Display/n4289 ),
    .b(\u2_Display/n4313 [21]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4324 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2817 (
    .a(\u2_Display/n4288 ),
    .b(\u2_Display/n4313 [22]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4323 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2818 (
    .a(\u2_Display/n4287 ),
    .b(\u2_Display/n4313 [23]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4322 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2819 (
    .a(\u2_Display/n4286 ),
    .b(\u2_Display/n4313 [24]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4321 ));
  EG_PHY_PAD #(
    //.LOCATION("M6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u282 (
    .ipad(on_off[4]),
    .di(on_off_pad[4]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2820 (
    .a(\u2_Display/n4285 ),
    .b(\u2_Display/n4313 [25]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4320 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2821 (
    .a(\u2_Display/n4284 ),
    .b(\u2_Display/n4313 [26]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4319 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2822 (
    .a(\u2_Display/n4283 ),
    .b(\u2_Display/n4313 [27]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4318 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2823 (
    .a(\u2_Display/n4282 ),
    .b(\u2_Display/n4313 [28]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4317 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2824 (
    .a(\u2_Display/n4281 ),
    .b(\u2_Display/n4313 [29]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4316 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2825 (
    .a(\u2_Display/n4280 ),
    .b(\u2_Display/n4313 [30]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4315 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2826 (
    .a(\u2_Display/n4279 ),
    .b(\u2_Display/n4313 [31]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4314 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2827 (
    .a(\u2_Display/n5433 ),
    .b(\u2_Display/n5436 [0]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5468 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2828 (
    .a(\u2_Display/n5432 ),
    .b(\u2_Display/n5436 [1]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5467 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2829 (
    .a(\u2_Display/n5431 ),
    .b(\u2_Display/n5436 [2]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5466 ));
  EG_PHY_PAD #(
    //.LOCATION("T6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u283 (
    .ipad(on_off[3]),
    .di(on_off_pad[3]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2830 (
    .a(\u2_Display/n5430 ),
    .b(\u2_Display/n5436 [3]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5465 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2831 (
    .a(\u2_Display/n5429 ),
    .b(\u2_Display/n5436 [4]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5464 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2832 (
    .a(\u2_Display/n5428 ),
    .b(\u2_Display/n5436 [5]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5463 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2833 (
    .a(\u2_Display/n5427 ),
    .b(\u2_Display/n5436 [6]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5462 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2834 (
    .a(\u2_Display/n5426 ),
    .b(\u2_Display/n5436 [7]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5461 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2835 (
    .a(\u2_Display/n5425 ),
    .b(\u2_Display/n5436 [8]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5460 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2836 (
    .a(\u2_Display/n5424 ),
    .b(\u2_Display/n5436 [9]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5459 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2837 (
    .a(\u2_Display/n5423 ),
    .b(\u2_Display/n5436 [10]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5458 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2838 (
    .a(\u2_Display/n5422 ),
    .b(\u2_Display/n5436 [11]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5457 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2839 (
    .a(\u2_Display/n5421 ),
    .b(\u2_Display/n5436 [12]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5456 ));
  EG_PHY_PAD #(
    //.LOCATION("T5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u284 (
    .ipad(on_off[2]),
    .di(on_off_pad[2]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2840 (
    .a(\u2_Display/n5420 ),
    .b(\u2_Display/n5436 [13]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5455 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2841 (
    .a(\u2_Display/n5419 ),
    .b(\u2_Display/n5436 [14]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5454 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2842 (
    .a(\u2_Display/n5418 ),
    .b(\u2_Display/n5436 [15]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5453 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2843 (
    .a(\u2_Display/n5417 ),
    .b(\u2_Display/n5436 [16]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5452 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2844 (
    .a(\u2_Display/n5416 ),
    .b(\u2_Display/n5436 [17]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5451 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2845 (
    .a(\u2_Display/n5415 ),
    .b(\u2_Display/n5436 [18]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5450 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2846 (
    .a(\u2_Display/n5414 ),
    .b(\u2_Display/n5436 [19]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5449 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2847 (
    .a(\u2_Display/n5413 ),
    .b(\u2_Display/n5436 [20]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5448 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2848 (
    .a(\u2_Display/n5412 ),
    .b(\u2_Display/n5436 [21]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5447 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2849 (
    .a(\u2_Display/n5411 ),
    .b(\u2_Display/n5436 [22]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5446 ));
  EG_PHY_PAD #(
    //.LOCATION("R5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u285 (
    .ipad(on_off[1]),
    .di(on_off_pad[1]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2850 (
    .a(\u2_Display/n5410 ),
    .b(\u2_Display/n5436 [23]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5445 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2851 (
    .a(\u2_Display/n5409 ),
    .b(\u2_Display/n5436 [24]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5444 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2852 (
    .a(\u2_Display/n5408 ),
    .b(\u2_Display/n5436 [25]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5443 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2853 (
    .a(\u2_Display/n5407 ),
    .b(\u2_Display/n5436 [26]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5442 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2854 (
    .a(\u2_Display/n5406 ),
    .b(\u2_Display/n5436 [27]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5441 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2855 (
    .a(\u2_Display/n5405 ),
    .b(\u2_Display/n5436 [28]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5440 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2856 (
    .a(\u2_Display/n5404 ),
    .b(\u2_Display/n5436 [29]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5439 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2857 (
    .a(\u2_Display/n5403 ),
    .b(\u2_Display/n5436 [30]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5438 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2858 (
    .a(\u2_Display/n5402 ),
    .b(\u2_Display/n5436 [31]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5437 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2859 (
    .a(\u2_Display/n941 ),
    .b(\u2_Display/n944 [0]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n976 ));
  EG_PHY_PAD #(
    //.LOCATION("T4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u286 (
    .ipad(on_off[0]),
    .di(on_off_pad[0]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2860 (
    .a(\u2_Display/n940 ),
    .b(\u2_Display/n944 [1]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n975 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2861 (
    .a(\u2_Display/n939 ),
    .b(\u2_Display/n944 [2]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n974 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2862 (
    .a(\u2_Display/n938 ),
    .b(\u2_Display/n944 [3]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n973 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2863 (
    .a(\u2_Display/n937 ),
    .b(\u2_Display/n944 [4]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n972 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2864 (
    .a(\u2_Display/n936 ),
    .b(\u2_Display/n944 [5]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n971 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2865 (
    .a(\u2_Display/n935 ),
    .b(\u2_Display/n944 [6]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n970 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2866 (
    .a(\u2_Display/n934 ),
    .b(\u2_Display/n944 [7]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n969 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2867 (
    .a(\u2_Display/n933 ),
    .b(\u2_Display/n944 [8]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n968 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2868 (
    .a(\u2_Display/n932 ),
    .b(\u2_Display/n944 [9]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n967 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2869 (
    .a(\u2_Display/n931 ),
    .b(\u2_Display/n944 [10]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n966 ));
  EG_PHY_PAD #(
    //.LOCATION("G11"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u287 (
    .ipad(rst_n),
    .di(rst_n_pad));  // source/rtl/VGA_Demo.v(5)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2870 (
    .a(\u2_Display/n930 ),
    .b(\u2_Display/n944 [11]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n965 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2871 (
    .a(\u2_Display/n929 ),
    .b(\u2_Display/n944 [12]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n964 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2872 (
    .a(\u2_Display/n928 ),
    .b(\u2_Display/n944 [13]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n963 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2873 (
    .a(\u2_Display/n927 ),
    .b(\u2_Display/n944 [14]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n962 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2874 (
    .a(\u2_Display/n926 ),
    .b(\u2_Display/n944 [15]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n961 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2875 (
    .a(\u2_Display/n925 ),
    .b(\u2_Display/n944 [16]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n960 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2876 (
    .a(\u2_Display/n924 ),
    .b(\u2_Display/n944 [17]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n959 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2877 (
    .a(\u2_Display/n923 ),
    .b(\u2_Display/n944 [18]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n958 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2878 (
    .a(\u2_Display/n922 ),
    .b(\u2_Display/n944 [19]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n957 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2879 (
    .a(\u2_Display/n921 ),
    .b(\u2_Display/n944 [20]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n956 ));
  EG_PHY_PAD #(
    //.LOCATION("C1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u288 (
    .do({open_n174,open_n175,open_n176,vga_b_pad[0]}),
    .opad(vga_b[7]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2880 (
    .a(\u2_Display/n920 ),
    .b(\u2_Display/n944 [21]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n955 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2881 (
    .a(\u2_Display/n919 ),
    .b(\u2_Display/n944 [22]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n954 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2882 (
    .a(\u2_Display/n918 ),
    .b(\u2_Display/n944 [23]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n953 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2883 (
    .a(\u2_Display/n917 ),
    .b(\u2_Display/n944 [24]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n952 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2884 (
    .a(\u2_Display/n916 ),
    .b(\u2_Display/n944 [25]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n951 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2885 (
    .a(\u2_Display/n915 ),
    .b(\u2_Display/n944 [26]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n950 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2886 (
    .a(\u2_Display/n914 ),
    .b(\u2_Display/n944 [27]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n949 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2887 (
    .a(\u2_Display/n913 ),
    .b(\u2_Display/n944 [28]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n948 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2888 (
    .a(\u2_Display/n912 ),
    .b(\u2_Display/n944 [29]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n947 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2889 (
    .a(\u2_Display/n911 ),
    .b(\u2_Display/n944 [30]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n946 ));
  EG_PHY_PAD #(
    //.LOCATION("D1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u289 (
    .do({open_n191,open_n192,open_n193,vga_b_pad[0]}),
    .opad(vga_b[6]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2890 (
    .a(\u2_Display/n910 ),
    .b(\u2_Display/n944 [31]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n945 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2891 (
    .a(\u2_Display/n2064 ),
    .b(\u2_Display/n2067 [0]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2099 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2892 (
    .a(\u2_Display/n2063 ),
    .b(\u2_Display/n2067 [1]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2098 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2893 (
    .a(\u2_Display/n2062 ),
    .b(\u2_Display/n2067 [2]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2097 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2894 (
    .a(\u2_Display/n2061 ),
    .b(\u2_Display/n2067 [3]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2096 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2895 (
    .a(\u2_Display/n2060 ),
    .b(\u2_Display/n2067 [4]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2095 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2896 (
    .a(\u2_Display/n2059 ),
    .b(\u2_Display/n2067 [5]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2094 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2897 (
    .a(\u2_Display/n2058 ),
    .b(\u2_Display/n2067 [6]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2093 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2898 (
    .a(\u2_Display/n2057 ),
    .b(\u2_Display/n2067 [7]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2092 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2899 (
    .a(\u2_Display/n2056 ),
    .b(\u2_Display/n2067 [8]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2091 ));
  EG_PHY_PAD #(
    //.LOCATION("E2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u290 (
    .do({open_n208,open_n209,open_n210,vga_b_pad[0]}),
    .opad(vga_b[5]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2900 (
    .a(\u2_Display/n2055 ),
    .b(\u2_Display/n2067 [9]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2090 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2901 (
    .a(\u2_Display/n2054 ),
    .b(\u2_Display/n2067 [10]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2089 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2902 (
    .a(\u2_Display/n2053 ),
    .b(\u2_Display/n2067 [11]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2088 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2903 (
    .a(\u2_Display/n2052 ),
    .b(\u2_Display/n2067 [12]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2087 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2904 (
    .a(\u2_Display/n2051 ),
    .b(\u2_Display/n2067 [13]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2086 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2905 (
    .a(\u2_Display/n2050 ),
    .b(\u2_Display/n2067 [14]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2085 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2906 (
    .a(\u2_Display/n2049 ),
    .b(\u2_Display/n2067 [15]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2084 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2907 (
    .a(\u2_Display/n2048 ),
    .b(\u2_Display/n2067 [16]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2083 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2908 (
    .a(\u2_Display/n2047 ),
    .b(\u2_Display/n2067 [17]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2082 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2909 (
    .a(\u2_Display/n2046 ),
    .b(\u2_Display/n2067 [18]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2081 ));
  EG_PHY_PAD #(
    //.LOCATION("G3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u291 (
    .do({open_n225,open_n226,open_n227,vga_b_pad[0]}),
    .opad(vga_b[4]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2910 (
    .a(\u2_Display/n2045 ),
    .b(\u2_Display/n2067 [19]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2080 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2911 (
    .a(\u2_Display/n2044 ),
    .b(\u2_Display/n2067 [20]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2079 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2912 (
    .a(\u2_Display/n2043 ),
    .b(\u2_Display/n2067 [21]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2078 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2913 (
    .a(\u2_Display/n2042 ),
    .b(\u2_Display/n2067 [22]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2077 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2914 (
    .a(\u2_Display/n2041 ),
    .b(\u2_Display/n2067 [23]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2076 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2915 (
    .a(\u2_Display/n2040 ),
    .b(\u2_Display/n2067 [24]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2075 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2916 (
    .a(\u2_Display/n2039 ),
    .b(\u2_Display/n2067 [25]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2074 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2917 (
    .a(\u2_Display/n2038 ),
    .b(\u2_Display/n2067 [26]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2073 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2918 (
    .a(\u2_Display/n2037 ),
    .b(\u2_Display/n2067 [27]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2072 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2919 (
    .a(\u2_Display/n2036 ),
    .b(\u2_Display/n2067 [28]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2071 ));
  EG_PHY_PAD #(
    //.LOCATION("E1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u292 (
    .do({open_n242,open_n243,open_n244,vga_b_pad[0]}),
    .opad(vga_b[3]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2920 (
    .a(\u2_Display/n2035 ),
    .b(\u2_Display/n2067 [29]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2070 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2921 (
    .a(\u2_Display/n2034 ),
    .b(\u2_Display/n2067 [30]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2069 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2922 (
    .a(\u2_Display/n2033 ),
    .b(\u2_Display/n2067 [31]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2068 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2923 (
    .a(\u2_Display/n3187 ),
    .b(\u2_Display/n3190 [0]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3222 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2924 (
    .a(\u2_Display/n3186 ),
    .b(\u2_Display/n3190 [1]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3221 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2925 (
    .a(\u2_Display/n3185 ),
    .b(\u2_Display/n3190 [2]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3220 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2926 (
    .a(\u2_Display/n3184 ),
    .b(\u2_Display/n3190 [3]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3219 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2927 (
    .a(\u2_Display/n3183 ),
    .b(\u2_Display/n3190 [4]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3218 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2928 (
    .a(\u2_Display/n3182 ),
    .b(\u2_Display/n3190 [5]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3217 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2929 (
    .a(\u2_Display/n3181 ),
    .b(\u2_Display/n3190 [6]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3216 ));
  EG_PHY_PAD #(
    //.LOCATION("F2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u293 (
    .do({open_n259,open_n260,open_n261,vga_b_pad[0]}),
    .opad(vga_b[2]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2930 (
    .a(\u2_Display/n3180 ),
    .b(\u2_Display/n3190 [7]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3215 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2931 (
    .a(\u2_Display/n3179 ),
    .b(\u2_Display/n3190 [8]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3214 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2932 (
    .a(\u2_Display/n3178 ),
    .b(\u2_Display/n3190 [9]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3213 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2933 (
    .a(\u2_Display/n3177 ),
    .b(\u2_Display/n3190 [10]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3212 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2934 (
    .a(\u2_Display/n3176 ),
    .b(\u2_Display/n3190 [11]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3211 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2935 (
    .a(\u2_Display/n3175 ),
    .b(\u2_Display/n3190 [12]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3210 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2936 (
    .a(\u2_Display/n3174 ),
    .b(\u2_Display/n3190 [13]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3209 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2937 (
    .a(\u2_Display/n3173 ),
    .b(\u2_Display/n3190 [14]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3208 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2938 (
    .a(\u2_Display/n3172 ),
    .b(\u2_Display/n3190 [15]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3207 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2939 (
    .a(\u2_Display/n3171 ),
    .b(\u2_Display/n3190 [16]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3206 ));
  EG_PHY_PAD #(
    //.LOCATION("F1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u294 (
    .do({open_n276,open_n277,open_n278,vga_b_pad[0]}),
    .opad(vga_b[1]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2940 (
    .a(\u2_Display/n3170 ),
    .b(\u2_Display/n3190 [17]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3205 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2941 (
    .a(\u2_Display/n3169 ),
    .b(\u2_Display/n3190 [18]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3204 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2942 (
    .a(\u2_Display/n3168 ),
    .b(\u2_Display/n3190 [19]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3203 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2943 (
    .a(\u2_Display/n3167 ),
    .b(\u2_Display/n3190 [20]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3202 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2944 (
    .a(\u2_Display/n3166 ),
    .b(\u2_Display/n3190 [21]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3201 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2945 (
    .a(\u2_Display/n3165 ),
    .b(\u2_Display/n3190 [22]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3200 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2946 (
    .a(\u2_Display/n3164 ),
    .b(\u2_Display/n3190 [23]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3199 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2947 (
    .a(\u2_Display/n3163 ),
    .b(\u2_Display/n3190 [24]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3198 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2948 (
    .a(\u2_Display/n3162 ),
    .b(\u2_Display/n3190 [25]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3197 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2949 (
    .a(\u2_Display/n3161 ),
    .b(\u2_Display/n3190 [26]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3196 ));
  EG_PHY_PAD #(
    //.LOCATION("G1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u295 (
    .do({open_n293,open_n294,open_n295,vga_b_pad[0]}),
    .opad(vga_b[0]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2950 (
    .a(\u2_Display/n3160 ),
    .b(\u2_Display/n3190 [27]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3195 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2951 (
    .a(\u2_Display/n3159 ),
    .b(\u2_Display/n3190 [28]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3194 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2952 (
    .a(\u2_Display/n3158 ),
    .b(\u2_Display/n3190 [29]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3193 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2953 (
    .a(\u2_Display/n3157 ),
    .b(\u2_Display/n3190 [30]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3192 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2954 (
    .a(\u2_Display/n3156 ),
    .b(\u2_Display/n3190 [31]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3191 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2955 (
    .a(\u2_Display/n4345 ),
    .b(\u2_Display/n4348 [0]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4380 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2956 (
    .a(\u2_Display/n4344 ),
    .b(\u2_Display/n4348 [1]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4379 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2957 (
    .a(\u2_Display/n4343 ),
    .b(\u2_Display/n4348 [2]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4378 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2958 (
    .a(\u2_Display/n4342 ),
    .b(\u2_Display/n4348 [3]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4377 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2959 (
    .a(\u2_Display/n4341 ),
    .b(\u2_Display/n4348 [4]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4376 ));
  EG_PHY_PAD #(
    //.LOCATION("H2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u296 (
    .do({open_n310,open_n311,open_n312,vga_clk_pad}),
    .opad(vga_clk));  // source/rtl/VGA_Demo.v(9)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2960 (
    .a(\u2_Display/n4340 ),
    .b(\u2_Display/n4348 [5]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4375 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2961 (
    .a(\u2_Display/n4339 ),
    .b(\u2_Display/n4348 [6]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4374 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2962 (
    .a(\u2_Display/n4338 ),
    .b(\u2_Display/n4348 [7]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4373 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2963 (
    .a(\u2_Display/n4337 ),
    .b(\u2_Display/n4348 [8]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4372 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2964 (
    .a(\u2_Display/n4336 ),
    .b(\u2_Display/n4348 [9]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4371 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2965 (
    .a(\u2_Display/n4335 ),
    .b(\u2_Display/n4348 [10]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4370 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2966 (
    .a(\u2_Display/n4334 ),
    .b(\u2_Display/n4348 [11]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4369 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2967 (
    .a(\u2_Display/n4333 ),
    .b(\u2_Display/n4348 [12]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4368 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2968 (
    .a(\u2_Display/n4332 ),
    .b(\u2_Display/n4348 [13]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4367 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2969 (
    .a(\u2_Display/n4331 ),
    .b(\u2_Display/n4348 [14]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4366 ));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u297 (
    .do({open_n327,open_n328,open_n329,vga_de_pad}),
    .opad(vga_de));  // source/rtl/VGA_Demo.v(13)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2970 (
    .a(\u2_Display/n4330 ),
    .b(\u2_Display/n4348 [15]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4365 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2971 (
    .a(\u2_Display/n4329 ),
    .b(\u2_Display/n4348 [16]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4364 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2972 (
    .a(\u2_Display/n4328 ),
    .b(\u2_Display/n4348 [17]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4363 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2973 (
    .a(\u2_Display/n4327 ),
    .b(\u2_Display/n4348 [18]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4362 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2974 (
    .a(\u2_Display/n4326 ),
    .b(\u2_Display/n4348 [19]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4361 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2975 (
    .a(\u2_Display/n4325 ),
    .b(\u2_Display/n4348 [20]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4360 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2976 (
    .a(\u2_Display/n4324 ),
    .b(\u2_Display/n4348 [21]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4359 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2977 (
    .a(\u2_Display/n4323 ),
    .b(\u2_Display/n4348 [22]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4358 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2978 (
    .a(\u2_Display/n4322 ),
    .b(\u2_Display/n4348 [23]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4357 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2979 (
    .a(\u2_Display/n4321 ),
    .b(\u2_Display/n4348 [24]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4356 ));
  EG_PHY_PAD #(
    //.LOCATION("H5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u298 (
    .do({open_n344,open_n345,open_n346,vga_b_pad[0]}),
    .opad(vga_g[7]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2980 (
    .a(\u2_Display/n4320 ),
    .b(\u2_Display/n4348 [25]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4355 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2981 (
    .a(\u2_Display/n4319 ),
    .b(\u2_Display/n4348 [26]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4354 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2982 (
    .a(\u2_Display/n4318 ),
    .b(\u2_Display/n4348 [27]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4353 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2983 (
    .a(\u2_Display/n4317 ),
    .b(\u2_Display/n4348 [28]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4352 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2984 (
    .a(\u2_Display/n4316 ),
    .b(\u2_Display/n4348 [29]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4351 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2985 (
    .a(\u2_Display/n4315 ),
    .b(\u2_Display/n4348 [30]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4350 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2986 (
    .a(\u2_Display/n4314 ),
    .b(\u2_Display/n4348 [31]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4349 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2987 (
    .a(\u2_Display/n5468 ),
    .b(\u2_Display/n5471 [0]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5503 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2988 (
    .a(\u2_Display/n5467 ),
    .b(\u2_Display/n5471 [1]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5502 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2989 (
    .a(\u2_Display/n5466 ),
    .b(\u2_Display/n5471 [2]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5501 ));
  EG_PHY_PAD #(
    //.LOCATION("H1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u299 (
    .do({open_n361,open_n362,open_n363,vga_b_pad[0]}),
    .opad(vga_g[6]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2990 (
    .a(\u2_Display/n5465 ),
    .b(\u2_Display/n5471 [3]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5500 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2991 (
    .a(\u2_Display/n5464 ),
    .b(\u2_Display/n5471 [4]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5499 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2992 (
    .a(\u2_Display/n5463 ),
    .b(\u2_Display/n5471 [5]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5498 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2993 (
    .a(\u2_Display/n5462 ),
    .b(\u2_Display/n5471 [6]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5497 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2994 (
    .a(\u2_Display/n5461 ),
    .b(\u2_Display/n5471 [7]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5496 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2995 (
    .a(\u2_Display/n5460 ),
    .b(\u2_Display/n5471 [8]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5495 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2996 (
    .a(\u2_Display/n5459 ),
    .b(\u2_Display/n5471 [9]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5494 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2997 (
    .a(\u2_Display/n5458 ),
    .b(\u2_Display/n5471 [10]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5493 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2998 (
    .a(\u2_Display/n5457 ),
    .b(\u2_Display/n5471 [11]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5492 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2999 (
    .a(\u2_Display/n5456 ),
    .b(\u2_Display/n5471 [12]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5491 ));
  EG_PHY_PAD #(
    //.LOCATION("J6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u300 (
    .do({open_n378,open_n379,open_n380,vga_b_pad[0]}),
    .opad(vga_g[5]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3000 (
    .a(\u2_Display/n5455 ),
    .b(\u2_Display/n5471 [13]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5490 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3001 (
    .a(\u2_Display/n5454 ),
    .b(\u2_Display/n5471 [14]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5489 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3002 (
    .a(\u2_Display/n5453 ),
    .b(\u2_Display/n5471 [15]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5488 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3003 (
    .a(\u2_Display/n5452 ),
    .b(\u2_Display/n5471 [16]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5487 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3004 (
    .a(\u2_Display/n5451 ),
    .b(\u2_Display/n5471 [17]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5486 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3005 (
    .a(\u2_Display/n5450 ),
    .b(\u2_Display/n5471 [18]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5485 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3006 (
    .a(\u2_Display/n5449 ),
    .b(\u2_Display/n5471 [19]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5484 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3007 (
    .a(\u2_Display/n5448 ),
    .b(\u2_Display/n5471 [20]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5483 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3008 (
    .a(\u2_Display/n5447 ),
    .b(\u2_Display/n5471 [21]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5482 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3009 (
    .a(\u2_Display/n5446 ),
    .b(\u2_Display/n5471 [22]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5481 ));
  EG_PHY_PAD #(
    //.LOCATION("H3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u301 (
    .do({open_n395,open_n396,open_n397,vga_b_pad[0]}),
    .opad(vga_g[4]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3010 (
    .a(\u2_Display/n5445 ),
    .b(\u2_Display/n5471 [23]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5480 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3011 (
    .a(\u2_Display/n5444 ),
    .b(\u2_Display/n5471 [24]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5479 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3012 (
    .a(\u2_Display/n5443 ),
    .b(\u2_Display/n5471 [25]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5478 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3013 (
    .a(\u2_Display/n5442 ),
    .b(\u2_Display/n5471 [26]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5477 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3014 (
    .a(\u2_Display/n5441 ),
    .b(\u2_Display/n5471 [27]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5476 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3015 (
    .a(\u2_Display/n5440 ),
    .b(\u2_Display/n5471 [28]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5475 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3016 (
    .a(\u2_Display/n5439 ),
    .b(\u2_Display/n5471 [29]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5474 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3017 (
    .a(\u2_Display/n5438 ),
    .b(\u2_Display/n5471 [30]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5473 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3018 (
    .a(\u2_Display/n5437 ),
    .b(\u2_Display/n5471 [31]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5472 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3019 (
    .a(\u2_Display/n976 ),
    .b(\u2_Display/n979 [0]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1011 ));
  EG_PHY_PAD #(
    //.LOCATION("J1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u302 (
    .do({open_n412,open_n413,open_n414,vga_b_pad[0]}),
    .opad(vga_g[3]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3020 (
    .a(\u2_Display/n975 ),
    .b(\u2_Display/n979 [1]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1010 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3021 (
    .a(\u2_Display/n974 ),
    .b(\u2_Display/n979 [2]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1009 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3022 (
    .a(\u2_Display/n973 ),
    .b(\u2_Display/n979 [3]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1008 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3023 (
    .a(\u2_Display/n972 ),
    .b(\u2_Display/n979 [4]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1007 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3024 (
    .a(\u2_Display/n971 ),
    .b(\u2_Display/n979 [5]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1006 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3025 (
    .a(\u2_Display/n970 ),
    .b(\u2_Display/n979 [6]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1005 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3026 (
    .a(\u2_Display/n969 ),
    .b(\u2_Display/n979 [7]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1004 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3027 (
    .a(\u2_Display/n968 ),
    .b(\u2_Display/n979 [8]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1003 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3028 (
    .a(\u2_Display/n967 ),
    .b(\u2_Display/n979 [9]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1002 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3029 (
    .a(\u2_Display/n966 ),
    .b(\u2_Display/n979 [10]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1001 ));
  EG_PHY_PAD #(
    //.LOCATION("K1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u303 (
    .do({open_n429,open_n430,open_n431,vga_b_pad[0]}),
    .opad(vga_g[2]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3030 (
    .a(\u2_Display/n965 ),
    .b(\u2_Display/n979 [11]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1000 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3031 (
    .a(\u2_Display/n964 ),
    .b(\u2_Display/n979 [12]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n999 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3032 (
    .a(\u2_Display/n963 ),
    .b(\u2_Display/n979 [13]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n998 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3033 (
    .a(\u2_Display/n962 ),
    .b(\u2_Display/n979 [14]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n997 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3034 (
    .a(\u2_Display/n961 ),
    .b(\u2_Display/n979 [15]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n996 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3035 (
    .a(\u2_Display/n960 ),
    .b(\u2_Display/n979 [16]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n995 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3036 (
    .a(\u2_Display/n959 ),
    .b(\u2_Display/n979 [17]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n994 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3037 (
    .a(\u2_Display/n958 ),
    .b(\u2_Display/n979 [18]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n993 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3038 (
    .a(\u2_Display/n957 ),
    .b(\u2_Display/n979 [19]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n992 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3039 (
    .a(\u2_Display/n956 ),
    .b(\u2_Display/n979 [20]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n991 ));
  EG_PHY_PAD #(
    //.LOCATION("K2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u304 (
    .do({open_n446,open_n447,open_n448,vga_b_pad[0]}),
    .opad(vga_g[1]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3040 (
    .a(\u2_Display/n955 ),
    .b(\u2_Display/n979 [21]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n990 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3041 (
    .a(\u2_Display/n954 ),
    .b(\u2_Display/n979 [22]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n989 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3042 (
    .a(\u2_Display/n953 ),
    .b(\u2_Display/n979 [23]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n988 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3043 (
    .a(\u2_Display/n952 ),
    .b(\u2_Display/n979 [24]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n987 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3044 (
    .a(\u2_Display/n951 ),
    .b(\u2_Display/n979 [25]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n986 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3045 (
    .a(\u2_Display/n950 ),
    .b(\u2_Display/n979 [26]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n985 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3046 (
    .a(\u2_Display/n949 ),
    .b(\u2_Display/n979 [27]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n984 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3047 (
    .a(\u2_Display/n948 ),
    .b(\u2_Display/n979 [28]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n983 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3048 (
    .a(\u2_Display/n947 ),
    .b(\u2_Display/n979 [29]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n982 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3049 (
    .a(\u2_Display/n946 ),
    .b(\u2_Display/n979 [30]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n981 ));
  EG_PHY_PAD #(
    //.LOCATION("L1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u305 (
    .do({open_n463,open_n464,open_n465,vga_b_pad[0]}),
    .opad(vga_g[0]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3050 (
    .a(\u2_Display/n945 ),
    .b(\u2_Display/n979 [31]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n980 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3051 (
    .a(\u2_Display/n2099 ),
    .b(\u2_Display/n2102 [0]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2134 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3052 (
    .a(\u2_Display/n2098 ),
    .b(\u2_Display/n2102 [1]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2133 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3053 (
    .a(\u2_Display/n2097 ),
    .b(\u2_Display/n2102 [2]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2132 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3054 (
    .a(\u2_Display/n2096 ),
    .b(\u2_Display/n2102 [3]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2131 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3055 (
    .a(\u2_Display/n2095 ),
    .b(\u2_Display/n2102 [4]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2130 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3056 (
    .a(\u2_Display/n2094 ),
    .b(\u2_Display/n2102 [5]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2129 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3057 (
    .a(\u2_Display/n2093 ),
    .b(\u2_Display/n2102 [6]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2128 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3058 (
    .a(\u2_Display/n2092 ),
    .b(\u2_Display/n2102 [7]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2127 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3059 (
    .a(\u2_Display/n2091 ),
    .b(\u2_Display/n2102 [8]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2126 ));
  EG_PHY_PAD #(
    //.LOCATION("J3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u306 (
    .do({open_n480,open_n481,open_n482,vga_hs_pad}),
    .opad(vga_hs));  // source/rtl/VGA_Demo.v(10)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3060 (
    .a(\u2_Display/n2090 ),
    .b(\u2_Display/n2102 [9]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2125 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3061 (
    .a(\u2_Display/n2089 ),
    .b(\u2_Display/n2102 [10]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2124 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3062 (
    .a(\u2_Display/n2088 ),
    .b(\u2_Display/n2102 [11]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2123 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3063 (
    .a(\u2_Display/n2087 ),
    .b(\u2_Display/n2102 [12]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2122 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3064 (
    .a(\u2_Display/n2086 ),
    .b(\u2_Display/n2102 [13]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2121 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3065 (
    .a(\u2_Display/n2085 ),
    .b(\u2_Display/n2102 [14]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2120 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3066 (
    .a(\u2_Display/n2084 ),
    .b(\u2_Display/n2102 [15]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2119 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3067 (
    .a(\u2_Display/n2083 ),
    .b(\u2_Display/n2102 [16]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2118 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3068 (
    .a(\u2_Display/n2082 ),
    .b(\u2_Display/n2102 [17]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2117 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3069 (
    .a(\u2_Display/n2081 ),
    .b(\u2_Display/n2102 [18]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2116 ));
  EG_PHY_PAD #(
    //.LOCATION("K6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u307 (
    .do({open_n497,open_n498,open_n499,vga_b_pad[0]}),
    .opad(vga_r[7]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3070 (
    .a(\u2_Display/n2080 ),
    .b(\u2_Display/n2102 [19]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2115 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3071 (
    .a(\u2_Display/n2079 ),
    .b(\u2_Display/n2102 [20]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2114 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3072 (
    .a(\u2_Display/n2078 ),
    .b(\u2_Display/n2102 [21]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2113 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3073 (
    .a(\u2_Display/n2077 ),
    .b(\u2_Display/n2102 [22]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2112 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3074 (
    .a(\u2_Display/n2076 ),
    .b(\u2_Display/n2102 [23]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2111 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3075 (
    .a(\u2_Display/n2075 ),
    .b(\u2_Display/n2102 [24]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2110 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3076 (
    .a(\u2_Display/n2074 ),
    .b(\u2_Display/n2102 [25]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2109 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3077 (
    .a(\u2_Display/n2073 ),
    .b(\u2_Display/n2102 [26]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2108 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3078 (
    .a(\u2_Display/n2072 ),
    .b(\u2_Display/n2102 [27]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2107 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3079 (
    .a(\u2_Display/n2071 ),
    .b(\u2_Display/n2102 [28]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2106 ));
  EG_PHY_PAD #(
    //.LOCATION("K3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u308 (
    .do({open_n514,open_n515,open_n516,vga_b_pad[0]}),
    .opad(vga_r[6]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3080 (
    .a(\u2_Display/n2070 ),
    .b(\u2_Display/n2102 [29]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2105 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3081 (
    .a(\u2_Display/n2069 ),
    .b(\u2_Display/n2102 [30]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2104 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3082 (
    .a(\u2_Display/n2068 ),
    .b(\u2_Display/n2102 [31]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2103 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3083 (
    .a(\u2_Display/n3222 ),
    .b(\u2_Display/n3225 [0]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3257 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3084 (
    .a(\u2_Display/n3221 ),
    .b(\u2_Display/n3225 [1]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3256 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3085 (
    .a(\u2_Display/n3220 ),
    .b(\u2_Display/n3225 [2]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3255 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3086 (
    .a(\u2_Display/n3219 ),
    .b(\u2_Display/n3225 [3]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3254 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3087 (
    .a(\u2_Display/n3218 ),
    .b(\u2_Display/n3225 [4]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3253 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3088 (
    .a(\u2_Display/n3217 ),
    .b(\u2_Display/n3225 [5]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3252 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3089 (
    .a(\u2_Display/n3216 ),
    .b(\u2_Display/n3225 [6]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3251 ));
  EG_PHY_PAD #(
    //.LOCATION("K5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u309 (
    .do({open_n531,open_n532,open_n533,vga_b_pad[0]}),
    .opad(vga_r[5]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3090 (
    .a(\u2_Display/n3215 ),
    .b(\u2_Display/n3225 [7]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3250 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3091 (
    .a(\u2_Display/n3214 ),
    .b(\u2_Display/n3225 [8]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3249 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3092 (
    .a(\u2_Display/n3213 ),
    .b(\u2_Display/n3225 [9]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3248 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3093 (
    .a(\u2_Display/n3212 ),
    .b(\u2_Display/n3225 [10]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3247 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3094 (
    .a(\u2_Display/n3211 ),
    .b(\u2_Display/n3225 [11]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3246 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3095 (
    .a(\u2_Display/n3210 ),
    .b(\u2_Display/n3225 [12]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3245 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3096 (
    .a(\u2_Display/n3209 ),
    .b(\u2_Display/n3225 [13]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3244 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3097 (
    .a(\u2_Display/n3208 ),
    .b(\u2_Display/n3225 [14]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3243 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3098 (
    .a(\u2_Display/n3207 ),
    .b(\u2_Display/n3225 [15]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3242 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3099 (
    .a(\u2_Display/n3206 ),
    .b(\u2_Display/n3225 [16]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3241 ));
  EG_PHY_PAD #(
    //.LOCATION("L4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u310 (
    .do({open_n548,open_n549,open_n550,vga_b_pad[0]}),
    .opad(vga_r[4]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3100 (
    .a(\u2_Display/n3205 ),
    .b(\u2_Display/n3225 [17]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3240 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3101 (
    .a(\u2_Display/n3204 ),
    .b(\u2_Display/n3225 [18]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3239 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3102 (
    .a(\u2_Display/n3203 ),
    .b(\u2_Display/n3225 [19]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3238 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3103 (
    .a(\u2_Display/n3202 ),
    .b(\u2_Display/n3225 [20]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3237 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3104 (
    .a(\u2_Display/n3201 ),
    .b(\u2_Display/n3225 [21]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3236 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3105 (
    .a(\u2_Display/n3200 ),
    .b(\u2_Display/n3225 [22]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3235 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3106 (
    .a(\u2_Display/n3199 ),
    .b(\u2_Display/n3225 [23]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3234 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3107 (
    .a(\u2_Display/n3198 ),
    .b(\u2_Display/n3225 [24]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3233 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3108 (
    .a(\u2_Display/n3197 ),
    .b(\u2_Display/n3225 [25]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3232 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3109 (
    .a(\u2_Display/n3196 ),
    .b(\u2_Display/n3225 [26]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3231 ));
  EG_PHY_PAD #(
    //.LOCATION("M1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u311 (
    .do({open_n565,open_n566,open_n567,vga_b_pad[0]}),
    .opad(vga_r[3]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3110 (
    .a(\u2_Display/n3195 ),
    .b(\u2_Display/n3225 [27]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3230 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3111 (
    .a(\u2_Display/n3194 ),
    .b(\u2_Display/n3225 [28]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3229 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3112 (
    .a(\u2_Display/n3193 ),
    .b(\u2_Display/n3225 [29]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3228 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3113 (
    .a(\u2_Display/n3192 ),
    .b(\u2_Display/n3225 [30]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3227 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3114 (
    .a(\u2_Display/n3191 ),
    .b(\u2_Display/n3225 [31]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3226 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3115 (
    .a(\u2_Display/n4380 ),
    .b(\u2_Display/n4383 [0]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4415 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3116 (
    .a(\u2_Display/n4379 ),
    .b(\u2_Display/n4383 [1]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4414 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3117 (
    .a(\u2_Display/n4378 ),
    .b(\u2_Display/n4383 [2]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4413 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3118 (
    .a(\u2_Display/n4377 ),
    .b(\u2_Display/n4383 [3]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4412 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3119 (
    .a(\u2_Display/n4376 ),
    .b(\u2_Display/n4383 [4]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4411 ));
  EG_PHY_PAD #(
    //.LOCATION("M2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u312 (
    .do({open_n582,open_n583,open_n584,vga_b_pad[0]}),
    .opad(vga_r[2]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3120 (
    .a(\u2_Display/n4375 ),
    .b(\u2_Display/n4383 [5]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4410 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3121 (
    .a(\u2_Display/n4374 ),
    .b(\u2_Display/n4383 [6]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4409 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3122 (
    .a(\u2_Display/n4373 ),
    .b(\u2_Display/n4383 [7]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4408 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3123 (
    .a(\u2_Display/n4372 ),
    .b(\u2_Display/n4383 [8]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4407 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3124 (
    .a(\u2_Display/n4371 ),
    .b(\u2_Display/n4383 [9]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4406 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3125 (
    .a(\u2_Display/n4370 ),
    .b(\u2_Display/n4383 [10]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4405 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3126 (
    .a(\u2_Display/n4369 ),
    .b(\u2_Display/n4383 [11]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4404 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3127 (
    .a(\u2_Display/n4368 ),
    .b(\u2_Display/n4383 [12]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4403 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3128 (
    .a(\u2_Display/n4367 ),
    .b(\u2_Display/n4383 [13]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4402 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3129 (
    .a(\u2_Display/n4366 ),
    .b(\u2_Display/n4383 [14]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4401 ));
  EG_PHY_PAD #(
    //.LOCATION("L3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u313 (
    .do({open_n599,open_n600,open_n601,vga_b_pad[0]}),
    .opad(vga_r[1]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3130 (
    .a(\u2_Display/n4365 ),
    .b(\u2_Display/n4383 [15]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4400 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3131 (
    .a(\u2_Display/n4364 ),
    .b(\u2_Display/n4383 [16]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4399 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3132 (
    .a(\u2_Display/n4363 ),
    .b(\u2_Display/n4383 [17]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4398 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3133 (
    .a(\u2_Display/n4362 ),
    .b(\u2_Display/n4383 [18]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4397 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3134 (
    .a(\u2_Display/n4361 ),
    .b(\u2_Display/n4383 [19]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4396 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3135 (
    .a(\u2_Display/n4360 ),
    .b(\u2_Display/n4383 [20]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4395 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3136 (
    .a(\u2_Display/n4359 ),
    .b(\u2_Display/n4383 [21]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4394 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3137 (
    .a(\u2_Display/n4358 ),
    .b(\u2_Display/n4383 [22]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4393 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3138 (
    .a(\u2_Display/n4357 ),
    .b(\u2_Display/n4383 [23]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4392 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3139 (
    .a(\u2_Display/n4356 ),
    .b(\u2_Display/n4383 [24]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4391 ));
  EG_PHY_PAD #(
    //.LOCATION("L5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u314 (
    .do({open_n616,open_n617,open_n618,vga_b_pad[0]}),
    .opad(vga_r[0]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3140 (
    .a(\u2_Display/n4355 ),
    .b(\u2_Display/n4383 [25]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4390 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3141 (
    .a(\u2_Display/n4354 ),
    .b(\u2_Display/n4383 [26]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4389 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3142 (
    .a(\u2_Display/n4353 ),
    .b(\u2_Display/n4383 [27]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4388 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3143 (
    .a(\u2_Display/n4352 ),
    .b(\u2_Display/n4383 [28]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4387 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3144 (
    .a(\u2_Display/n4351 ),
    .b(\u2_Display/n4383 [29]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4386 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3145 (
    .a(\u2_Display/n4350 ),
    .b(\u2_Display/n4383 [30]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4385 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3146 (
    .a(\u2_Display/n4349 ),
    .b(\u2_Display/n4383 [31]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4384 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3147 (
    .a(\u2_Display/n5503 ),
    .b(\u2_Display/n5506 [0]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5538 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3148 (
    .a(\u2_Display/n5502 ),
    .b(\u2_Display/n5506 [1]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5537 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3149 (
    .a(\u2_Display/n5501 ),
    .b(\u2_Display/n5506 [2]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5536 ));
  EG_PHY_PAD #(
    //.LOCATION("J4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u315 (
    .do({open_n633,open_n634,open_n635,vga_vs_pad}),
    .opad(vga_vs));  // source/rtl/VGA_Demo.v(11)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3150 (
    .a(\u2_Display/n5500 ),
    .b(\u2_Display/n5506 [3]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5535 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3151 (
    .a(\u2_Display/n5499 ),
    .b(\u2_Display/n5506 [4]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5534 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3152 (
    .a(\u2_Display/n5498 ),
    .b(\u2_Display/n5506 [5]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5533 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3153 (
    .a(\u2_Display/n5497 ),
    .b(\u2_Display/n5506 [6]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5532 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3154 (
    .a(\u2_Display/n5496 ),
    .b(\u2_Display/n5506 [7]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5531 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3155 (
    .a(\u2_Display/n5495 ),
    .b(\u2_Display/n5506 [8]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5530 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3156 (
    .a(\u2_Display/n5494 ),
    .b(\u2_Display/n5506 [9]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5529 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3157 (
    .a(\u2_Display/n5493 ),
    .b(\u2_Display/n5506 [10]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5528 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3158 (
    .a(\u2_Display/n5492 ),
    .b(\u2_Display/n5506 [11]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5527 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3159 (
    .a(\u2_Display/n5491 ),
    .b(\u2_Display/n5506 [12]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5526 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u316 (
    .a(\u1_Driver/n2 [9]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3160 (
    .a(\u2_Display/n5490 ),
    .b(\u2_Display/n5506 [13]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5525 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3161 (
    .a(\u2_Display/n5489 ),
    .b(\u2_Display/n5506 [14]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5524 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3162 (
    .a(\u2_Display/n5488 ),
    .b(\u2_Display/n5506 [15]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5523 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3163 (
    .a(\u2_Display/n5487 ),
    .b(\u2_Display/n5506 [16]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5522 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3164 (
    .a(\u2_Display/n5486 ),
    .b(\u2_Display/n5506 [17]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5521 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3165 (
    .a(\u2_Display/n5485 ),
    .b(\u2_Display/n5506 [18]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5520 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3166 (
    .a(\u2_Display/n5484 ),
    .b(\u2_Display/n5506 [19]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5519 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3167 (
    .a(\u2_Display/n5483 ),
    .b(\u2_Display/n5506 [20]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5518 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3168 (
    .a(\u2_Display/n5482 ),
    .b(\u2_Display/n5506 [21]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5517 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3169 (
    .a(\u2_Display/n5481 ),
    .b(\u2_Display/n5506 [22]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5516 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u317 (
    .a(\u1_Driver/n2 [8]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3170 (
    .a(\u2_Display/n5480 ),
    .b(\u2_Display/n5506 [23]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5515 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3171 (
    .a(\u2_Display/n5479 ),
    .b(\u2_Display/n5506 [24]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5514 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3172 (
    .a(\u2_Display/n5478 ),
    .b(\u2_Display/n5506 [25]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5513 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3173 (
    .a(\u2_Display/n5477 ),
    .b(\u2_Display/n5506 [26]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5512 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3174 (
    .a(\u2_Display/n5476 ),
    .b(\u2_Display/n5506 [27]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5511 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3175 (
    .a(\u2_Display/n5475 ),
    .b(\u2_Display/n5506 [28]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5510 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3176 (
    .a(\u2_Display/n5474 ),
    .b(\u2_Display/n5506 [29]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5509 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3177 (
    .a(\u2_Display/n5473 ),
    .b(\u2_Display/n5506 [30]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5508 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3178 (
    .a(\u2_Display/n5472 ),
    .b(\u2_Display/n5506 [31]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5507 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3179 (
    .a(\u2_Display/n1011 ),
    .b(\u2_Display/n1014 [0]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1046 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u318 (
    .a(\u1_Driver/n2 [7]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3180 (
    .a(\u2_Display/n1010 ),
    .b(\u2_Display/n1014 [1]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1045 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3181 (
    .a(\u2_Display/n1009 ),
    .b(\u2_Display/n1014 [2]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1044 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3182 (
    .a(\u2_Display/n1008 ),
    .b(\u2_Display/n1014 [3]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1043 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3183 (
    .a(\u2_Display/n1007 ),
    .b(\u2_Display/n1014 [4]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1042 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3184 (
    .a(\u2_Display/n1006 ),
    .b(\u2_Display/n1014 [5]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1041 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3185 (
    .a(\u2_Display/n1005 ),
    .b(\u2_Display/n1014 [6]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1040 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3186 (
    .a(\u2_Display/n1004 ),
    .b(\u2_Display/n1014 [7]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1039 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3187 (
    .a(\u2_Display/n1003 ),
    .b(\u2_Display/n1014 [8]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1038 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3188 (
    .a(\u2_Display/n1002 ),
    .b(\u2_Display/n1014 [9]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1037 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3189 (
    .a(\u2_Display/n1001 ),
    .b(\u2_Display/n1014 [10]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1036 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u319 (
    .a(\u1_Driver/n2 [6]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3190 (
    .a(\u2_Display/n1000 ),
    .b(\u2_Display/n1014 [11]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1035 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3191 (
    .a(\u2_Display/n999 ),
    .b(\u2_Display/n1014 [12]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1034 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3192 (
    .a(\u2_Display/n998 ),
    .b(\u2_Display/n1014 [13]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1033 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3193 (
    .a(\u2_Display/n997 ),
    .b(\u2_Display/n1014 [14]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1032 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3194 (
    .a(\u2_Display/n996 ),
    .b(\u2_Display/n1014 [15]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1031 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3195 (
    .a(\u2_Display/n995 ),
    .b(\u2_Display/n1014 [16]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1030 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3196 (
    .a(\u2_Display/n994 ),
    .b(\u2_Display/n1014 [17]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1029 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3197 (
    .a(\u2_Display/n993 ),
    .b(\u2_Display/n1014 [18]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1028 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3198 (
    .a(\u2_Display/n992 ),
    .b(\u2_Display/n1014 [19]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1027 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3199 (
    .a(\u2_Display/n991 ),
    .b(\u2_Display/n1014 [20]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1026 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u320 (
    .a(\u1_Driver/n2 [5]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3200 (
    .a(\u2_Display/n990 ),
    .b(\u2_Display/n1014 [21]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1025 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3201 (
    .a(\u2_Display/n989 ),
    .b(\u2_Display/n1014 [22]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1024 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3202 (
    .a(\u2_Display/n988 ),
    .b(\u2_Display/n1014 [23]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1023 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3203 (
    .a(\u2_Display/n987 ),
    .b(\u2_Display/n1014 [24]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1022 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3204 (
    .a(\u2_Display/n986 ),
    .b(\u2_Display/n1014 [25]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1021 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3205 (
    .a(\u2_Display/n985 ),
    .b(\u2_Display/n1014 [26]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1020 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3206 (
    .a(\u2_Display/n984 ),
    .b(\u2_Display/n1014 [27]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1019 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3207 (
    .a(\u2_Display/n983 ),
    .b(\u2_Display/n1014 [28]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1018 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3208 (
    .a(\u2_Display/n982 ),
    .b(\u2_Display/n1014 [29]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1017 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3209 (
    .a(\u2_Display/n981 ),
    .b(\u2_Display/n1014 [30]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1016 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u321 (
    .a(\u1_Driver/n2 [4]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3210 (
    .a(\u2_Display/n980 ),
    .b(\u2_Display/n1014 [31]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1015 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3211 (
    .a(\u2_Display/n2134 ),
    .b(\u2_Display/n2137 [0]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2169 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3212 (
    .a(\u2_Display/n2133 ),
    .b(\u2_Display/n2137 [1]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2168 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3213 (
    .a(\u2_Display/n2132 ),
    .b(\u2_Display/n2137 [2]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2167 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3214 (
    .a(\u2_Display/n2131 ),
    .b(\u2_Display/n2137 [3]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2166 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3215 (
    .a(\u2_Display/n2130 ),
    .b(\u2_Display/n2137 [4]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2165 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3216 (
    .a(\u2_Display/n2129 ),
    .b(\u2_Display/n2137 [5]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2164 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3217 (
    .a(\u2_Display/n2128 ),
    .b(\u2_Display/n2137 [6]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2163 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3218 (
    .a(\u2_Display/n2127 ),
    .b(\u2_Display/n2137 [7]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2162 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3219 (
    .a(\u2_Display/n2126 ),
    .b(\u2_Display/n2137 [8]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2161 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u322 (
    .a(\u1_Driver/n2 [3]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3220 (
    .a(\u2_Display/n2125 ),
    .b(\u2_Display/n2137 [9]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2160 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3221 (
    .a(\u2_Display/n2124 ),
    .b(\u2_Display/n2137 [10]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2159 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3222 (
    .a(\u2_Display/n2123 ),
    .b(\u2_Display/n2137 [11]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2158 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3223 (
    .a(\u2_Display/n2122 ),
    .b(\u2_Display/n2137 [12]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2157 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3224 (
    .a(\u2_Display/n2121 ),
    .b(\u2_Display/n2137 [13]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2156 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3225 (
    .a(\u2_Display/n2120 ),
    .b(\u2_Display/n2137 [14]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2155 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3226 (
    .a(\u2_Display/n2119 ),
    .b(\u2_Display/n2137 [15]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2154 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3227 (
    .a(\u2_Display/n2118 ),
    .b(\u2_Display/n2137 [16]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2153 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3228 (
    .a(\u2_Display/n2117 ),
    .b(\u2_Display/n2137 [17]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2152 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3229 (
    .a(\u2_Display/n2116 ),
    .b(\u2_Display/n2137 [18]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2151 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u323 (
    .a(\u1_Driver/n2 [2]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3230 (
    .a(\u2_Display/n2115 ),
    .b(\u2_Display/n2137 [19]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2150 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3231 (
    .a(\u2_Display/n2114 ),
    .b(\u2_Display/n2137 [20]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2149 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3232 (
    .a(\u2_Display/n2113 ),
    .b(\u2_Display/n2137 [21]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2148 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3233 (
    .a(\u2_Display/n2112 ),
    .b(\u2_Display/n2137 [22]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2147 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3234 (
    .a(\u2_Display/n2111 ),
    .b(\u2_Display/n2137 [23]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2146 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3235 (
    .a(\u2_Display/n2110 ),
    .b(\u2_Display/n2137 [24]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2145 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3236 (
    .a(\u2_Display/n2109 ),
    .b(\u2_Display/n2137 [25]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2144 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3237 (
    .a(\u2_Display/n2108 ),
    .b(\u2_Display/n2137 [26]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2143 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3238 (
    .a(\u2_Display/n2107 ),
    .b(\u2_Display/n2137 [27]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2142 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3239 (
    .a(\u2_Display/n2106 ),
    .b(\u2_Display/n2137 [28]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2141 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u324 (
    .a(\u1_Driver/n2 [11]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3240 (
    .a(\u2_Display/n2105 ),
    .b(\u2_Display/n2137 [29]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2140 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3241 (
    .a(\u2_Display/n2104 ),
    .b(\u2_Display/n2137 [30]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2139 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3242 (
    .a(\u2_Display/n2103 ),
    .b(\u2_Display/n2137 [31]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2138 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3243 (
    .a(\u2_Display/n3257 ),
    .b(\u2_Display/n3260 [0]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3292 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3244 (
    .a(\u2_Display/n3256 ),
    .b(\u2_Display/n3260 [1]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3291 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3245 (
    .a(\u2_Display/n3255 ),
    .b(\u2_Display/n3260 [2]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3290 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3246 (
    .a(\u2_Display/n3254 ),
    .b(\u2_Display/n3260 [3]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3289 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3247 (
    .a(\u2_Display/n3253 ),
    .b(\u2_Display/n3260 [4]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3288 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3248 (
    .a(\u2_Display/n3252 ),
    .b(\u2_Display/n3260 [5]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3287 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3249 (
    .a(\u2_Display/n3251 ),
    .b(\u2_Display/n3260 [6]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3286 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u325 (
    .a(\u1_Driver/n2 [10]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3250 (
    .a(\u2_Display/n3250 ),
    .b(\u2_Display/n3260 [7]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3285 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3251 (
    .a(\u2_Display/n3249 ),
    .b(\u2_Display/n3260 [8]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3284 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3252 (
    .a(\u2_Display/n3248 ),
    .b(\u2_Display/n3260 [9]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3283 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3253 (
    .a(\u2_Display/n3247 ),
    .b(\u2_Display/n3260 [10]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3282 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3254 (
    .a(\u2_Display/n3246 ),
    .b(\u2_Display/n3260 [11]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3281 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3255 (
    .a(\u2_Display/n3245 ),
    .b(\u2_Display/n3260 [12]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3280 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3256 (
    .a(\u2_Display/n3244 ),
    .b(\u2_Display/n3260 [13]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3279 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3257 (
    .a(\u2_Display/n3243 ),
    .b(\u2_Display/n3260 [14]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3278 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3258 (
    .a(\u2_Display/n3242 ),
    .b(\u2_Display/n3260 [15]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3277 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3259 (
    .a(\u2_Display/n3241 ),
    .b(\u2_Display/n3260 [16]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3276 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u326 (
    .a(\u1_Driver/n2 [1]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3260 (
    .a(\u2_Display/n3240 ),
    .b(\u2_Display/n3260 [17]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3275 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3261 (
    .a(\u2_Display/n3239 ),
    .b(\u2_Display/n3260 [18]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3274 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3262 (
    .a(\u2_Display/n3238 ),
    .b(\u2_Display/n3260 [19]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3273 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3263 (
    .a(\u2_Display/n3237 ),
    .b(\u2_Display/n3260 [20]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3272 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3264 (
    .a(\u2_Display/n3236 ),
    .b(\u2_Display/n3260 [21]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3271 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3265 (
    .a(\u2_Display/n3235 ),
    .b(\u2_Display/n3260 [22]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3270 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3266 (
    .a(\u2_Display/n3234 ),
    .b(\u2_Display/n3260 [23]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3269 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3267 (
    .a(\u2_Display/n3233 ),
    .b(\u2_Display/n3260 [24]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3268 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3268 (
    .a(\u2_Display/n3232 ),
    .b(\u2_Display/n3260 [25]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3267 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3269 (
    .a(\u2_Display/n3231 ),
    .b(\u2_Display/n3260 [26]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3266 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u327 (
    .a(\u1_Driver/n2 [0]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3270 (
    .a(\u2_Display/n3230 ),
    .b(\u2_Display/n3260 [27]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3265 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3271 (
    .a(\u2_Display/n3229 ),
    .b(\u2_Display/n3260 [28]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3264 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3272 (
    .a(\u2_Display/n3228 ),
    .b(\u2_Display/n3260 [29]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3263 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3273 (
    .a(\u2_Display/n3227 ),
    .b(\u2_Display/n3260 [30]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3262 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3274 (
    .a(\u2_Display/n3226 ),
    .b(\u2_Display/n3260 [31]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3261 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3275 (
    .a(\u2_Display/n4415 ),
    .b(\u2_Display/n4418 [0]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4450 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3276 (
    .a(\u2_Display/n4414 ),
    .b(\u2_Display/n4418 [1]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4449 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3277 (
    .a(\u2_Display/n4413 ),
    .b(\u2_Display/n4418 [2]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4448 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3278 (
    .a(\u2_Display/n4412 ),
    .b(\u2_Display/n4418 [3]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4447 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3279 (
    .a(\u2_Display/n4411 ),
    .b(\u2_Display/n4418 [4]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4446 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u328 (
    .a(\u2_Display/i [10]),
    .b(\u2_Display/i [9]),
    .o(\u2_Display/add7_2_co ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3280 (
    .a(\u2_Display/n4410 ),
    .b(\u2_Display/n4418 [5]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4445 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3281 (
    .a(\u2_Display/n4409 ),
    .b(\u2_Display/n4418 [6]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4444 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3282 (
    .a(\u2_Display/n4408 ),
    .b(\u2_Display/n4418 [7]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4443 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3283 (
    .a(\u2_Display/n4407 ),
    .b(\u2_Display/n4418 [8]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4442 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3284 (
    .a(\u2_Display/n4406 ),
    .b(\u2_Display/n4418 [9]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4441 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3285 (
    .a(\u2_Display/n4405 ),
    .b(\u2_Display/n4418 [10]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4440 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3286 (
    .a(\u2_Display/n4404 ),
    .b(\u2_Display/n4418 [11]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4439 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3287 (
    .a(\u2_Display/n4403 ),
    .b(\u2_Display/n4418 [12]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4438 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3288 (
    .a(\u2_Display/n4402 ),
    .b(\u2_Display/n4418 [13]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4437 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3289 (
    .a(\u2_Display/n4401 ),
    .b(\u2_Display/n4418 [14]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4436 ));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u329 (
    .a(\u2_Display/i [10]),
    .b(\u2_Display/i [9]),
    .o(\u2_Display/n140 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3290 (
    .a(\u2_Display/n4400 ),
    .b(\u2_Display/n4418 [15]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4435 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3291 (
    .a(\u2_Display/n4399 ),
    .b(\u2_Display/n4418 [16]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4434 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3292 (
    .a(\u2_Display/n4398 ),
    .b(\u2_Display/n4418 [17]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4433 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3293 (
    .a(\u2_Display/n4397 ),
    .b(\u2_Display/n4418 [18]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4432 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3294 (
    .a(\u2_Display/n4396 ),
    .b(\u2_Display/n4418 [19]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4431 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3295 (
    .a(\u2_Display/n4395 ),
    .b(\u2_Display/n4418 [20]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4430 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3296 (
    .a(\u2_Display/n4394 ),
    .b(\u2_Display/n4418 [21]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4429 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3297 (
    .a(\u2_Display/n4393 ),
    .b(\u2_Display/n4418 [22]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4428 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3298 (
    .a(\u2_Display/n4392 ),
    .b(\u2_Display/n4418 [23]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4427 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3299 (
    .a(\u2_Display/n4391 ),
    .b(\u2_Display/n4418 [24]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4426 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u330 (
    .a(\u1_Driver/n11 ),
    .b(\u1_Driver/n12 ),
    .c(\u1_Driver/n14 ),
    .d(\u1_Driver/n15 ),
    .o(vga_de_pad));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3300 (
    .a(\u2_Display/n4390 ),
    .b(\u2_Display/n4418 [25]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4425 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3301 (
    .a(\u2_Display/n4389 ),
    .b(\u2_Display/n4418 [26]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4424 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3302 (
    .a(\u2_Display/n4388 ),
    .b(\u2_Display/n4418 [27]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4423 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3303 (
    .a(\u2_Display/n4387 ),
    .b(\u2_Display/n4418 [28]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4422 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3304 (
    .a(\u2_Display/n4386 ),
    .b(\u2_Display/n4418 [29]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4421 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3305 (
    .a(\u2_Display/n4385 ),
    .b(\u2_Display/n4418 [30]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4420 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3306 (
    .a(\u2_Display/n4384 ),
    .b(\u2_Display/n4418 [31]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4419 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3307 (
    .a(\u2_Display/n5538 ),
    .b(\u2_Display/n5541 [0]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5573 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3308 (
    .a(\u2_Display/n5537 ),
    .b(\u2_Display/n5541 [1]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5572 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3309 (
    .a(\u2_Display/n5536 ),
    .b(\u2_Display/n5541 [2]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5571 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u331 (
    .a(\u2_Display/n3788 [0]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [0]),
    .o(\u2_Display/n3820 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3310 (
    .a(\u2_Display/n5535 ),
    .b(\u2_Display/n5541 [3]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5570 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3311 (
    .a(\u2_Display/n5534 ),
    .b(\u2_Display/n5541 [4]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5569 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3312 (
    .a(\u2_Display/n5533 ),
    .b(\u2_Display/n5541 [5]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5568 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3313 (
    .a(\u2_Display/n5532 ),
    .b(\u2_Display/n5541 [6]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5567 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3314 (
    .a(\u2_Display/n5531 ),
    .b(\u2_Display/n5541 [7]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5566 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3315 (
    .a(\u2_Display/n5530 ),
    .b(\u2_Display/n5541 [8]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5565 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3316 (
    .a(\u2_Display/n5529 ),
    .b(\u2_Display/n5541 [9]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5564 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3317 (
    .a(\u2_Display/n5528 ),
    .b(\u2_Display/n5541 [10]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5563 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3318 (
    .a(\u2_Display/n5527 ),
    .b(\u2_Display/n5541 [11]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5562 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3319 (
    .a(\u2_Display/n5526 ),
    .b(\u2_Display/n5541 [12]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5561 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u332 (
    .a(\u2_Display/n3788 [1]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [1]),
    .o(\u2_Display/n3819 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3320 (
    .a(\u2_Display/n5525 ),
    .b(\u2_Display/n5541 [13]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5560 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3321 (
    .a(\u2_Display/n5524 ),
    .b(\u2_Display/n5541 [14]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5559 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3322 (
    .a(\u2_Display/n5523 ),
    .b(\u2_Display/n5541 [15]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5558 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3323 (
    .a(\u2_Display/n5522 ),
    .b(\u2_Display/n5541 [16]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5557 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3324 (
    .a(\u2_Display/n5521 ),
    .b(\u2_Display/n5541 [17]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5556 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3325 (
    .a(\u2_Display/n5520 ),
    .b(\u2_Display/n5541 [18]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5555 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3326 (
    .a(\u2_Display/n5519 ),
    .b(\u2_Display/n5541 [19]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5554 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3327 (
    .a(\u2_Display/n5518 ),
    .b(\u2_Display/n5541 [20]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5553 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3328 (
    .a(\u2_Display/n5517 ),
    .b(\u2_Display/n5541 [21]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5552 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3329 (
    .a(\u2_Display/n5516 ),
    .b(\u2_Display/n5541 [22]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5551 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u333 (
    .a(\u2_Display/n3788 [2]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [2]),
    .o(\u2_Display/n3818 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3330 (
    .a(\u2_Display/n5515 ),
    .b(\u2_Display/n5541 [23]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5550 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3331 (
    .a(\u2_Display/n5514 ),
    .b(\u2_Display/n5541 [24]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5549 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3332 (
    .a(\u2_Display/n5513 ),
    .b(\u2_Display/n5541 [25]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5548 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3333 (
    .a(\u2_Display/n5512 ),
    .b(\u2_Display/n5541 [26]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5547 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3334 (
    .a(\u2_Display/n5511 ),
    .b(\u2_Display/n5541 [27]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5546 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3335 (
    .a(\u2_Display/n5510 ),
    .b(\u2_Display/n5541 [28]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5545 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3336 (
    .a(\u2_Display/n5509 ),
    .b(\u2_Display/n5541 [29]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5544 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3337 (
    .a(\u2_Display/n5508 ),
    .b(\u2_Display/n5541 [30]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5543 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3338 (
    .a(\u2_Display/n5507 ),
    .b(\u2_Display/n5541 [31]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5542 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3339 (
    .a(\u2_Display/n1046 ),
    .b(\u2_Display/n1049 [0]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1081 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u334 (
    .a(\u2_Display/n3788 [3]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [3]),
    .o(\u2_Display/n3817 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3340 (
    .a(\u2_Display/n1045 ),
    .b(\u2_Display/n1049 [1]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1080 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3341 (
    .a(\u2_Display/n1044 ),
    .b(\u2_Display/n1049 [2]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1079 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3342 (
    .a(\u2_Display/n1043 ),
    .b(\u2_Display/n1049 [3]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1078 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3343 (
    .a(\u2_Display/n1042 ),
    .b(\u2_Display/n1049 [4]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1077 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3344 (
    .a(\u2_Display/n1041 ),
    .b(\u2_Display/n1049 [5]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1076 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3345 (
    .a(\u2_Display/n1040 ),
    .b(\u2_Display/n1049 [6]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1075 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3346 (
    .a(\u2_Display/n1039 ),
    .b(\u2_Display/n1049 [7]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1074 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3347 (
    .a(\u2_Display/n1038 ),
    .b(\u2_Display/n1049 [8]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1073 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3348 (
    .a(\u2_Display/n1037 ),
    .b(\u2_Display/n1049 [9]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1072 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3349 (
    .a(\u2_Display/n1036 ),
    .b(\u2_Display/n1049 [10]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1071 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u335 (
    .a(\u2_Display/n3788 [4]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [4]),
    .o(\u2_Display/n3816 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3350 (
    .a(\u2_Display/n1035 ),
    .b(\u2_Display/n1049 [11]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1070 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3351 (
    .a(\u2_Display/n1034 ),
    .b(\u2_Display/n1049 [12]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1069 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3352 (
    .a(\u2_Display/n1033 ),
    .b(\u2_Display/n1049 [13]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1068 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3353 (
    .a(\u2_Display/n1032 ),
    .b(\u2_Display/n1049 [14]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1067 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3354 (
    .a(\u2_Display/n1031 ),
    .b(\u2_Display/n1049 [15]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1066 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3355 (
    .a(\u2_Display/n1030 ),
    .b(\u2_Display/n1049 [16]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1065 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3356 (
    .a(\u2_Display/n1029 ),
    .b(\u2_Display/n1049 [17]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1064 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3357 (
    .a(\u2_Display/n1028 ),
    .b(\u2_Display/n1049 [18]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1063 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3358 (
    .a(\u2_Display/n1027 ),
    .b(\u2_Display/n1049 [19]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1062 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3359 (
    .a(\u2_Display/n1026 ),
    .b(\u2_Display/n1049 [20]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1061 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u336 (
    .a(\u2_Display/n3788 [5]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [5]),
    .o(\u2_Display/n3815 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3360 (
    .a(\u2_Display/n1025 ),
    .b(\u2_Display/n1049 [21]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1060 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3361 (
    .a(\u2_Display/n1024 ),
    .b(\u2_Display/n1049 [22]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1059 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3362 (
    .a(\u2_Display/n1023 ),
    .b(\u2_Display/n1049 [23]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1058 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3363 (
    .a(\u2_Display/n1022 ),
    .b(\u2_Display/n1049 [24]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1057 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3364 (
    .a(\u2_Display/n1021 ),
    .b(\u2_Display/n1049 [25]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1056 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3365 (
    .a(\u2_Display/n1020 ),
    .b(\u2_Display/n1049 [26]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1055 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3366 (
    .a(\u2_Display/n1019 ),
    .b(\u2_Display/n1049 [27]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1054 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3367 (
    .a(\u2_Display/n1018 ),
    .b(\u2_Display/n1049 [28]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1053 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3368 (
    .a(\u2_Display/n1017 ),
    .b(\u2_Display/n1049 [29]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1052 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3369 (
    .a(\u2_Display/n1016 ),
    .b(\u2_Display/n1049 [30]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1051 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u337 (
    .a(\u2_Display/n3788 [6]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [6]),
    .o(\u2_Display/n3814 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3370 (
    .a(\u2_Display/n1015 ),
    .b(\u2_Display/n1049 [31]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1050 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3371 (
    .a(\u2_Display/n2169 ),
    .b(\u2_Display/n2172 [0]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2204 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3372 (
    .a(\u2_Display/n2168 ),
    .b(\u2_Display/n2172 [1]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2203 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3373 (
    .a(\u2_Display/n2167 ),
    .b(\u2_Display/n2172 [2]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2202 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3374 (
    .a(\u2_Display/n2166 ),
    .b(\u2_Display/n2172 [3]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2201 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3375 (
    .a(\u2_Display/n2165 ),
    .b(\u2_Display/n2172 [4]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2200 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3376 (
    .a(\u2_Display/n2164 ),
    .b(\u2_Display/n2172 [5]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2199 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3377 (
    .a(\u2_Display/n2163 ),
    .b(\u2_Display/n2172 [6]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2198 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3378 (
    .a(\u2_Display/n2162 ),
    .b(\u2_Display/n2172 [7]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2197 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3379 (
    .a(\u2_Display/n2161 ),
    .b(\u2_Display/n2172 [8]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2196 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u338 (
    .a(\u2_Display/n3788 [7]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [7]),
    .o(\u2_Display/n3813 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3380 (
    .a(\u2_Display/n2160 ),
    .b(\u2_Display/n2172 [9]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2195 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3381 (
    .a(\u2_Display/n2159 ),
    .b(\u2_Display/n2172 [10]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2194 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3382 (
    .a(\u2_Display/n2158 ),
    .b(\u2_Display/n2172 [11]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2193 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3383 (
    .a(\u2_Display/n2157 ),
    .b(\u2_Display/n2172 [12]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2192 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3384 (
    .a(\u2_Display/n2156 ),
    .b(\u2_Display/n2172 [13]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2191 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3385 (
    .a(\u2_Display/n2155 ),
    .b(\u2_Display/n2172 [14]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2190 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3386 (
    .a(\u2_Display/n2154 ),
    .b(\u2_Display/n2172 [15]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2189 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3387 (
    .a(\u2_Display/n2153 ),
    .b(\u2_Display/n2172 [16]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2188 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3388 (
    .a(\u2_Display/n2152 ),
    .b(\u2_Display/n2172 [17]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2187 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3389 (
    .a(\u2_Display/n2151 ),
    .b(\u2_Display/n2172 [18]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2186 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u339 (
    .a(\u2_Display/n3788 [8]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [8]),
    .o(\u2_Display/n3812 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3390 (
    .a(\u2_Display/n2150 ),
    .b(\u2_Display/n2172 [19]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2185 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3391 (
    .a(\u2_Display/n2149 ),
    .b(\u2_Display/n2172 [20]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2184 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3392 (
    .a(\u2_Display/n2148 ),
    .b(\u2_Display/n2172 [21]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2183 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3393 (
    .a(\u2_Display/n2147 ),
    .b(\u2_Display/n2172 [22]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2182 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3394 (
    .a(\u2_Display/n2146 ),
    .b(\u2_Display/n2172 [23]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2181 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3395 (
    .a(\u2_Display/n2145 ),
    .b(\u2_Display/n2172 [24]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2180 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3396 (
    .a(\u2_Display/n2144 ),
    .b(\u2_Display/n2172 [25]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2179 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3397 (
    .a(\u2_Display/n2143 ),
    .b(\u2_Display/n2172 [26]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2178 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3398 (
    .a(\u2_Display/n2142 ),
    .b(\u2_Display/n2172 [27]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2177 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3399 (
    .a(\u2_Display/n2141 ),
    .b(\u2_Display/n2172 [28]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2176 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u340 (
    .a(\u2_Display/n3788 [9]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [9]),
    .o(\u2_Display/n3811 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3400 (
    .a(\u2_Display/n2140 ),
    .b(\u2_Display/n2172 [29]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2175 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3401 (
    .a(\u2_Display/n2139 ),
    .b(\u2_Display/n2172 [30]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2174 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3402 (
    .a(\u2_Display/n2138 ),
    .b(\u2_Display/n2172 [31]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2173 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3403 (
    .a(\u2_Display/n3292 ),
    .b(\u2_Display/n3295 [0]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3327 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3404 (
    .a(\u2_Display/n3291 ),
    .b(\u2_Display/n3295 [1]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3326 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3405 (
    .a(\u2_Display/n3290 ),
    .b(\u2_Display/n3295 [2]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3325 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3406 (
    .a(\u2_Display/n3289 ),
    .b(\u2_Display/n3295 [3]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3324 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3407 (
    .a(\u2_Display/n3288 ),
    .b(\u2_Display/n3295 [4]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3323 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3408 (
    .a(\u2_Display/n3287 ),
    .b(\u2_Display/n3295 [5]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3322 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3409 (
    .a(\u2_Display/n3286 ),
    .b(\u2_Display/n3295 [6]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3321 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u341 (
    .a(\u2_Display/n3788 [10]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [10]),
    .o(\u2_Display/n3810 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3410 (
    .a(\u2_Display/n3285 ),
    .b(\u2_Display/n3295 [7]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3320 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3411 (
    .a(\u2_Display/n3284 ),
    .b(\u2_Display/n3295 [8]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3319 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3412 (
    .a(\u2_Display/n3283 ),
    .b(\u2_Display/n3295 [9]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3318 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3413 (
    .a(\u2_Display/n3282 ),
    .b(\u2_Display/n3295 [10]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3317 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3414 (
    .a(\u2_Display/n3281 ),
    .b(\u2_Display/n3295 [11]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3316 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3415 (
    .a(\u2_Display/n3280 ),
    .b(\u2_Display/n3295 [12]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3315 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3416 (
    .a(\u2_Display/n3279 ),
    .b(\u2_Display/n3295 [13]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3314 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3417 (
    .a(\u2_Display/n3278 ),
    .b(\u2_Display/n3295 [14]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3313 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3418 (
    .a(\u2_Display/n3277 ),
    .b(\u2_Display/n3295 [15]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3312 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3419 (
    .a(\u2_Display/n3276 ),
    .b(\u2_Display/n3295 [16]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3311 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u342 (
    .a(\u2_Display/n3788 [11]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [11]),
    .o(\u2_Display/n3809 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3420 (
    .a(\u2_Display/n3275 ),
    .b(\u2_Display/n3295 [17]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3310 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3421 (
    .a(\u2_Display/n3274 ),
    .b(\u2_Display/n3295 [18]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3309 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3422 (
    .a(\u2_Display/n3273 ),
    .b(\u2_Display/n3295 [19]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3308 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3423 (
    .a(\u2_Display/n3272 ),
    .b(\u2_Display/n3295 [20]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3307 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3424 (
    .a(\u2_Display/n3271 ),
    .b(\u2_Display/n3295 [21]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3306 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3425 (
    .a(\u2_Display/n3270 ),
    .b(\u2_Display/n3295 [22]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3305 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3426 (
    .a(\u2_Display/n3269 ),
    .b(\u2_Display/n3295 [23]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3304 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3427 (
    .a(\u2_Display/n3268 ),
    .b(\u2_Display/n3295 [24]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3303 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3428 (
    .a(\u2_Display/n3267 ),
    .b(\u2_Display/n3295 [25]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3302 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3429 (
    .a(\u2_Display/n3266 ),
    .b(\u2_Display/n3295 [26]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3301 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u343 (
    .a(\u2_Display/n3788 [12]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [12]),
    .o(\u2_Display/n3808 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3430 (
    .a(\u2_Display/n3265 ),
    .b(\u2_Display/n3295 [27]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3300 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3431 (
    .a(\u2_Display/n3264 ),
    .b(\u2_Display/n3295 [28]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3299 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3432 (
    .a(\u2_Display/n3263 ),
    .b(\u2_Display/n3295 [29]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3298 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3433 (
    .a(\u2_Display/n3262 ),
    .b(\u2_Display/n3295 [30]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3297 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3434 (
    .a(\u2_Display/n3261 ),
    .b(\u2_Display/n3295 [31]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3296 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3435 (
    .a(\u2_Display/n4450 ),
    .b(\u2_Display/n4453 [0]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4485 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3436 (
    .a(\u2_Display/n4449 ),
    .b(\u2_Display/n4453 [1]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4484 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3437 (
    .a(\u2_Display/n4448 ),
    .b(\u2_Display/n4453 [2]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4483 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3438 (
    .a(\u2_Display/n4447 ),
    .b(\u2_Display/n4453 [3]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4482 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3439 (
    .a(\u2_Display/n4446 ),
    .b(\u2_Display/n4453 [4]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4481 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u344 (
    .a(\u2_Display/n3788 [13]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [13]),
    .o(\u2_Display/n3807 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3440 (
    .a(\u2_Display/n4445 ),
    .b(\u2_Display/n4453 [5]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4480 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3441 (
    .a(\u2_Display/n4444 ),
    .b(\u2_Display/n4453 [6]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4479 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3442 (
    .a(\u2_Display/n4443 ),
    .b(\u2_Display/n4453 [7]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4478 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3443 (
    .a(\u2_Display/n4442 ),
    .b(\u2_Display/n4453 [8]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4477 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3444 (
    .a(\u2_Display/n4441 ),
    .b(\u2_Display/n4453 [9]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4476 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3445 (
    .a(\u2_Display/n4440 ),
    .b(\u2_Display/n4453 [10]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4475 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3446 (
    .a(\u2_Display/n4439 ),
    .b(\u2_Display/n4453 [11]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4474 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3447 (
    .a(\u2_Display/n4438 ),
    .b(\u2_Display/n4453 [12]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4473 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3448 (
    .a(\u2_Display/n4437 ),
    .b(\u2_Display/n4453 [13]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4472 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3449 (
    .a(\u2_Display/n4436 ),
    .b(\u2_Display/n4453 [14]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4471 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u345 (
    .a(\u2_Display/n3788 [14]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [14]),
    .o(\u2_Display/n3806 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3450 (
    .a(\u2_Display/n4435 ),
    .b(\u2_Display/n4453 [15]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4470 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3451 (
    .a(\u2_Display/n4434 ),
    .b(\u2_Display/n4453 [16]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4469 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3452 (
    .a(\u2_Display/n4433 ),
    .b(\u2_Display/n4453 [17]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4468 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3453 (
    .a(\u2_Display/n4432 ),
    .b(\u2_Display/n4453 [18]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4467 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3454 (
    .a(\u2_Display/n4431 ),
    .b(\u2_Display/n4453 [19]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4466 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3455 (
    .a(\u2_Display/n4430 ),
    .b(\u2_Display/n4453 [20]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4465 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3456 (
    .a(\u2_Display/n4429 ),
    .b(\u2_Display/n4453 [21]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4464 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3457 (
    .a(\u2_Display/n4428 ),
    .b(\u2_Display/n4453 [22]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4463 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3458 (
    .a(\u2_Display/n4427 ),
    .b(\u2_Display/n4453 [23]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4462 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3459 (
    .a(\u2_Display/n4426 ),
    .b(\u2_Display/n4453 [24]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4461 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u346 (
    .a(\u2_Display/n3788 [15]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [15]),
    .o(\u2_Display/n3805 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3460 (
    .a(\u2_Display/n4425 ),
    .b(\u2_Display/n4453 [25]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4460 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3461 (
    .a(\u2_Display/n4424 ),
    .b(\u2_Display/n4453 [26]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4459 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3462 (
    .a(\u2_Display/n4423 ),
    .b(\u2_Display/n4453 [27]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4458 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3463 (
    .a(\u2_Display/n4422 ),
    .b(\u2_Display/n4453 [28]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4457 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3464 (
    .a(\u2_Display/n4421 ),
    .b(\u2_Display/n4453 [29]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4456 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3465 (
    .a(\u2_Display/n4420 ),
    .b(\u2_Display/n4453 [30]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4455 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3466 (
    .a(\u2_Display/n4419 ),
    .b(\u2_Display/n4453 [31]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4454 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3467 (
    .a(\u2_Display/n5573 ),
    .b(\u2_Display/n5576 [0]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5608 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3468 (
    .a(\u2_Display/n5572 ),
    .b(\u2_Display/n5576 [1]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5607 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3469 (
    .a(\u2_Display/n5571 ),
    .b(\u2_Display/n5576 [2]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5606 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u347 (
    .a(\u2_Display/n3788 [16]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [16]),
    .o(\u2_Display/n3804 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3470 (
    .a(\u2_Display/n5570 ),
    .b(\u2_Display/n5576 [3]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5605 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3471 (
    .a(\u2_Display/n5569 ),
    .b(\u2_Display/n5576 [4]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5604 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3472 (
    .a(\u2_Display/n5568 ),
    .b(\u2_Display/n5576 [5]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5603 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3473 (
    .a(\u2_Display/n5567 ),
    .b(\u2_Display/n5576 [6]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5602 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3474 (
    .a(\u2_Display/n5566 ),
    .b(\u2_Display/n5576 [7]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5601 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3475 (
    .a(\u2_Display/n5565 ),
    .b(\u2_Display/n5576 [8]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5600 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3476 (
    .a(\u2_Display/n5564 ),
    .b(\u2_Display/n5576 [9]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5599 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3477 (
    .a(\u2_Display/n5563 ),
    .b(\u2_Display/n5576 [10]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5598 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3478 (
    .a(\u2_Display/n5562 ),
    .b(\u2_Display/n5576 [11]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5597 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3479 (
    .a(\u2_Display/n5561 ),
    .b(\u2_Display/n5576 [12]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5596 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u348 (
    .a(\u2_Display/n3788 [17]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [17]),
    .o(\u2_Display/n3803 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3480 (
    .a(\u2_Display/n5560 ),
    .b(\u2_Display/n5576 [13]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5595 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3481 (
    .a(\u2_Display/n5559 ),
    .b(\u2_Display/n5576 [14]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5594 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3482 (
    .a(\u2_Display/n5558 ),
    .b(\u2_Display/n5576 [15]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5593 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3483 (
    .a(\u2_Display/n5557 ),
    .b(\u2_Display/n5576 [16]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5592 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3484 (
    .a(\u2_Display/n5556 ),
    .b(\u2_Display/n5576 [17]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5591 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3485 (
    .a(\u2_Display/n5555 ),
    .b(\u2_Display/n5576 [18]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5590 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3486 (
    .a(\u2_Display/n5554 ),
    .b(\u2_Display/n5576 [19]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5589 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3487 (
    .a(\u2_Display/n5553 ),
    .b(\u2_Display/n5576 [20]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5588 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3488 (
    .a(\u2_Display/n5552 ),
    .b(\u2_Display/n5576 [21]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5587 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3489 (
    .a(\u2_Display/n5551 ),
    .b(\u2_Display/n5576 [22]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5586 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u349 (
    .a(\u2_Display/n3788 [18]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [18]),
    .o(\u2_Display/n3802 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3490 (
    .a(\u2_Display/n5550 ),
    .b(\u2_Display/n5576 [23]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5585 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3491 (
    .a(\u2_Display/n5549 ),
    .b(\u2_Display/n5576 [24]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5584 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3492 (
    .a(\u2_Display/n5548 ),
    .b(\u2_Display/n5576 [25]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5583 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3493 (
    .a(\u2_Display/n5547 ),
    .b(\u2_Display/n5576 [26]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5582 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3494 (
    .a(\u2_Display/n5546 ),
    .b(\u2_Display/n5576 [27]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5581 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3495 (
    .a(\u2_Display/n5545 ),
    .b(\u2_Display/n5576 [28]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5580 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3496 (
    .a(\u2_Display/n5544 ),
    .b(\u2_Display/n5576 [29]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5579 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3497 (
    .a(\u2_Display/n5543 ),
    .b(\u2_Display/n5576 [30]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5578 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3498 (
    .a(\u2_Display/n5542 ),
    .b(\u2_Display/n5576 [31]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5577 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3499 (
    .a(\u2_Display/n1081 ),
    .b(\u2_Display/n1084 [0]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1116 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u350 (
    .a(\u2_Display/n3788 [19]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [19]),
    .o(\u2_Display/n3801 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3500 (
    .a(\u2_Display/n1080 ),
    .b(\u2_Display/n1084 [1]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1115 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3501 (
    .a(\u2_Display/n1079 ),
    .b(\u2_Display/n1084 [2]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1114 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3502 (
    .a(\u2_Display/n1078 ),
    .b(\u2_Display/n1084 [3]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1113 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3503 (
    .a(\u2_Display/n1077 ),
    .b(\u2_Display/n1084 [4]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1112 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3504 (
    .a(\u2_Display/n1076 ),
    .b(\u2_Display/n1084 [5]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1111 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3505 (
    .a(\u2_Display/n1075 ),
    .b(\u2_Display/n1084 [6]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1110 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3506 (
    .a(\u2_Display/n1074 ),
    .b(\u2_Display/n1084 [7]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1109 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3507 (
    .a(\u2_Display/n1073 ),
    .b(\u2_Display/n1084 [8]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1108 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3508 (
    .a(\u2_Display/n1072 ),
    .b(\u2_Display/n1084 [9]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1107 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3509 (
    .a(\u2_Display/n1071 ),
    .b(\u2_Display/n1084 [10]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1106 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u351 (
    .a(\u2_Display/n3788 [20]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [20]),
    .o(\u2_Display/n3800 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3510 (
    .a(\u2_Display/n1070 ),
    .b(\u2_Display/n1084 [11]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1105 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3511 (
    .a(\u2_Display/n1069 ),
    .b(\u2_Display/n1084 [12]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1104 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3512 (
    .a(\u2_Display/n1068 ),
    .b(\u2_Display/n1084 [13]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1103 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3513 (
    .a(\u2_Display/n1067 ),
    .b(\u2_Display/n1084 [14]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1102 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3514 (
    .a(\u2_Display/n1066 ),
    .b(\u2_Display/n1084 [15]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1101 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3515 (
    .a(\u2_Display/n1065 ),
    .b(\u2_Display/n1084 [16]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1100 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3516 (
    .a(\u2_Display/n1064 ),
    .b(\u2_Display/n1084 [17]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1099 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3517 (
    .a(\u2_Display/n1063 ),
    .b(\u2_Display/n1084 [18]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1098 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3518 (
    .a(\u2_Display/n1062 ),
    .b(\u2_Display/n1084 [19]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1097 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3519 (
    .a(\u2_Display/n1061 ),
    .b(\u2_Display/n1084 [20]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1096 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u352 (
    .a(\u2_Display/n3788 [21]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [21]),
    .o(\u2_Display/n3799 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3520 (
    .a(\u2_Display/n1060 ),
    .b(\u2_Display/n1084 [21]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1095 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3521 (
    .a(\u2_Display/n1059 ),
    .b(\u2_Display/n1084 [22]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1094 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3522 (
    .a(\u2_Display/n1058 ),
    .b(\u2_Display/n1084 [23]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1093 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3523 (
    .a(\u2_Display/n1057 ),
    .b(\u2_Display/n1084 [24]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1092 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3524 (
    .a(\u2_Display/n1056 ),
    .b(\u2_Display/n1084 [25]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1091 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3525 (
    .a(\u2_Display/n1055 ),
    .b(\u2_Display/n1084 [26]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1090 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3526 (
    .a(\u2_Display/n1054 ),
    .b(\u2_Display/n1084 [27]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1089 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3527 (
    .a(\u2_Display/n1053 ),
    .b(\u2_Display/n1084 [28]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1088 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3528 (
    .a(\u2_Display/n1052 ),
    .b(\u2_Display/n1084 [29]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1087 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3529 (
    .a(\u2_Display/n1051 ),
    .b(\u2_Display/n1084 [30]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1086 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u353 (
    .a(\u2_Display/n3788 [22]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [22]),
    .o(\u2_Display/n3798 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3530 (
    .a(\u2_Display/n1050 ),
    .b(\u2_Display/n1084 [31]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1085 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3531 (
    .a(\u2_Display/n2204 ),
    .b(\u2_Display/n2207 [0]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2239 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3532 (
    .a(\u2_Display/n2203 ),
    .b(\u2_Display/n2207 [1]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2238 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3533 (
    .a(\u2_Display/n2202 ),
    .b(\u2_Display/n2207 [2]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2237 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3534 (
    .a(\u2_Display/n2201 ),
    .b(\u2_Display/n2207 [3]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2236 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3535 (
    .a(\u2_Display/n2200 ),
    .b(\u2_Display/n2207 [4]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2235 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3536 (
    .a(\u2_Display/n2199 ),
    .b(\u2_Display/n2207 [5]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2234 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3537 (
    .a(\u2_Display/n2198 ),
    .b(\u2_Display/n2207 [6]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2233 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3538 (
    .a(\u2_Display/n2197 ),
    .b(\u2_Display/n2207 [7]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2232 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3539 (
    .a(\u2_Display/n2196 ),
    .b(\u2_Display/n2207 [8]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2231 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u354 (
    .a(\u2_Display/n3788 [23]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [23]),
    .o(\u2_Display/n3797 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3540 (
    .a(\u2_Display/n2195 ),
    .b(\u2_Display/n2207 [9]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2230 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3541 (
    .a(\u2_Display/n2194 ),
    .b(\u2_Display/n2207 [10]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2229 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3542 (
    .a(\u2_Display/n2193 ),
    .b(\u2_Display/n2207 [11]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2228 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3543 (
    .a(\u2_Display/n2192 ),
    .b(\u2_Display/n2207 [12]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2227 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3544 (
    .a(\u2_Display/n2191 ),
    .b(\u2_Display/n2207 [13]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2226 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3545 (
    .a(\u2_Display/n2190 ),
    .b(\u2_Display/n2207 [14]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2225 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3546 (
    .a(\u2_Display/n2189 ),
    .b(\u2_Display/n2207 [15]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2224 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3547 (
    .a(\u2_Display/n2188 ),
    .b(\u2_Display/n2207 [16]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2223 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3548 (
    .a(\u2_Display/n2187 ),
    .b(\u2_Display/n2207 [17]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2222 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3549 (
    .a(\u2_Display/n2186 ),
    .b(\u2_Display/n2207 [18]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2221 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u355 (
    .a(\u2_Display/n3788 [24]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [24]),
    .o(\u2_Display/n3796 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3550 (
    .a(\u2_Display/n2185 ),
    .b(\u2_Display/n2207 [19]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2220 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3551 (
    .a(\u2_Display/n2184 ),
    .b(\u2_Display/n2207 [20]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2219 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3552 (
    .a(\u2_Display/n2183 ),
    .b(\u2_Display/n2207 [21]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2218 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3553 (
    .a(\u2_Display/n2182 ),
    .b(\u2_Display/n2207 [22]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2217 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3554 (
    .a(\u2_Display/n2181 ),
    .b(\u2_Display/n2207 [23]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2216 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3555 (
    .a(\u2_Display/n2180 ),
    .b(\u2_Display/n2207 [24]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2215 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3556 (
    .a(\u2_Display/n2179 ),
    .b(\u2_Display/n2207 [25]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2214 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3557 (
    .a(\u2_Display/n2178 ),
    .b(\u2_Display/n2207 [26]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2213 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3558 (
    .a(\u2_Display/n2177 ),
    .b(\u2_Display/n2207 [27]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2212 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3559 (
    .a(\u2_Display/n2176 ),
    .b(\u2_Display/n2207 [28]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2211 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u356 (
    .a(\u2_Display/n3788 [25]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [25]),
    .o(\u2_Display/n3795 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3560 (
    .a(\u2_Display/n2175 ),
    .b(\u2_Display/n2207 [29]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2210 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3561 (
    .a(\u2_Display/n2174 ),
    .b(\u2_Display/n2207 [30]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2209 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3562 (
    .a(\u2_Display/n2173 ),
    .b(\u2_Display/n2207 [31]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2208 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3563 (
    .a(\u2_Display/n3327 ),
    .b(\u2_Display/n3330 [0]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3362 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3564 (
    .a(\u2_Display/n3326 ),
    .b(\u2_Display/n3330 [1]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3361 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3565 (
    .a(\u2_Display/n3325 ),
    .b(\u2_Display/n3330 [2]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3360 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3566 (
    .a(\u2_Display/n3324 ),
    .b(\u2_Display/n3330 [3]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3359 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3567 (
    .a(\u2_Display/n3323 ),
    .b(\u2_Display/n3330 [4]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3358 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3568 (
    .a(\u2_Display/n3322 ),
    .b(\u2_Display/n3330 [5]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3357 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3569 (
    .a(\u2_Display/n3321 ),
    .b(\u2_Display/n3330 [6]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3356 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u357 (
    .a(\u2_Display/n3788 [26]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [26]),
    .o(\u2_Display/n3794 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3570 (
    .a(\u2_Display/n3320 ),
    .b(\u2_Display/n3330 [7]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3355 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3571 (
    .a(\u2_Display/n3319 ),
    .b(\u2_Display/n3330 [8]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3354 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3572 (
    .a(\u2_Display/n3318 ),
    .b(\u2_Display/n3330 [9]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3353 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3573 (
    .a(\u2_Display/n3317 ),
    .b(\u2_Display/n3330 [10]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3352 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3574 (
    .a(\u2_Display/n3316 ),
    .b(\u2_Display/n3330 [11]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3351 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3575 (
    .a(\u2_Display/n3315 ),
    .b(\u2_Display/n3330 [12]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3350 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3576 (
    .a(\u2_Display/n3314 ),
    .b(\u2_Display/n3330 [13]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3349 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3577 (
    .a(\u2_Display/n3313 ),
    .b(\u2_Display/n3330 [14]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3348 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3578 (
    .a(\u2_Display/n3312 ),
    .b(\u2_Display/n3330 [15]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3347 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3579 (
    .a(\u2_Display/n3311 ),
    .b(\u2_Display/n3330 [16]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3346 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u358 (
    .a(\u2_Display/n3788 [27]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [27]),
    .o(\u2_Display/n3793 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3580 (
    .a(\u2_Display/n3310 ),
    .b(\u2_Display/n3330 [17]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3345 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3581 (
    .a(\u2_Display/n3309 ),
    .b(\u2_Display/n3330 [18]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3344 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3582 (
    .a(\u2_Display/n3308 ),
    .b(\u2_Display/n3330 [19]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3343 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3583 (
    .a(\u2_Display/n3307 ),
    .b(\u2_Display/n3330 [20]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3342 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3584 (
    .a(\u2_Display/n3306 ),
    .b(\u2_Display/n3330 [21]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3341 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3585 (
    .a(\u2_Display/n3305 ),
    .b(\u2_Display/n3330 [22]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3340 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3586 (
    .a(\u2_Display/n3304 ),
    .b(\u2_Display/n3330 [23]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3339 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3587 (
    .a(\u2_Display/n3303 ),
    .b(\u2_Display/n3330 [24]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3338 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3588 (
    .a(\u2_Display/n3302 ),
    .b(\u2_Display/n3330 [25]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3337 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3589 (
    .a(\u2_Display/n3301 ),
    .b(\u2_Display/n3330 [26]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3336 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u359 (
    .a(\u2_Display/n3788 [28]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [28]),
    .o(\u2_Display/n3792 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3590 (
    .a(\u2_Display/n3300 ),
    .b(\u2_Display/n3330 [27]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3335 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3591 (
    .a(\u2_Display/n3299 ),
    .b(\u2_Display/n3330 [28]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3334 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3592 (
    .a(\u2_Display/n3298 ),
    .b(\u2_Display/n3330 [29]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3333 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3593 (
    .a(\u2_Display/n3297 ),
    .b(\u2_Display/n3330 [30]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3332 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3594 (
    .a(\u2_Display/n3296 ),
    .b(\u2_Display/n3330 [31]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3331 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3595 (
    .a(\u2_Display/n4485 ),
    .b(\u2_Display/n4488 [0]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4520 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3596 (
    .a(\u2_Display/n4484 ),
    .b(\u2_Display/n4488 [1]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4519 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3597 (
    .a(\u2_Display/n4483 ),
    .b(\u2_Display/n4488 [2]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4518 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3598 (
    .a(\u2_Display/n4482 ),
    .b(\u2_Display/n4488 [3]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4517 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3599 (
    .a(\u2_Display/n4481 ),
    .b(\u2_Display/n4488 [4]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4516 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u360 (
    .a(\u2_Display/n3788 [29]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [29]),
    .o(\u2_Display/n3791 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3600 (
    .a(\u2_Display/n4480 ),
    .b(\u2_Display/n4488 [5]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4515 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3601 (
    .a(\u2_Display/n4479 ),
    .b(\u2_Display/n4488 [6]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4514 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3602 (
    .a(\u2_Display/n4478 ),
    .b(\u2_Display/n4488 [7]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4513 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3603 (
    .a(\u2_Display/n4477 ),
    .b(\u2_Display/n4488 [8]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4512 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3604 (
    .a(\u2_Display/n4476 ),
    .b(\u2_Display/n4488 [9]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4511 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3605 (
    .a(\u2_Display/n4475 ),
    .b(\u2_Display/n4488 [10]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4510 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3606 (
    .a(\u2_Display/n4474 ),
    .b(\u2_Display/n4488 [11]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4509 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3607 (
    .a(\u2_Display/n4473 ),
    .b(\u2_Display/n4488 [12]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4508 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3608 (
    .a(\u2_Display/n4472 ),
    .b(\u2_Display/n4488 [13]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4507 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3609 (
    .a(\u2_Display/n4471 ),
    .b(\u2_Display/n4488 [14]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4506 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u361 (
    .a(\u2_Display/n3788 [30]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [30]),
    .o(\u2_Display/n3790 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3610 (
    .a(\u2_Display/n4470 ),
    .b(\u2_Display/n4488 [15]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4505 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3611 (
    .a(\u2_Display/n4469 ),
    .b(\u2_Display/n4488 [16]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4504 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3612 (
    .a(\u2_Display/n4468 ),
    .b(\u2_Display/n4488 [17]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4503 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3613 (
    .a(\u2_Display/n4467 ),
    .b(\u2_Display/n4488 [18]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4502 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3614 (
    .a(\u2_Display/n4466 ),
    .b(\u2_Display/n4488 [19]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4501 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3615 (
    .a(\u2_Display/n4465 ),
    .b(\u2_Display/n4488 [20]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4500 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3616 (
    .a(\u2_Display/n4464 ),
    .b(\u2_Display/n4488 [21]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4499 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3617 (
    .a(\u2_Display/n4463 ),
    .b(\u2_Display/n4488 [22]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4498 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3618 (
    .a(\u2_Display/n4462 ),
    .b(\u2_Display/n4488 [23]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4497 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3619 (
    .a(\u2_Display/n4461 ),
    .b(\u2_Display/n4488 [24]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4496 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u362 (
    .a(\u2_Display/n3788 [31]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [31]),
    .o(\u2_Display/n3789 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3620 (
    .a(\u2_Display/n4460 ),
    .b(\u2_Display/n4488 [25]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4495 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3621 (
    .a(\u2_Display/n4459 ),
    .b(\u2_Display/n4488 [26]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4494 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3622 (
    .a(\u2_Display/n4458 ),
    .b(\u2_Display/n4488 [27]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4493 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3623 (
    .a(\u2_Display/n4457 ),
    .b(\u2_Display/n4488 [28]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4492 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3624 (
    .a(\u2_Display/n4456 ),
    .b(\u2_Display/n4488 [29]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4491 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3625 (
    .a(\u2_Display/n4455 ),
    .b(\u2_Display/n4488 [30]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4490 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3626 (
    .a(\u2_Display/n4454 ),
    .b(\u2_Display/n4488 [31]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4489 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3627 (
    .a(\u2_Display/n5608 ),
    .b(\u2_Display/n5611 [0]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5643 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3628 (
    .a(\u2_Display/n5607 ),
    .b(\u2_Display/n5611 [1]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5642 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3629 (
    .a(\u2_Display/n5606 ),
    .b(\u2_Display/n5611 [2]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5641 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u363 (
    .a(\u2_Display/n4911 [0]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [0]),
    .o(\u2_Display/n6101 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3630 (
    .a(\u2_Display/n5605 ),
    .b(\u2_Display/n5611 [3]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5640 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3631 (
    .a(\u2_Display/n5604 ),
    .b(\u2_Display/n5611 [4]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5639 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3632 (
    .a(\u2_Display/n5603 ),
    .b(\u2_Display/n5611 [5]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5638 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3633 (
    .a(\u2_Display/n5602 ),
    .b(\u2_Display/n5611 [6]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5637 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3634 (
    .a(\u2_Display/n5601 ),
    .b(\u2_Display/n5611 [7]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5636 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3635 (
    .a(\u2_Display/n5600 ),
    .b(\u2_Display/n5611 [8]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5635 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3636 (
    .a(\u2_Display/n5599 ),
    .b(\u2_Display/n5611 [9]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5634 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3637 (
    .a(\u2_Display/n5598 ),
    .b(\u2_Display/n5611 [10]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5633 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3638 (
    .a(\u2_Display/n5597 ),
    .b(\u2_Display/n5611 [11]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5632 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3639 (
    .a(\u2_Display/n5596 ),
    .b(\u2_Display/n5611 [12]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5631 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u364 (
    .a(\u2_Display/n4911 [1]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [1]),
    .o(\u2_Display/n6100 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3640 (
    .a(\u2_Display/n5595 ),
    .b(\u2_Display/n5611 [13]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5630 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3641 (
    .a(\u2_Display/n5594 ),
    .b(\u2_Display/n5611 [14]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5629 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3642 (
    .a(\u2_Display/n5593 ),
    .b(\u2_Display/n5611 [15]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5628 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3643 (
    .a(\u2_Display/n5592 ),
    .b(\u2_Display/n5611 [16]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5627 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3644 (
    .a(\u2_Display/n5591 ),
    .b(\u2_Display/n5611 [17]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5626 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3645 (
    .a(\u2_Display/n5590 ),
    .b(\u2_Display/n5611 [18]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5625 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3646 (
    .a(\u2_Display/n5589 ),
    .b(\u2_Display/n5611 [19]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5624 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3647 (
    .a(\u2_Display/n5588 ),
    .b(\u2_Display/n5611 [20]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5623 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3648 (
    .a(\u2_Display/n5587 ),
    .b(\u2_Display/n5611 [21]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5622 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3649 (
    .a(\u2_Display/n5586 ),
    .b(\u2_Display/n5611 [22]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5621 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u365 (
    .a(\u2_Display/n4911 [2]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [2]),
    .o(\u2_Display/n6099 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3650 (
    .a(\u2_Display/n5585 ),
    .b(\u2_Display/n5611 [23]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5620 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3651 (
    .a(\u2_Display/n5584 ),
    .b(\u2_Display/n5611 [24]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5619 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3652 (
    .a(\u2_Display/n5583 ),
    .b(\u2_Display/n5611 [25]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5618 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3653 (
    .a(\u2_Display/n5582 ),
    .b(\u2_Display/n5611 [26]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5617 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3654 (
    .a(\u2_Display/n5581 ),
    .b(\u2_Display/n5611 [27]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5616 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3655 (
    .a(\u2_Display/n5580 ),
    .b(\u2_Display/n5611 [28]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5615 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3656 (
    .a(\u2_Display/n5579 ),
    .b(\u2_Display/n5611 [29]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5614 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3657 (
    .a(\u2_Display/n5578 ),
    .b(\u2_Display/n5611 [30]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5613 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3658 (
    .a(\u2_Display/n5577 ),
    .b(\u2_Display/n5611 [31]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5612 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3659 (
    .a(\u2_Display/n1116 ),
    .b(\u2_Display/n1119 [0]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1151 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u366 (
    .a(\u2_Display/n4911 [3]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [3]),
    .o(\u2_Display/n6098 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3660 (
    .a(\u2_Display/n1115 ),
    .b(\u2_Display/n1119 [1]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1150 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3661 (
    .a(\u2_Display/n1114 ),
    .b(\u2_Display/n1119 [2]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1149 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3662 (
    .a(\u2_Display/n1113 ),
    .b(\u2_Display/n1119 [3]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1148 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3663 (
    .a(\u2_Display/n1112 ),
    .b(\u2_Display/n1119 [4]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1147 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3664 (
    .a(\u2_Display/n1111 ),
    .b(\u2_Display/n1119 [5]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1146 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3665 (
    .a(\u2_Display/n1110 ),
    .b(\u2_Display/n1119 [6]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1145 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3666 (
    .a(\u2_Display/n1109 ),
    .b(\u2_Display/n1119 [7]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1144 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3667 (
    .a(\u2_Display/n1108 ),
    .b(\u2_Display/n1119 [8]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1143 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3668 (
    .a(\u2_Display/n1107 ),
    .b(\u2_Display/n1119 [9]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1142 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3669 (
    .a(\u2_Display/n1106 ),
    .b(\u2_Display/n1119 [10]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1141 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u367 (
    .a(\u2_Display/n4911 [4]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [4]),
    .o(\u2_Display/n6097 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3670 (
    .a(\u2_Display/n1105 ),
    .b(\u2_Display/n1119 [11]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1140 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3671 (
    .a(\u2_Display/n1104 ),
    .b(\u2_Display/n1119 [12]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1139 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3672 (
    .a(\u2_Display/n1103 ),
    .b(\u2_Display/n1119 [13]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1138 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3673 (
    .a(\u2_Display/n1102 ),
    .b(\u2_Display/n1119 [14]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1137 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3674 (
    .a(\u2_Display/n1101 ),
    .b(\u2_Display/n1119 [15]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1136 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3675 (
    .a(\u2_Display/n1100 ),
    .b(\u2_Display/n1119 [16]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1135 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3676 (
    .a(\u2_Display/n1099 ),
    .b(\u2_Display/n1119 [17]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1134 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3677 (
    .a(\u2_Display/n1098 ),
    .b(\u2_Display/n1119 [18]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1133 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3678 (
    .a(\u2_Display/n1097 ),
    .b(\u2_Display/n1119 [19]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1132 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3679 (
    .a(\u2_Display/n1096 ),
    .b(\u2_Display/n1119 [20]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1131 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u368 (
    .a(\u2_Display/n4911 [5]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [5]),
    .o(\u2_Display/n6096 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3680 (
    .a(\u2_Display/n1095 ),
    .b(\u2_Display/n1119 [21]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1130 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3681 (
    .a(\u2_Display/n1094 ),
    .b(\u2_Display/n1119 [22]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1129 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3682 (
    .a(\u2_Display/n1093 ),
    .b(\u2_Display/n1119 [23]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1128 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3683 (
    .a(\u2_Display/n1092 ),
    .b(\u2_Display/n1119 [24]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1127 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3684 (
    .a(\u2_Display/n1091 ),
    .b(\u2_Display/n1119 [25]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1126 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3685 (
    .a(\u2_Display/n1090 ),
    .b(\u2_Display/n1119 [26]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1125 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3686 (
    .a(\u2_Display/n1089 ),
    .b(\u2_Display/n1119 [27]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1124 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3687 (
    .a(\u2_Display/n1088 ),
    .b(\u2_Display/n1119 [28]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1123 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3688 (
    .a(\u2_Display/n1087 ),
    .b(\u2_Display/n1119 [29]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1122 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3689 (
    .a(\u2_Display/n1086 ),
    .b(\u2_Display/n1119 [30]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1121 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u369 (
    .a(\u2_Display/n4911 [6]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [6]),
    .o(\u2_Display/n6095 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3690 (
    .a(\u2_Display/n1085 ),
    .b(\u2_Display/n1119 [31]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1120 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3691 (
    .a(\u2_Display/n2239 ),
    .b(\u2_Display/n2242 [0]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2274 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3692 (
    .a(\u2_Display/n2238 ),
    .b(\u2_Display/n2242 [1]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2273 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3693 (
    .a(\u2_Display/n2237 ),
    .b(\u2_Display/n2242 [2]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2272 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3694 (
    .a(\u2_Display/n2236 ),
    .b(\u2_Display/n2242 [3]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2271 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3695 (
    .a(\u2_Display/n2235 ),
    .b(\u2_Display/n2242 [4]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2270 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3696 (
    .a(\u2_Display/n2234 ),
    .b(\u2_Display/n2242 [5]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2269 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3697 (
    .a(\u2_Display/n2233 ),
    .b(\u2_Display/n2242 [6]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2268 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3698 (
    .a(\u2_Display/n2232 ),
    .b(\u2_Display/n2242 [7]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2267 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3699 (
    .a(\u2_Display/n2231 ),
    .b(\u2_Display/n2242 [8]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2266 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u370 (
    .a(\u2_Display/n4911 [7]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [7]),
    .o(\u2_Display/n6094 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3700 (
    .a(\u2_Display/n2230 ),
    .b(\u2_Display/n2242 [9]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2265 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3701 (
    .a(\u2_Display/n2229 ),
    .b(\u2_Display/n2242 [10]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2264 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3702 (
    .a(\u2_Display/n2228 ),
    .b(\u2_Display/n2242 [11]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2263 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3703 (
    .a(\u2_Display/n2227 ),
    .b(\u2_Display/n2242 [12]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2262 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3704 (
    .a(\u2_Display/n2226 ),
    .b(\u2_Display/n2242 [13]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2261 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3705 (
    .a(\u2_Display/n2225 ),
    .b(\u2_Display/n2242 [14]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2260 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3706 (
    .a(\u2_Display/n2224 ),
    .b(\u2_Display/n2242 [15]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2259 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3707 (
    .a(\u2_Display/n2223 ),
    .b(\u2_Display/n2242 [16]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2258 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3708 (
    .a(\u2_Display/n2222 ),
    .b(\u2_Display/n2242 [17]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2257 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3709 (
    .a(\u2_Display/n2221 ),
    .b(\u2_Display/n2242 [18]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2256 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u371 (
    .a(\u2_Display/n4911 [8]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [8]),
    .o(\u2_Display/n6093 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3710 (
    .a(\u2_Display/n2220 ),
    .b(\u2_Display/n2242 [19]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2255 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3711 (
    .a(\u2_Display/n2219 ),
    .b(\u2_Display/n2242 [20]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2254 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3712 (
    .a(\u2_Display/n2218 ),
    .b(\u2_Display/n2242 [21]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2253 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3713 (
    .a(\u2_Display/n2217 ),
    .b(\u2_Display/n2242 [22]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2252 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3714 (
    .a(\u2_Display/n2216 ),
    .b(\u2_Display/n2242 [23]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2251 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3715 (
    .a(\u2_Display/n2215 ),
    .b(\u2_Display/n2242 [24]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2250 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3716 (
    .a(\u2_Display/n2214 ),
    .b(\u2_Display/n2242 [25]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2249 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3717 (
    .a(\u2_Display/n2213 ),
    .b(\u2_Display/n2242 [26]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2248 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3718 (
    .a(\u2_Display/n2212 ),
    .b(\u2_Display/n2242 [27]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2247 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3719 (
    .a(\u2_Display/n2211 ),
    .b(\u2_Display/n2242 [28]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2246 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u372 (
    .a(\u2_Display/n4911 [9]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [9]),
    .o(\u2_Display/n6092 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3720 (
    .a(\u2_Display/n2210 ),
    .b(\u2_Display/n2242 [29]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2245 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3721 (
    .a(\u2_Display/n2209 ),
    .b(\u2_Display/n2242 [30]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2244 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3722 (
    .a(\u2_Display/n2208 ),
    .b(\u2_Display/n2242 [31]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2243 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3723 (
    .a(\u2_Display/n3362 ),
    .b(\u2_Display/n3365 [0]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3397 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3724 (
    .a(\u2_Display/n3361 ),
    .b(\u2_Display/n3365 [1]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3396 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3725 (
    .a(\u2_Display/n3360 ),
    .b(\u2_Display/n3365 [2]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3395 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3726 (
    .a(\u2_Display/n3359 ),
    .b(\u2_Display/n3365 [3]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3394 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3727 (
    .a(\u2_Display/n3358 ),
    .b(\u2_Display/n3365 [4]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3393 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3728 (
    .a(\u2_Display/n3357 ),
    .b(\u2_Display/n3365 [5]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3392 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3729 (
    .a(\u2_Display/n3356 ),
    .b(\u2_Display/n3365 [6]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3391 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u373 (
    .a(\u2_Display/n4911 [10]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [10]),
    .o(\u2_Display/n6091 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3730 (
    .a(\u2_Display/n3355 ),
    .b(\u2_Display/n3365 [7]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3390 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3731 (
    .a(\u2_Display/n3354 ),
    .b(\u2_Display/n3365 [8]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3389 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3732 (
    .a(\u2_Display/n3353 ),
    .b(\u2_Display/n3365 [9]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3388 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3733 (
    .a(\u2_Display/n3352 ),
    .b(\u2_Display/n3365 [10]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3387 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3734 (
    .a(\u2_Display/n3351 ),
    .b(\u2_Display/n3365 [11]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3386 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3735 (
    .a(\u2_Display/n3350 ),
    .b(\u2_Display/n3365 [12]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3385 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3736 (
    .a(\u2_Display/n3349 ),
    .b(\u2_Display/n3365 [13]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3384 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3737 (
    .a(\u2_Display/n3348 ),
    .b(\u2_Display/n3365 [14]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3383 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3738 (
    .a(\u2_Display/n3347 ),
    .b(\u2_Display/n3365 [15]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3382 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3739 (
    .a(\u2_Display/n3346 ),
    .b(\u2_Display/n3365 [16]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3381 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u374 (
    .a(\u2_Display/n4911 [11]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [11]),
    .o(\u2_Display/n6090 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3740 (
    .a(\u2_Display/n3345 ),
    .b(\u2_Display/n3365 [17]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3380 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3741 (
    .a(\u2_Display/n3344 ),
    .b(\u2_Display/n3365 [18]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3379 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3742 (
    .a(\u2_Display/n3343 ),
    .b(\u2_Display/n3365 [19]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3378 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3743 (
    .a(\u2_Display/n3342 ),
    .b(\u2_Display/n3365 [20]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3377 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3744 (
    .a(\u2_Display/n3341 ),
    .b(\u2_Display/n3365 [21]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3376 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3745 (
    .a(\u2_Display/n3340 ),
    .b(\u2_Display/n3365 [22]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3375 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3746 (
    .a(\u2_Display/n3339 ),
    .b(\u2_Display/n3365 [23]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3374 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3747 (
    .a(\u2_Display/n3338 ),
    .b(\u2_Display/n3365 [24]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3373 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3748 (
    .a(\u2_Display/n3337 ),
    .b(\u2_Display/n3365 [25]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3372 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3749 (
    .a(\u2_Display/n3336 ),
    .b(\u2_Display/n3365 [26]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3371 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u375 (
    .a(\u2_Display/n4911 [12]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [12]),
    .o(\u2_Display/n6089 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3750 (
    .a(\u2_Display/n3335 ),
    .b(\u2_Display/n3365 [27]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3370 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3751 (
    .a(\u2_Display/n3334 ),
    .b(\u2_Display/n3365 [28]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3369 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3752 (
    .a(\u2_Display/n3333 ),
    .b(\u2_Display/n3365 [29]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3368 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3753 (
    .a(\u2_Display/n3332 ),
    .b(\u2_Display/n3365 [30]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3367 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3754 (
    .a(\u2_Display/n3331 ),
    .b(\u2_Display/n3365 [31]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3366 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3755 (
    .a(\u2_Display/n4520 ),
    .b(\u2_Display/n4523 [0]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4555 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3756 (
    .a(\u2_Display/n4519 ),
    .b(\u2_Display/n4523 [1]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4554 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3757 (
    .a(\u2_Display/n4518 ),
    .b(\u2_Display/n4523 [2]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4553 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3758 (
    .a(\u2_Display/n4517 ),
    .b(\u2_Display/n4523 [3]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4552 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3759 (
    .a(\u2_Display/n4516 ),
    .b(\u2_Display/n4523 [4]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4551 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u376 (
    .a(\u2_Display/n4911 [13]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [13]),
    .o(\u2_Display/n6088 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3760 (
    .a(\u2_Display/n4515 ),
    .b(\u2_Display/n4523 [5]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4550 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3761 (
    .a(\u2_Display/n4514 ),
    .b(\u2_Display/n4523 [6]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4549 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3762 (
    .a(\u2_Display/n4513 ),
    .b(\u2_Display/n4523 [7]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4548 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3763 (
    .a(\u2_Display/n4512 ),
    .b(\u2_Display/n4523 [8]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4547 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3764 (
    .a(\u2_Display/n4511 ),
    .b(\u2_Display/n4523 [9]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4546 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3765 (
    .a(\u2_Display/n4510 ),
    .b(\u2_Display/n4523 [10]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4545 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3766 (
    .a(\u2_Display/n4509 ),
    .b(\u2_Display/n4523 [11]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4544 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3767 (
    .a(\u2_Display/n4508 ),
    .b(\u2_Display/n4523 [12]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4543 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3768 (
    .a(\u2_Display/n4507 ),
    .b(\u2_Display/n4523 [13]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4542 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3769 (
    .a(\u2_Display/n4506 ),
    .b(\u2_Display/n4523 [14]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4541 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u377 (
    .a(\u2_Display/n4911 [14]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [14]),
    .o(\u2_Display/n6087 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3770 (
    .a(\u2_Display/n4505 ),
    .b(\u2_Display/n4523 [15]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4540 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3771 (
    .a(\u2_Display/n4504 ),
    .b(\u2_Display/n4523 [16]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4539 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3772 (
    .a(\u2_Display/n4503 ),
    .b(\u2_Display/n4523 [17]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4538 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3773 (
    .a(\u2_Display/n4502 ),
    .b(\u2_Display/n4523 [18]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4537 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3774 (
    .a(\u2_Display/n4501 ),
    .b(\u2_Display/n4523 [19]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4536 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3775 (
    .a(\u2_Display/n4500 ),
    .b(\u2_Display/n4523 [20]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4535 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3776 (
    .a(\u2_Display/n4499 ),
    .b(\u2_Display/n4523 [21]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4534 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3777 (
    .a(\u2_Display/n4498 ),
    .b(\u2_Display/n4523 [22]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4533 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3778 (
    .a(\u2_Display/n4497 ),
    .b(\u2_Display/n4523 [23]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4532 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3779 (
    .a(\u2_Display/n4496 ),
    .b(\u2_Display/n4523 [24]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4531 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u378 (
    .a(\u2_Display/n4911 [15]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [15]),
    .o(\u2_Display/n6086 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3780 (
    .a(\u2_Display/n4495 ),
    .b(\u2_Display/n4523 [25]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4530 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3781 (
    .a(\u2_Display/n4494 ),
    .b(\u2_Display/n4523 [26]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4529 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3782 (
    .a(\u2_Display/n4493 ),
    .b(\u2_Display/n4523 [27]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4528 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3783 (
    .a(\u2_Display/n4492 ),
    .b(\u2_Display/n4523 [28]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4527 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3784 (
    .a(\u2_Display/n4491 ),
    .b(\u2_Display/n4523 [29]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4526 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3785 (
    .a(\u2_Display/n4490 ),
    .b(\u2_Display/n4523 [30]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4525 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3786 (
    .a(\u2_Display/n4489 ),
    .b(\u2_Display/n4523 [31]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4524 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3787 (
    .a(\u2_Display/n5643 ),
    .b(\u2_Display/n5646 [0]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5678 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3788 (
    .a(\u2_Display/n5642 ),
    .b(\u2_Display/n5646 [1]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5677 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3789 (
    .a(\u2_Display/n5641 ),
    .b(\u2_Display/n5646 [2]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5676 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u379 (
    .a(\u2_Display/n4911 [16]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [16]),
    .o(\u2_Display/n6085 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3790 (
    .a(\u2_Display/n5640 ),
    .b(\u2_Display/n5646 [3]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5675 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3791 (
    .a(\u2_Display/n5639 ),
    .b(\u2_Display/n5646 [4]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5674 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3792 (
    .a(\u2_Display/n5638 ),
    .b(\u2_Display/n5646 [5]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5673 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3793 (
    .a(\u2_Display/n5637 ),
    .b(\u2_Display/n5646 [6]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5672 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3794 (
    .a(\u2_Display/n5636 ),
    .b(\u2_Display/n5646 [7]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5671 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3795 (
    .a(\u2_Display/n5635 ),
    .b(\u2_Display/n5646 [8]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5670 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3796 (
    .a(\u2_Display/n5634 ),
    .b(\u2_Display/n5646 [9]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5669 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3797 (
    .a(\u2_Display/n5633 ),
    .b(\u2_Display/n5646 [10]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5668 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3798 (
    .a(\u2_Display/n5632 ),
    .b(\u2_Display/n5646 [11]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5667 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3799 (
    .a(\u2_Display/n5631 ),
    .b(\u2_Display/n5646 [12]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5666 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u380 (
    .a(\u2_Display/n4911 [17]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [17]),
    .o(\u2_Display/n6084 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3800 (
    .a(\u2_Display/n5630 ),
    .b(\u2_Display/n5646 [13]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5665 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3801 (
    .a(\u2_Display/n5629 ),
    .b(\u2_Display/n5646 [14]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5664 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3802 (
    .a(\u2_Display/n5628 ),
    .b(\u2_Display/n5646 [15]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5663 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3803 (
    .a(\u2_Display/n5627 ),
    .b(\u2_Display/n5646 [16]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5662 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3804 (
    .a(\u2_Display/n5626 ),
    .b(\u2_Display/n5646 [17]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5661 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3805 (
    .a(\u2_Display/n5625 ),
    .b(\u2_Display/n5646 [18]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5660 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3806 (
    .a(\u2_Display/n5624 ),
    .b(\u2_Display/n5646 [19]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5659 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3807 (
    .a(\u2_Display/n5623 ),
    .b(\u2_Display/n5646 [20]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5658 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3808 (
    .a(\u2_Display/n5622 ),
    .b(\u2_Display/n5646 [21]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5657 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3809 (
    .a(\u2_Display/n5621 ),
    .b(\u2_Display/n5646 [22]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5656 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u381 (
    .a(\u2_Display/n4911 [18]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [18]),
    .o(\u2_Display/n6083 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3810 (
    .a(\u2_Display/n5620 ),
    .b(\u2_Display/n5646 [23]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5655 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3811 (
    .a(\u2_Display/n5619 ),
    .b(\u2_Display/n5646 [24]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5654 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3812 (
    .a(\u2_Display/n5618 ),
    .b(\u2_Display/n5646 [25]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5653 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3813 (
    .a(\u2_Display/n5617 ),
    .b(\u2_Display/n5646 [26]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5652 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3814 (
    .a(\u2_Display/n5616 ),
    .b(\u2_Display/n5646 [27]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5651 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3815 (
    .a(\u2_Display/n5615 ),
    .b(\u2_Display/n5646 [28]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5650 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3816 (
    .a(\u2_Display/n5614 ),
    .b(\u2_Display/n5646 [29]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5649 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3817 (
    .a(\u2_Display/n5613 ),
    .b(\u2_Display/n5646 [30]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5648 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3818 (
    .a(\u2_Display/n5612 ),
    .b(\u2_Display/n5646 [31]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5647 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3819 (
    .a(\u2_Display/n1151 ),
    .b(\u2_Display/n1154 [0]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1186 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u382 (
    .a(\u2_Display/n4911 [19]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [19]),
    .o(\u2_Display/n6082 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3820 (
    .a(\u2_Display/n1150 ),
    .b(\u2_Display/n1154 [1]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1185 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3821 (
    .a(\u2_Display/n1149 ),
    .b(\u2_Display/n1154 [2]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1184 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3822 (
    .a(\u2_Display/n1148 ),
    .b(\u2_Display/n1154 [3]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1183 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3823 (
    .a(\u2_Display/n1147 ),
    .b(\u2_Display/n1154 [4]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1182 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3824 (
    .a(\u2_Display/n1146 ),
    .b(\u2_Display/n1154 [5]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1181 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3825 (
    .a(\u2_Display/n1145 ),
    .b(\u2_Display/n1154 [6]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1180 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3826 (
    .a(\u2_Display/n1144 ),
    .b(\u2_Display/n1154 [7]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1179 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3827 (
    .a(\u2_Display/n1143 ),
    .b(\u2_Display/n1154 [8]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1178 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3828 (
    .a(\u2_Display/n1142 ),
    .b(\u2_Display/n1154 [9]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1177 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3829 (
    .a(\u2_Display/n1141 ),
    .b(\u2_Display/n1154 [10]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1176 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u383 (
    .a(\u2_Display/n4911 [20]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [20]),
    .o(\u2_Display/n6081 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3830 (
    .a(\u2_Display/n1140 ),
    .b(\u2_Display/n1154 [11]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1175 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3831 (
    .a(\u2_Display/n1139 ),
    .b(\u2_Display/n1154 [12]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1174 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3832 (
    .a(\u2_Display/n1138 ),
    .b(\u2_Display/n1154 [13]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1173 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3833 (
    .a(\u2_Display/n1137 ),
    .b(\u2_Display/n1154 [14]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1172 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3834 (
    .a(\u2_Display/n1136 ),
    .b(\u2_Display/n1154 [15]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1171 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3835 (
    .a(\u2_Display/n1135 ),
    .b(\u2_Display/n1154 [16]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1170 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3836 (
    .a(\u2_Display/n1134 ),
    .b(\u2_Display/n1154 [17]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1169 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3837 (
    .a(\u2_Display/n1133 ),
    .b(\u2_Display/n1154 [18]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1168 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3838 (
    .a(\u2_Display/n1132 ),
    .b(\u2_Display/n1154 [19]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1167 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3839 (
    .a(\u2_Display/n1131 ),
    .b(\u2_Display/n1154 [20]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1166 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u384 (
    .a(\u2_Display/n4911 [21]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [21]),
    .o(\u2_Display/n6080 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3840 (
    .a(\u2_Display/n1130 ),
    .b(\u2_Display/n1154 [21]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1165 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3841 (
    .a(\u2_Display/n1129 ),
    .b(\u2_Display/n1154 [22]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1164 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3842 (
    .a(\u2_Display/n1128 ),
    .b(\u2_Display/n1154 [23]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1163 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3843 (
    .a(\u2_Display/n1127 ),
    .b(\u2_Display/n1154 [24]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1162 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3844 (
    .a(\u2_Display/n1126 ),
    .b(\u2_Display/n1154 [25]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1161 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3845 (
    .a(\u2_Display/n1125 ),
    .b(\u2_Display/n1154 [26]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1160 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3846 (
    .a(\u2_Display/n1124 ),
    .b(\u2_Display/n1154 [27]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1159 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3847 (
    .a(\u2_Display/n1123 ),
    .b(\u2_Display/n1154 [28]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1158 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3848 (
    .a(\u2_Display/n1122 ),
    .b(\u2_Display/n1154 [29]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1157 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3849 (
    .a(\u2_Display/n1121 ),
    .b(\u2_Display/n1154 [30]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1156 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u385 (
    .a(\u2_Display/n4911 [22]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [22]),
    .o(\u2_Display/n6079 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3850 (
    .a(\u2_Display/n1120 ),
    .b(\u2_Display/n1154 [31]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1155 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3851 (
    .a(\u2_Display/n2274 ),
    .b(\u2_Display/n2277 [0]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2309 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3852 (
    .a(\u2_Display/n2273 ),
    .b(\u2_Display/n2277 [1]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2308 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3853 (
    .a(\u2_Display/n2272 ),
    .b(\u2_Display/n2277 [2]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2307 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3854 (
    .a(\u2_Display/n2271 ),
    .b(\u2_Display/n2277 [3]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2306 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3855 (
    .a(\u2_Display/n2270 ),
    .b(\u2_Display/n2277 [4]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2305 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3856 (
    .a(\u2_Display/n2269 ),
    .b(\u2_Display/n2277 [5]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2304 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3857 (
    .a(\u2_Display/n2268 ),
    .b(\u2_Display/n2277 [6]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2303 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3858 (
    .a(\u2_Display/n2267 ),
    .b(\u2_Display/n2277 [7]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2302 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3859 (
    .a(\u2_Display/n2266 ),
    .b(\u2_Display/n2277 [8]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2301 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u386 (
    .a(\u2_Display/n4911 [23]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [23]),
    .o(\u2_Display/n6078 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3860 (
    .a(\u2_Display/n2265 ),
    .b(\u2_Display/n2277 [9]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2300 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3861 (
    .a(\u2_Display/n2264 ),
    .b(\u2_Display/n2277 [10]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2299 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3862 (
    .a(\u2_Display/n2263 ),
    .b(\u2_Display/n2277 [11]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2298 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3863 (
    .a(\u2_Display/n2262 ),
    .b(\u2_Display/n2277 [12]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2297 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3864 (
    .a(\u2_Display/n2261 ),
    .b(\u2_Display/n2277 [13]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2296 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3865 (
    .a(\u2_Display/n2260 ),
    .b(\u2_Display/n2277 [14]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2295 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3866 (
    .a(\u2_Display/n2259 ),
    .b(\u2_Display/n2277 [15]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2294 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3867 (
    .a(\u2_Display/n2258 ),
    .b(\u2_Display/n2277 [16]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2293 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3868 (
    .a(\u2_Display/n2257 ),
    .b(\u2_Display/n2277 [17]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2292 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3869 (
    .a(\u2_Display/n2256 ),
    .b(\u2_Display/n2277 [18]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2291 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u387 (
    .a(\u2_Display/n4911 [24]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [24]),
    .o(\u2_Display/n6077 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3870 (
    .a(\u2_Display/n2255 ),
    .b(\u2_Display/n2277 [19]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2290 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3871 (
    .a(\u2_Display/n2254 ),
    .b(\u2_Display/n2277 [20]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2289 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3872 (
    .a(\u2_Display/n2253 ),
    .b(\u2_Display/n2277 [21]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2288 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3873 (
    .a(\u2_Display/n2252 ),
    .b(\u2_Display/n2277 [22]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2287 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3874 (
    .a(\u2_Display/n2251 ),
    .b(\u2_Display/n2277 [23]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2286 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3875 (
    .a(\u2_Display/n2250 ),
    .b(\u2_Display/n2277 [24]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2285 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3876 (
    .a(\u2_Display/n2249 ),
    .b(\u2_Display/n2277 [25]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2284 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3877 (
    .a(\u2_Display/n2248 ),
    .b(\u2_Display/n2277 [26]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2283 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3878 (
    .a(\u2_Display/n2247 ),
    .b(\u2_Display/n2277 [27]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2282 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3879 (
    .a(\u2_Display/n2246 ),
    .b(\u2_Display/n2277 [28]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2281 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u388 (
    .a(\u2_Display/n4911 [25]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [25]),
    .o(\u2_Display/n6076 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3880 (
    .a(\u2_Display/n2245 ),
    .b(\u2_Display/n2277 [29]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2280 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3881 (
    .a(\u2_Display/n2244 ),
    .b(\u2_Display/n2277 [30]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2279 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3882 (
    .a(\u2_Display/n2243 ),
    .b(\u2_Display/n2277 [31]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2278 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3883 (
    .a(\u2_Display/n3397 ),
    .b(\u2_Display/n3400 [0]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3432 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3884 (
    .a(\u2_Display/n3396 ),
    .b(\u2_Display/n3400 [1]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3431 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3885 (
    .a(\u2_Display/n3395 ),
    .b(\u2_Display/n3400 [2]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3430 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3886 (
    .a(\u2_Display/n3394 ),
    .b(\u2_Display/n3400 [3]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3429 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3887 (
    .a(\u2_Display/n3393 ),
    .b(\u2_Display/n3400 [4]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3428 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3888 (
    .a(\u2_Display/n3392 ),
    .b(\u2_Display/n3400 [5]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3427 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3889 (
    .a(\u2_Display/n3391 ),
    .b(\u2_Display/n3400 [6]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3426 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u389 (
    .a(\u2_Display/n4911 [26]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [26]),
    .o(\u2_Display/n6075 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3890 (
    .a(\u2_Display/n3390 ),
    .b(\u2_Display/n3400 [7]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3425 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3891 (
    .a(\u2_Display/n3389 ),
    .b(\u2_Display/n3400 [8]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3424 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3892 (
    .a(\u2_Display/n3388 ),
    .b(\u2_Display/n3400 [9]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3423 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3893 (
    .a(\u2_Display/n3387 ),
    .b(\u2_Display/n3400 [10]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3422 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3894 (
    .a(\u2_Display/n3386 ),
    .b(\u2_Display/n3400 [11]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3421 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3895 (
    .a(\u2_Display/n3385 ),
    .b(\u2_Display/n3400 [12]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3420 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3896 (
    .a(\u2_Display/n3384 ),
    .b(\u2_Display/n3400 [13]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3419 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3897 (
    .a(\u2_Display/n3383 ),
    .b(\u2_Display/n3400 [14]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3418 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3898 (
    .a(\u2_Display/n3382 ),
    .b(\u2_Display/n3400 [15]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3417 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3899 (
    .a(\u2_Display/n3381 ),
    .b(\u2_Display/n3400 [16]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3416 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u390 (
    .a(\u2_Display/n4911 [27]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [27]),
    .o(\u2_Display/n6074 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3900 (
    .a(\u2_Display/n3380 ),
    .b(\u2_Display/n3400 [17]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3415 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3901 (
    .a(\u2_Display/n3379 ),
    .b(\u2_Display/n3400 [18]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3414 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3902 (
    .a(\u2_Display/n3378 ),
    .b(\u2_Display/n3400 [19]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3413 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3903 (
    .a(\u2_Display/n3377 ),
    .b(\u2_Display/n3400 [20]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3412 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3904 (
    .a(\u2_Display/n3376 ),
    .b(\u2_Display/n3400 [21]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3411 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3905 (
    .a(\u2_Display/n3375 ),
    .b(\u2_Display/n3400 [22]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3410 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3906 (
    .a(\u2_Display/n3374 ),
    .b(\u2_Display/n3400 [23]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3409 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3907 (
    .a(\u2_Display/n3373 ),
    .b(\u2_Display/n3400 [24]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3408 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3908 (
    .a(\u2_Display/n3372 ),
    .b(\u2_Display/n3400 [25]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3407 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3909 (
    .a(\u2_Display/n3371 ),
    .b(\u2_Display/n3400 [26]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3406 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u391 (
    .a(\u2_Display/n4911 [28]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [28]),
    .o(\u2_Display/n6073 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3910 (
    .a(\u2_Display/n3370 ),
    .b(\u2_Display/n3400 [27]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3405 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3911 (
    .a(\u2_Display/n3369 ),
    .b(\u2_Display/n3400 [28]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3404 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3912 (
    .a(\u2_Display/n3368 ),
    .b(\u2_Display/n3400 [29]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3403 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3913 (
    .a(\u2_Display/n3367 ),
    .b(\u2_Display/n3400 [30]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3402 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3914 (
    .a(\u2_Display/n3366 ),
    .b(\u2_Display/n3400 [31]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3401 ));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u3915 (
    .a(\u2_Display/n5668 ),
    .b(_al_u1168_o),
    .c(on_off_pad[0]),
    .d(\u2_Display/i [10]),
    .o(\u2_Display/n238 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3916 (
    .a(\u2_Display/n3432 ),
    .b(\u2_Display/n3435 [0]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3916_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3917 (
    .a(\u2_Display/n1186 ),
    .b(\u2_Display/n1189 [0]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3917_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3918 (
    .a(_al_u3916_o),
    .b(_al_u3917_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [0]),
    .o(_al_u3918_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3919 (
    .a(_al_u3918_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [0]),
    .o(\u2_Display/n239 [0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u392 (
    .a(\u2_Display/n4911 [29]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [29]),
    .o(\u2_Display/n6072 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3920 (
    .a(\u2_Display/n3431 ),
    .b(\u2_Display/n3435 [1]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3920_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3921 (
    .a(\u2_Display/n1185 ),
    .b(\u2_Display/n1189 [1]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3921_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3922 (
    .a(_al_u3920_o),
    .b(_al_u3921_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [1]),
    .o(_al_u3922_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3923 (
    .a(_al_u3922_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [1]),
    .o(\u2_Display/n239 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3924 (
    .a(\u2_Display/n1184 ),
    .b(\u2_Display/n1189 [2]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3924_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3925 (
    .a(\u2_Display/n3430 ),
    .b(\u2_Display/n3435 [2]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3925_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~((E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D))*~(C)+B*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*~(C)+~(B)*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*C+B*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*C)"),
    .INIT(32'hacfcac0c))
    _al_u3926 (
    .a(_al_u3924_o),
    .b(_al_u3925_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [2]),
    .o(_al_u3926_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u3927 (
    .a(_al_u3926_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [2]),
    .o(\u2_Display/n239 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3928 (
    .a(\u2_Display/n3429 ),
    .b(\u2_Display/n3435 [3]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3928_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3929 (
    .a(\u2_Display/n1183 ),
    .b(\u2_Display/n1189 [3]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3929_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u393 (
    .a(\u2_Display/n4911 [30]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [30]),
    .o(\u2_Display/n6071 ));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3930 (
    .a(_al_u3928_o),
    .b(_al_u3929_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [3]),
    .o(_al_u3930_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3931 (
    .a(_al_u3930_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [3]),
    .o(\u2_Display/n239 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3932 (
    .a(\u2_Display/n3428 ),
    .b(\u2_Display/n3435 [4]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3932_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3933 (
    .a(\u2_Display/n1182 ),
    .b(\u2_Display/n1189 [4]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3933_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3934 (
    .a(_al_u3932_o),
    .b(_al_u3933_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [4]),
    .o(_al_u3934_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3935 (
    .a(_al_u3934_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [4]),
    .o(\u2_Display/n239 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3936 (
    .a(\u2_Display/n3427 ),
    .b(\u2_Display/n3435 [5]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3936_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3937 (
    .a(\u2_Display/n1181 ),
    .b(\u2_Display/n1189 [5]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3937_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3938 (
    .a(_al_u3936_o),
    .b(_al_u3937_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [5]),
    .o(_al_u3938_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3939 (
    .a(_al_u3938_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [5]),
    .o(\u2_Display/n239 [5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u394 (
    .a(\u2_Display/n4911 [31]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [31]),
    .o(\u2_Display/n6070 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3940 (
    .a(\u2_Display/n1180 ),
    .b(\u2_Display/n1189 [6]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3940_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3941 (
    .a(\u2_Display/n3426 ),
    .b(\u2_Display/n3435 [6]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3941_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~((E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D))*~(C)+B*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*~(C)+~(B)*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*C+B*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*C)"),
    .INIT(32'hacfcac0c))
    _al_u3942 (
    .a(_al_u3940_o),
    .b(_al_u3941_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [6]),
    .o(_al_u3942_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u3943 (
    .a(_al_u3942_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [6]),
    .o(\u2_Display/n239 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3944 (
    .a(\u2_Display/n3425 ),
    .b(\u2_Display/n3435 [7]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3944_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3945 (
    .a(\u2_Display/n1179 ),
    .b(\u2_Display/n1189 [7]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3945_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3946 (
    .a(_al_u3944_o),
    .b(_al_u3945_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [7]),
    .o(_al_u3946_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3947 (
    .a(_al_u3946_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [7]),
    .o(\u2_Display/n239 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3948 (
    .a(\u2_Display/n1178 ),
    .b(\u2_Display/n1189 [8]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3948_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3949 (
    .a(\u2_Display/n3424 ),
    .b(\u2_Display/n3435 [8]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3949_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u395 (
    .a(\u2_Display/n419 [0]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [0]),
    .o(\u2_Display/n451 ));
  AL_MAP_LUT5 #(
    .EQN("(B*~((E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D))*~(C)+B*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*~(C)+~(B)*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*C+B*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*C)"),
    .INIT(32'hacfcac0c))
    _al_u3950 (
    .a(_al_u3948_o),
    .b(_al_u3949_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [8]),
    .o(_al_u3950_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u3951 (
    .a(_al_u3950_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [8]),
    .o(\u2_Display/n239 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3952 (
    .a(\u2_Display/n3423 ),
    .b(\u2_Display/n3435 [9]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3952_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3953 (
    .a(\u2_Display/n1177 ),
    .b(\u2_Display/n1189 [9]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3953_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3954 (
    .a(_al_u3952_o),
    .b(_al_u3953_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [9]),
    .o(_al_u3954_o));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    _al_u3955 (
    .a(_al_u3954_o),
    .b(on_off_pad[1]),
    .c(on_off_pad[0]),
    .d(\u2_Display/counta [9]),
    .o(\u2_Display/n239 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .INIT(16'haab8))
    _al_u3956 (
    .a(\u2_Display/n5678 ),
    .b(on_off_pad[0]),
    .c(\u2_Display/n5681 [0]),
    .d(\u2_Display/n5679 ),
    .o(_al_u3956_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3957 (
    .a(\u2_Display/n2309 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [0]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [0]),
    .o(_al_u3957_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*~(C)+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(C)+~(~A)*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C)"),
    .INIT(32'h3a3a0afa))
    _al_u3958 (
    .a(_al_u3957_o),
    .b(\u2_Display/n4555 ),
    .c(on_off_pad[2]),
    .d(\u2_Display/n4558 [0]),
    .e(\u2_Display/n4556 ),
    .o(_al_u3958_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u3959 (
    .a(_al_u3958_o),
    .b(_al_u3956_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u396 (
    .a(\u2_Display/n419 [1]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [1]),
    .o(\u2_Display/n450 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3960 (
    .a(\u2_Display/n2308 ),
    .b(\u2_Display/n2312 [1]),
    .c(\u2_Display/n2310 ),
    .o(_al_u3960_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3961 (
    .a(\u2_Display/n4554 ),
    .b(\u2_Display/n4558 [1]),
    .c(\u2_Display/n4556 ),
    .o(_al_u3961_o));
  AL_MAP_LUT5 #(
    .EQN("~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'h330533f5))
    _al_u3962 (
    .a(_al_u3960_o),
    .b(_al_u3961_o),
    .c(\u2_Display/mux5_b0_sel_is_0_o ),
    .d(on_off_pad[2]),
    .e(\u2_Display/i [1]),
    .o(_al_u3962_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h5757535f))
    _al_u3963 (
    .a(\u2_Display/n5677 ),
    .b(on_off_pad[1]),
    .c(on_off_pad[0]),
    .d(\u2_Display/n5681 [1]),
    .e(\u2_Display/n5679 ),
    .o(_al_u3963_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u3964 (
    .a(_al_u3962_o),
    .b(_al_u3963_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .INIT(16'haab8))
    _al_u3965 (
    .a(\u2_Display/n5676 ),
    .b(on_off_pad[0]),
    .c(\u2_Display/n5681 [2]),
    .d(\u2_Display/n5679 ),
    .o(_al_u3965_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3966 (
    .a(\u2_Display/n2307 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [2]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [2]),
    .o(_al_u3966_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*~(C)+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(C)+~(~A)*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C)"),
    .INIT(32'h3a3a0afa))
    _al_u3967 (
    .a(_al_u3966_o),
    .b(\u2_Display/n4553 ),
    .c(on_off_pad[2]),
    .d(\u2_Display/n4558 [2]),
    .e(\u2_Display/n4556 ),
    .o(_al_u3967_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u3968 (
    .a(_al_u3967_o),
    .b(_al_u3965_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3969 (
    .a(\u2_Display/n2306 ),
    .b(\u2_Display/n2312 [3]),
    .c(\u2_Display/n2310 ),
    .o(_al_u3969_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u397 (
    .a(\u2_Display/n419 [2]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [2]),
    .o(\u2_Display/n449 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3970 (
    .a(\u2_Display/n4552 ),
    .b(\u2_Display/n4558 [3]),
    .c(\u2_Display/n4556 ),
    .o(_al_u3970_o));
  AL_MAP_LUT5 #(
    .EQN("~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'h330533f5))
    _al_u3971 (
    .a(_al_u3969_o),
    .b(_al_u3970_o),
    .c(\u2_Display/mux5_b0_sel_is_0_o ),
    .d(on_off_pad[2]),
    .e(\u2_Display/i [3]),
    .o(_al_u3971_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h5757535f))
    _al_u3972 (
    .a(\u2_Display/n5675 ),
    .b(on_off_pad[1]),
    .c(on_off_pad[0]),
    .d(\u2_Display/n5681 [3]),
    .e(\u2_Display/n5679 ),
    .o(_al_u3972_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u3973 (
    .a(_al_u3971_o),
    .b(_al_u3972_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3974 (
    .a(\u2_Display/n4551 ),
    .b(\u2_Display/n4558 [4]),
    .c(\u2_Display/n4556 ),
    .o(_al_u3974_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3975 (
    .a(\u2_Display/n2305 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [4]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [4]),
    .o(_al_u3975_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h5757535f))
    _al_u3976 (
    .a(\u2_Display/n5674 ),
    .b(on_off_pad[1]),
    .c(on_off_pad[0]),
    .d(\u2_Display/n5681 [4]),
    .e(\u2_Display/n5679 ),
    .o(_al_u3976_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*(~B*~(A)*~(E)+~B*A*~(E)+~(~B)*A*E+~B*A*E)))"),
    .INIT(32'haf0f3f0f))
    _al_u3977 (
    .a(_al_u3974_o),
    .b(_al_u3975_o),
    .c(_al_u3976_o),
    .d(\u2_Display/mux19_b0_sel_is_0_o ),
    .e(on_off_pad[2]),
    .o(\u2_Display/n238 [4]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hababafa3))
    _al_u3978 (
    .a(\u2_Display/n5673 ),
    .b(on_off_pad[1]),
    .c(on_off_pad[0]),
    .d(\u2_Display/n5681 [5]),
    .e(\u2_Display/n5679 ),
    .o(_al_u3978_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3979 (
    .a(\u2_Display/n2304 ),
    .b(\u2_Display/n2312 [5]),
    .c(\u2_Display/n2310 ),
    .o(_al_u3979_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u398 (
    .a(\u2_Display/n419 [3]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [3]),
    .o(\u2_Display/n448 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u3980 (
    .a(_al_u3979_o),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(on_off_pad[2]),
    .d(\u2_Display/i [5]),
    .o(_al_u3980_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    .INIT(16'h88c0))
    _al_u3981 (
    .a(\u2_Display/n4550 ),
    .b(on_off_pad[2]),
    .c(\u2_Display/n4558 [5]),
    .d(\u2_Display/n4556 ),
    .o(_al_u3981_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u3982 (
    .a(_al_u3980_o),
    .b(_al_u3978_o),
    .c(_al_u3981_o),
    .d(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3983 (
    .a(\u2_Display/n4549 ),
    .b(\u2_Display/n4558 [6]),
    .c(\u2_Display/n4556 ),
    .o(_al_u3983_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3984 (
    .a(\u2_Display/n2303 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [6]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [6]),
    .o(_al_u3984_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h5757535f))
    _al_u3985 (
    .a(\u2_Display/n5672 ),
    .b(on_off_pad[1]),
    .c(on_off_pad[0]),
    .d(\u2_Display/n5681 [6]),
    .e(\u2_Display/n5679 ),
    .o(_al_u3985_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*(~B*~(A)*~(E)+~B*A*~(E)+~(~B)*A*E+~B*A*E)))"),
    .INIT(32'haf0f3f0f))
    _al_u3986 (
    .a(_al_u3983_o),
    .b(_al_u3984_o),
    .c(_al_u3985_o),
    .d(\u2_Display/mux19_b0_sel_is_0_o ),
    .e(on_off_pad[2]),
    .o(\u2_Display/n238 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .INIT(16'haab8))
    _al_u3987 (
    .a(\u2_Display/n5671 ),
    .b(on_off_pad[0]),
    .c(\u2_Display/n5681 [7]),
    .d(\u2_Display/n5679 ),
    .o(_al_u3987_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3988 (
    .a(\u2_Display/n2302 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [7]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [7]),
    .o(_al_u3988_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*~(C)+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(C)+~(~A)*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C)"),
    .INIT(32'h3a3a0afa))
    _al_u3989 (
    .a(_al_u3988_o),
    .b(\u2_Display/n4548 ),
    .c(on_off_pad[2]),
    .d(\u2_Display/n4558 [7]),
    .e(\u2_Display/n4556 ),
    .o(_al_u3989_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u399 (
    .a(\u2_Display/n419 [4]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [4]),
    .o(\u2_Display/n447 ));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u3990 (
    .a(_al_u3989_o),
    .b(_al_u3987_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .INIT(16'haab8))
    _al_u3991 (
    .a(\u2_Display/n5670 ),
    .b(on_off_pad[0]),
    .c(\u2_Display/n5681 [8]),
    .d(\u2_Display/n5679 ),
    .o(_al_u3991_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3992 (
    .a(\u2_Display/n2301 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [8]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [8]),
    .o(_al_u3992_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*~(C)+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(C)+~(~A)*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C)"),
    .INIT(32'h3a3a0afa))
    _al_u3993 (
    .a(_al_u3992_o),
    .b(\u2_Display/n4547 ),
    .c(on_off_pad[2]),
    .d(\u2_Display/n4558 [8]),
    .e(\u2_Display/n4556 ),
    .o(_al_u3993_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u3994 (
    .a(_al_u3993_o),
    .b(_al_u3991_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .INIT(16'haab8))
    _al_u3995 (
    .a(\u2_Display/n5669 ),
    .b(on_off_pad[0]),
    .c(\u2_Display/n5681 [9]),
    .d(\u2_Display/n5679 ),
    .o(_al_u3995_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3996 (
    .a(\u2_Display/n2300 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [9]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [9]),
    .o(_al_u3996_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*~(C)+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(C)+~(~A)*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C)"),
    .INIT(32'h3a3a0afa))
    _al_u3997 (
    .a(_al_u3996_o),
    .b(\u2_Display/n4546 ),
    .c(on_off_pad[2]),
    .d(\u2_Display/n4558 [9]),
    .e(\u2_Display/n4556 ),
    .o(_al_u3997_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u3998 (
    .a(_al_u3997_o),
    .b(_al_u3995_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [9]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u3999 (
    .a(rst_n_pad),
    .o(\u0_PLL/n0 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u400 (
    .a(\u2_Display/n419 [5]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [5]),
    .o(\u2_Display/n446 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u4000 (
    .a(clk_vga),
    .o(vga_clk_pad));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u4001 (
    .a(\u1_Driver/n4 ),
    .o(vga_hs_pad));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u4002 (
    .a(\u1_Driver/n10 ),
    .o(vga_vs_pad));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u4003 (
    .a(\u2_Display/clk1s ),
    .o(\u2_Display/n36 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u4004 (
    .a(\u2_Display/i [9]),
    .o(\u2_Display/n140 [0]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u4005 (
    .a(\u2_Display/j [9]),
    .o(\u2_Display/n99 [0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u401 (
    .a(\u2_Display/n419 [6]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [6]),
    .o(\u2_Display/n445 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u402 (
    .a(\u2_Display/n419 [7]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [7]),
    .o(\u2_Display/n444 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u403 (
    .a(\u2_Display/n419 [8]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [8]),
    .o(\u2_Display/n443 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u404 (
    .a(\u2_Display/n419 [9]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [9]),
    .o(\u2_Display/n442 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u405 (
    .a(\u2_Display/n419 [10]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [10]),
    .o(\u2_Display/n441 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u406 (
    .a(\u2_Display/n419 [11]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [11]),
    .o(\u2_Display/n440 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u407 (
    .a(\u2_Display/n419 [12]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [12]),
    .o(\u2_Display/n439 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u408 (
    .a(\u2_Display/n419 [13]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [13]),
    .o(\u2_Display/n438 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u409 (
    .a(\u2_Display/n419 [14]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [14]),
    .o(\u2_Display/n437 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u410 (
    .a(\u2_Display/n419 [15]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [15]),
    .o(\u2_Display/n436 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u411 (
    .a(\u2_Display/n419 [16]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [16]),
    .o(\u2_Display/n435 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u412 (
    .a(\u2_Display/n419 [17]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [17]),
    .o(\u2_Display/n434 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u413 (
    .a(\u2_Display/n419 [18]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [18]),
    .o(\u2_Display/n433 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u414 (
    .a(\u2_Display/n419 [19]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [19]),
    .o(\u2_Display/n432 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u415 (
    .a(\u2_Display/n419 [20]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [20]),
    .o(\u2_Display/n431 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u416 (
    .a(\u2_Display/n419 [21]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [21]),
    .o(\u2_Display/n430 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u417 (
    .a(\u2_Display/n419 [22]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [22]),
    .o(\u2_Display/n429 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u418 (
    .a(\u2_Display/n419 [23]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [23]),
    .o(\u2_Display/n428 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u419 (
    .a(\u2_Display/n419 [24]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [24]),
    .o(\u2_Display/n427 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u420 (
    .a(\u2_Display/n419 [25]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [25]),
    .o(\u2_Display/n426 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u421 (
    .a(\u2_Display/n419 [26]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [26]),
    .o(\u2_Display/n425 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u422 (
    .a(\u2_Display/n419 [27]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [27]),
    .o(\u2_Display/n424 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u423 (
    .a(\u2_Display/n419 [28]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [28]),
    .o(\u2_Display/n423 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u424 (
    .a(\u2_Display/n419 [29]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [29]),
    .o(\u2_Display/n422 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u425 (
    .a(\u2_Display/n419 [30]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [30]),
    .o(\u2_Display/n421 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u426 (
    .a(\u2_Display/n419 [31]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [31]),
    .o(\u2_Display/n420 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u427 (
    .a(\u2_Display/n1542 [0]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [0]),
    .o(\u2_Display/n1574 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u428 (
    .a(\u2_Display/n1542 [1]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [1]),
    .o(\u2_Display/n1573 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u429 (
    .a(\u2_Display/n1542 [2]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [2]),
    .o(\u2_Display/n1572 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u430 (
    .a(\u2_Display/n1542 [3]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [3]),
    .o(\u2_Display/n1571 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u431 (
    .a(\u2_Display/n1542 [4]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [4]),
    .o(\u2_Display/n1570 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u432 (
    .a(\u2_Display/n1542 [5]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [5]),
    .o(\u2_Display/n1569 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u433 (
    .a(\u2_Display/n1542 [6]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [6]),
    .o(\u2_Display/n1568 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u434 (
    .a(\u2_Display/n1542 [7]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [7]),
    .o(\u2_Display/n1567 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u435 (
    .a(\u2_Display/n1542 [8]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [8]),
    .o(\u2_Display/n1566 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u436 (
    .a(\u2_Display/n1542 [9]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [9]),
    .o(\u2_Display/n1565 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u437 (
    .a(\u2_Display/n1542 [10]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [10]),
    .o(\u2_Display/n1564 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u438 (
    .a(\u2_Display/n1542 [11]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [11]),
    .o(\u2_Display/n1563 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u439 (
    .a(\u2_Display/n1542 [12]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [12]),
    .o(\u2_Display/n1562 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u440 (
    .a(\u2_Display/n1542 [13]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [13]),
    .o(\u2_Display/n1561 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u441 (
    .a(\u2_Display/n1542 [14]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [14]),
    .o(\u2_Display/n1560 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u442 (
    .a(\u2_Display/n1542 [15]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [15]),
    .o(\u2_Display/n1559 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u443 (
    .a(\u2_Display/n1542 [16]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [16]),
    .o(\u2_Display/n1558 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u444 (
    .a(\u2_Display/n1542 [17]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [17]),
    .o(\u2_Display/n1557 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u445 (
    .a(\u2_Display/n1542 [18]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [18]),
    .o(\u2_Display/n1556 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u446 (
    .a(\u2_Display/n1542 [19]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [19]),
    .o(\u2_Display/n1555 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u447 (
    .a(\u2_Display/n1542 [20]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [20]),
    .o(\u2_Display/n1554 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u448 (
    .a(\u2_Display/n1542 [21]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [21]),
    .o(\u2_Display/n1553 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u449 (
    .a(\u2_Display/n1542 [22]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [22]),
    .o(\u2_Display/n1552 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u450 (
    .a(\u2_Display/n1542 [23]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [23]),
    .o(\u2_Display/n1551 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u451 (
    .a(\u2_Display/n1542 [24]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [24]),
    .o(\u2_Display/n1550 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u452 (
    .a(\u2_Display/n1542 [25]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [25]),
    .o(\u2_Display/n1549 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u453 (
    .a(\u2_Display/n1542 [26]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [26]),
    .o(\u2_Display/n1548 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u454 (
    .a(\u2_Display/n1542 [27]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [27]),
    .o(\u2_Display/n1547 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u455 (
    .a(\u2_Display/n1542 [28]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [28]),
    .o(\u2_Display/n1546 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u456 (
    .a(\u2_Display/n1542 [29]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [29]),
    .o(\u2_Display/n1545 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u457 (
    .a(\u2_Display/n1542 [30]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [30]),
    .o(\u2_Display/n1544 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u458 (
    .a(\u2_Display/n1542 [31]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [31]),
    .o(\u2_Display/n1543 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u459 (
    .a(\u2_Display/n2665 [0]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [0]),
    .o(\u2_Display/n2697 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u460 (
    .a(\u2_Display/n2665 [1]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [1]),
    .o(\u2_Display/n2696 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u461 (
    .a(\u2_Display/n2665 [2]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [2]),
    .o(\u2_Display/n2695 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u462 (
    .a(\u2_Display/n2665 [3]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [3]),
    .o(\u2_Display/n2694 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u463 (
    .a(\u2_Display/n2665 [4]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [4]),
    .o(\u2_Display/n2693 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u464 (
    .a(\u2_Display/n2665 [5]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [5]),
    .o(\u2_Display/n2692 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u465 (
    .a(\u2_Display/n2665 [6]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [6]),
    .o(\u2_Display/n2691 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u466 (
    .a(\u2_Display/n2665 [7]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [7]),
    .o(\u2_Display/n2690 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u467 (
    .a(\u2_Display/n2665 [8]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [8]),
    .o(\u2_Display/n2689 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u468 (
    .a(\u2_Display/n2665 [9]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [9]),
    .o(\u2_Display/n2688 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u469 (
    .a(\u2_Display/n2665 [10]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [10]),
    .o(\u2_Display/n2687 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u470 (
    .a(\u2_Display/n2665 [11]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [11]),
    .o(\u2_Display/n2686 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u471 (
    .a(\u2_Display/n2665 [12]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [12]),
    .o(\u2_Display/n2685 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u472 (
    .a(\u2_Display/n2665 [13]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [13]),
    .o(\u2_Display/n2684 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u473 (
    .a(\u2_Display/n2665 [14]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [14]),
    .o(\u2_Display/n2683 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u474 (
    .a(\u2_Display/n2665 [15]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [15]),
    .o(\u2_Display/n2682 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u475 (
    .a(\u2_Display/n2665 [16]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [16]),
    .o(\u2_Display/n2681 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u476 (
    .a(\u2_Display/n2665 [17]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [17]),
    .o(\u2_Display/n2680 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u477 (
    .a(\u2_Display/n2665 [18]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [18]),
    .o(\u2_Display/n2679 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u478 (
    .a(\u2_Display/n2665 [19]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [19]),
    .o(\u2_Display/n2678 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u479 (
    .a(\u2_Display/n2665 [20]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [20]),
    .o(\u2_Display/n2677 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u480 (
    .a(\u2_Display/n2665 [21]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [21]),
    .o(\u2_Display/n2676 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u481 (
    .a(\u2_Display/n2665 [22]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [22]),
    .o(\u2_Display/n2675 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u482 (
    .a(\u2_Display/n2665 [23]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [23]),
    .o(\u2_Display/n2674 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u483 (
    .a(\u2_Display/n2665 [24]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [24]),
    .o(\u2_Display/n2673 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u484 (
    .a(\u2_Display/n2665 [25]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [25]),
    .o(\u2_Display/n2672 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u485 (
    .a(\u2_Display/n2665 [26]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [26]),
    .o(\u2_Display/n2671 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u486 (
    .a(\u2_Display/n2665 [27]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [27]),
    .o(\u2_Display/n2670 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u487 (
    .a(\u2_Display/n2665 [28]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [28]),
    .o(\u2_Display/n2669 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u488 (
    .a(\u2_Display/n2665 [29]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [29]),
    .o(\u2_Display/n2668 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u489 (
    .a(\u2_Display/n2665 [30]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [30]),
    .o(\u2_Display/n2667 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u490 (
    .a(\u2_Display/n2665 [31]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [31]),
    .o(\u2_Display/n2666 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u491 (
    .a(vga_de_pad),
    .b(lcd_data[23]),
    .o(vga_b_pad[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u492 (
    .a(\u1_Driver/n14 ),
    .b(\u1_Driver/n15 ),
    .c(\u1_Driver/n17 ),
    .d(\u1_Driver/n18 ),
    .o(\u1_Driver/lcd_request ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u493 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [9]),
    .o(lcd_ypos[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u494 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [8]),
    .o(lcd_ypos[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u495 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [7]),
    .o(lcd_ypos[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u496 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [6]),
    .o(lcd_ypos[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u497 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [5]),
    .o(lcd_ypos[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u498 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [4]),
    .o(lcd_ypos[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u499 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [3]),
    .o(lcd_ypos[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u500 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [2]),
    .o(lcd_ypos[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u501 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [11]),
    .o(lcd_ypos[11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u502 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [10]),
    .o(lcd_ypos[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u503 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [1]),
    .o(lcd_ypos[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u504 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [0]),
    .o(lcd_ypos[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u505 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [9]),
    .o(lcd_xpos[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u506 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [8]),
    .o(lcd_xpos[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u507 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [7]),
    .o(lcd_xpos[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u508 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [6]),
    .o(lcd_xpos[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u509 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [5]),
    .o(lcd_xpos[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u510 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [4]),
    .o(lcd_xpos[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u511 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [3]),
    .o(lcd_xpos[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u512 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [2]),
    .o(lcd_xpos[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u513 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [11]),
    .o(lcd_xpos[11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u514 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [10]),
    .o(lcd_xpos[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u515 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [1]),
    .o(lcd_xpos[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u516 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [0]),
    .o(lcd_xpos[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u517 (
    .a(\u2_Display/n3820 ),
    .b(\u2_Display/n3823 [0]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3855 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u518 (
    .a(\u2_Display/n3819 ),
    .b(\u2_Display/n3823 [1]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3854 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u519 (
    .a(\u2_Display/n3818 ),
    .b(\u2_Display/n3823 [2]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3853 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u520 (
    .a(\u2_Display/n3817 ),
    .b(\u2_Display/n3823 [3]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3852 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u521 (
    .a(\u2_Display/n3816 ),
    .b(\u2_Display/n3823 [4]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3851 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u522 (
    .a(\u2_Display/n3815 ),
    .b(\u2_Display/n3823 [5]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3850 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u523 (
    .a(\u2_Display/n3814 ),
    .b(\u2_Display/n3823 [6]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3849 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u524 (
    .a(\u2_Display/n3813 ),
    .b(\u2_Display/n3823 [7]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3848 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u525 (
    .a(\u2_Display/n3812 ),
    .b(\u2_Display/n3823 [8]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3847 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u526 (
    .a(\u2_Display/n3811 ),
    .b(\u2_Display/n3823 [9]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3846 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u527 (
    .a(\u2_Display/n3810 ),
    .b(\u2_Display/n3823 [10]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3845 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u528 (
    .a(\u2_Display/n3809 ),
    .b(\u2_Display/n3823 [11]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3844 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u529 (
    .a(\u2_Display/n3808 ),
    .b(\u2_Display/n3823 [12]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3843 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u530 (
    .a(\u2_Display/n3807 ),
    .b(\u2_Display/n3823 [13]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3842 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u531 (
    .a(\u2_Display/n3806 ),
    .b(\u2_Display/n3823 [14]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3841 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u532 (
    .a(\u2_Display/n3805 ),
    .b(\u2_Display/n3823 [15]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3840 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u533 (
    .a(\u2_Display/n3804 ),
    .b(\u2_Display/n3823 [16]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3839 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u534 (
    .a(\u2_Display/n3803 ),
    .b(\u2_Display/n3823 [17]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3838 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u535 (
    .a(\u2_Display/n3802 ),
    .b(\u2_Display/n3823 [18]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3837 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u536 (
    .a(\u2_Display/n3801 ),
    .b(\u2_Display/n3823 [19]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3836 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u537 (
    .a(\u2_Display/n3800 ),
    .b(\u2_Display/n3823 [20]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3835 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u538 (
    .a(\u2_Display/n3799 ),
    .b(\u2_Display/n3823 [21]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3834 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u539 (
    .a(\u2_Display/n3798 ),
    .b(\u2_Display/n3823 [22]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3833 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u540 (
    .a(\u2_Display/n3797 ),
    .b(\u2_Display/n3823 [23]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3832 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u541 (
    .a(\u2_Display/n3796 ),
    .b(\u2_Display/n3823 [24]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3831 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u542 (
    .a(\u2_Display/n3795 ),
    .b(\u2_Display/n3823 [25]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3830 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u543 (
    .a(\u2_Display/n3794 ),
    .b(\u2_Display/n3823 [26]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3829 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u544 (
    .a(\u2_Display/n3793 ),
    .b(\u2_Display/n3823 [27]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3828 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u545 (
    .a(\u2_Display/n3792 ),
    .b(\u2_Display/n3823 [28]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3827 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u546 (
    .a(\u2_Display/n3791 ),
    .b(\u2_Display/n3823 [29]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3826 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u547 (
    .a(\u2_Display/n3790 ),
    .b(\u2_Display/n3823 [30]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3825 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u548 (
    .a(\u2_Display/n3789 ),
    .b(\u2_Display/n3823 [31]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3824 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u549 (
    .a(\u2_Display/n6101 ),
    .b(\u2_Display/n4946 [0]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6136 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u550 (
    .a(\u2_Display/n6100 ),
    .b(\u2_Display/n4946 [1]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6135 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u551 (
    .a(\u2_Display/n6099 ),
    .b(\u2_Display/n4946 [2]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6134 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u552 (
    .a(\u2_Display/n6098 ),
    .b(\u2_Display/n4946 [3]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6133 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u553 (
    .a(\u2_Display/n6097 ),
    .b(\u2_Display/n4946 [4]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6132 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u554 (
    .a(\u2_Display/n6096 ),
    .b(\u2_Display/n4946 [5]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6131 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u555 (
    .a(\u2_Display/n6095 ),
    .b(\u2_Display/n4946 [6]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6130 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u556 (
    .a(\u2_Display/n6094 ),
    .b(\u2_Display/n4946 [7]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6129 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u557 (
    .a(\u2_Display/n6093 ),
    .b(\u2_Display/n4946 [8]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6128 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u558 (
    .a(\u2_Display/n6092 ),
    .b(\u2_Display/n4946 [9]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6127 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u559 (
    .a(\u2_Display/n6091 ),
    .b(\u2_Display/n4946 [10]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6126 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u560 (
    .a(\u2_Display/n6090 ),
    .b(\u2_Display/n4946 [11]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6125 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u561 (
    .a(\u2_Display/n6089 ),
    .b(\u2_Display/n4946 [12]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6124 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u562 (
    .a(\u2_Display/n6088 ),
    .b(\u2_Display/n4946 [13]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6123 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u563 (
    .a(\u2_Display/n6087 ),
    .b(\u2_Display/n4946 [14]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6122 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u564 (
    .a(\u2_Display/n6086 ),
    .b(\u2_Display/n4946 [15]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6121 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u565 (
    .a(\u2_Display/n6085 ),
    .b(\u2_Display/n4946 [16]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6120 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u566 (
    .a(\u2_Display/n6084 ),
    .b(\u2_Display/n4946 [17]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6119 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u567 (
    .a(\u2_Display/n6083 ),
    .b(\u2_Display/n4946 [18]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6118 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u568 (
    .a(\u2_Display/n6082 ),
    .b(\u2_Display/n4946 [19]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6117 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u569 (
    .a(\u2_Display/n6081 ),
    .b(\u2_Display/n4946 [20]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6116 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u570 (
    .a(\u2_Display/n6080 ),
    .b(\u2_Display/n4946 [21]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6115 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u571 (
    .a(\u2_Display/n6079 ),
    .b(\u2_Display/n4946 [22]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6114 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u572 (
    .a(\u2_Display/n6078 ),
    .b(\u2_Display/n4946 [23]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6113 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u573 (
    .a(\u2_Display/n6077 ),
    .b(\u2_Display/n4946 [24]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6112 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u574 (
    .a(\u2_Display/n6076 ),
    .b(\u2_Display/n4946 [25]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6111 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u575 (
    .a(\u2_Display/n6075 ),
    .b(\u2_Display/n4946 [26]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6110 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u576 (
    .a(\u2_Display/n6074 ),
    .b(\u2_Display/n4946 [27]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6109 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u577 (
    .a(\u2_Display/n6073 ),
    .b(\u2_Display/n4946 [28]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6108 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u578 (
    .a(\u2_Display/n6072 ),
    .b(\u2_Display/n4946 [29]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6107 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u579 (
    .a(\u2_Display/n6071 ),
    .b(\u2_Display/n4946 [30]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6106 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u580 (
    .a(\u2_Display/n6070 ),
    .b(\u2_Display/n4946 [31]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6105 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u581 (
    .a(\u2_Display/n451 ),
    .b(\u2_Display/n454 [0]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n486 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u582 (
    .a(\u2_Display/n450 ),
    .b(\u2_Display/n454 [1]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n485 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u583 (
    .a(\u2_Display/n449 ),
    .b(\u2_Display/n454 [2]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n484 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u584 (
    .a(\u2_Display/n448 ),
    .b(\u2_Display/n454 [3]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n483 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u585 (
    .a(\u2_Display/n447 ),
    .b(\u2_Display/n454 [4]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n482 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u586 (
    .a(\u2_Display/n446 ),
    .b(\u2_Display/n454 [5]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n481 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u587 (
    .a(\u2_Display/n445 ),
    .b(\u2_Display/n454 [6]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n480 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u588 (
    .a(\u2_Display/n444 ),
    .b(\u2_Display/n454 [7]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n479 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u589 (
    .a(\u2_Display/n443 ),
    .b(\u2_Display/n454 [8]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n478 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u590 (
    .a(\u2_Display/n442 ),
    .b(\u2_Display/n454 [9]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n477 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u591 (
    .a(\u2_Display/n441 ),
    .b(\u2_Display/n454 [10]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n476 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u592 (
    .a(\u2_Display/n440 ),
    .b(\u2_Display/n454 [11]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n475 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u593 (
    .a(\u2_Display/n439 ),
    .b(\u2_Display/n454 [12]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n474 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u594 (
    .a(\u2_Display/n438 ),
    .b(\u2_Display/n454 [13]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n473 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u595 (
    .a(\u2_Display/n437 ),
    .b(\u2_Display/n454 [14]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n472 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u596 (
    .a(\u2_Display/n436 ),
    .b(\u2_Display/n454 [15]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n471 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u597 (
    .a(\u2_Display/n435 ),
    .b(\u2_Display/n454 [16]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n470 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u598 (
    .a(\u2_Display/n434 ),
    .b(\u2_Display/n454 [17]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n469 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u599 (
    .a(\u2_Display/n433 ),
    .b(\u2_Display/n454 [18]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n468 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u600 (
    .a(\u2_Display/n432 ),
    .b(\u2_Display/n454 [19]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n467 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u601 (
    .a(\u2_Display/n431 ),
    .b(\u2_Display/n454 [20]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n466 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u602 (
    .a(\u2_Display/n430 ),
    .b(\u2_Display/n454 [21]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n465 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u603 (
    .a(\u2_Display/n429 ),
    .b(\u2_Display/n454 [22]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n464 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u604 (
    .a(\u2_Display/n428 ),
    .b(\u2_Display/n454 [23]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n463 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u605 (
    .a(\u2_Display/n427 ),
    .b(\u2_Display/n454 [24]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n462 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u606 (
    .a(\u2_Display/n426 ),
    .b(\u2_Display/n454 [25]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n461 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u607 (
    .a(\u2_Display/n425 ),
    .b(\u2_Display/n454 [26]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n460 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u608 (
    .a(\u2_Display/n424 ),
    .b(\u2_Display/n454 [27]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n459 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u609 (
    .a(\u2_Display/n423 ),
    .b(\u2_Display/n454 [28]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n458 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u610 (
    .a(\u2_Display/n422 ),
    .b(\u2_Display/n454 [29]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n457 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u611 (
    .a(\u2_Display/n421 ),
    .b(\u2_Display/n454 [30]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n456 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u612 (
    .a(\u2_Display/n420 ),
    .b(\u2_Display/n454 [31]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n455 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u613 (
    .a(\u2_Display/n1574 ),
    .b(\u2_Display/n1577 [0]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1609 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u614 (
    .a(\u2_Display/n1573 ),
    .b(\u2_Display/n1577 [1]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1608 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u615 (
    .a(\u2_Display/n1572 ),
    .b(\u2_Display/n1577 [2]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1607 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u616 (
    .a(\u2_Display/n1571 ),
    .b(\u2_Display/n1577 [3]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1606 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u617 (
    .a(\u2_Display/n1570 ),
    .b(\u2_Display/n1577 [4]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1605 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u618 (
    .a(\u2_Display/n1569 ),
    .b(\u2_Display/n1577 [5]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1604 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u619 (
    .a(\u2_Display/n1568 ),
    .b(\u2_Display/n1577 [6]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1603 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u620 (
    .a(\u2_Display/n1567 ),
    .b(\u2_Display/n1577 [7]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1602 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u621 (
    .a(\u2_Display/n1566 ),
    .b(\u2_Display/n1577 [8]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1601 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u622 (
    .a(\u2_Display/n1565 ),
    .b(\u2_Display/n1577 [9]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1600 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u623 (
    .a(\u2_Display/n1564 ),
    .b(\u2_Display/n1577 [10]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1599 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u624 (
    .a(\u2_Display/n1563 ),
    .b(\u2_Display/n1577 [11]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1598 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u625 (
    .a(\u2_Display/n1562 ),
    .b(\u2_Display/n1577 [12]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1597 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u626 (
    .a(\u2_Display/n1561 ),
    .b(\u2_Display/n1577 [13]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1596 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u627 (
    .a(\u2_Display/n1560 ),
    .b(\u2_Display/n1577 [14]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1595 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u628 (
    .a(\u2_Display/n1559 ),
    .b(\u2_Display/n1577 [15]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1594 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u629 (
    .a(\u2_Display/n1558 ),
    .b(\u2_Display/n1577 [16]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1593 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u630 (
    .a(\u2_Display/n1557 ),
    .b(\u2_Display/n1577 [17]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1592 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u631 (
    .a(\u2_Display/n1556 ),
    .b(\u2_Display/n1577 [18]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1591 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u632 (
    .a(\u2_Display/n1555 ),
    .b(\u2_Display/n1577 [19]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1590 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u633 (
    .a(\u2_Display/n1554 ),
    .b(\u2_Display/n1577 [20]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1589 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u634 (
    .a(\u2_Display/n1553 ),
    .b(\u2_Display/n1577 [21]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1588 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u635 (
    .a(\u2_Display/n1552 ),
    .b(\u2_Display/n1577 [22]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1587 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u636 (
    .a(\u2_Display/n1551 ),
    .b(\u2_Display/n1577 [23]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1586 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u637 (
    .a(\u2_Display/n1550 ),
    .b(\u2_Display/n1577 [24]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1585 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u638 (
    .a(\u2_Display/n1549 ),
    .b(\u2_Display/n1577 [25]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1584 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u639 (
    .a(\u2_Display/n1548 ),
    .b(\u2_Display/n1577 [26]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1583 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u640 (
    .a(\u2_Display/n1547 ),
    .b(\u2_Display/n1577 [27]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1582 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u641 (
    .a(\u2_Display/n1546 ),
    .b(\u2_Display/n1577 [28]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1581 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u642 (
    .a(\u2_Display/n1545 ),
    .b(\u2_Display/n1577 [29]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1580 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u643 (
    .a(\u2_Display/n1544 ),
    .b(\u2_Display/n1577 [30]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1579 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u644 (
    .a(\u2_Display/n1543 ),
    .b(\u2_Display/n1577 [31]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1578 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u645 (
    .a(\u2_Display/n2697 ),
    .b(\u2_Display/n2700 [0]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2732 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u646 (
    .a(\u2_Display/n2696 ),
    .b(\u2_Display/n2700 [1]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2731 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u647 (
    .a(\u2_Display/n2695 ),
    .b(\u2_Display/n2700 [2]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2730 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u648 (
    .a(\u2_Display/n2694 ),
    .b(\u2_Display/n2700 [3]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2729 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u649 (
    .a(\u2_Display/n2693 ),
    .b(\u2_Display/n2700 [4]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2728 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u650 (
    .a(\u2_Display/n2692 ),
    .b(\u2_Display/n2700 [5]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2727 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u651 (
    .a(\u2_Display/n2691 ),
    .b(\u2_Display/n2700 [6]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2726 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u652 (
    .a(\u2_Display/n2690 ),
    .b(\u2_Display/n2700 [7]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2725 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u653 (
    .a(\u2_Display/n2689 ),
    .b(\u2_Display/n2700 [8]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2724 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u654 (
    .a(\u2_Display/n2688 ),
    .b(\u2_Display/n2700 [9]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2723 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u655 (
    .a(\u2_Display/n2687 ),
    .b(\u2_Display/n2700 [10]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2722 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u656 (
    .a(\u2_Display/n2686 ),
    .b(\u2_Display/n2700 [11]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2721 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u657 (
    .a(\u2_Display/n2685 ),
    .b(\u2_Display/n2700 [12]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2720 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u658 (
    .a(\u2_Display/n2684 ),
    .b(\u2_Display/n2700 [13]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2719 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u659 (
    .a(\u2_Display/n2683 ),
    .b(\u2_Display/n2700 [14]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2718 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u660 (
    .a(\u2_Display/n2682 ),
    .b(\u2_Display/n2700 [15]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2717 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u661 (
    .a(\u2_Display/n2681 ),
    .b(\u2_Display/n2700 [16]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2716 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u662 (
    .a(\u2_Display/n2680 ),
    .b(\u2_Display/n2700 [17]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2715 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u663 (
    .a(\u2_Display/n2679 ),
    .b(\u2_Display/n2700 [18]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2714 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u664 (
    .a(\u2_Display/n2678 ),
    .b(\u2_Display/n2700 [19]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2713 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u665 (
    .a(\u2_Display/n2677 ),
    .b(\u2_Display/n2700 [20]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2712 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u666 (
    .a(\u2_Display/n2676 ),
    .b(\u2_Display/n2700 [21]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2711 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u667 (
    .a(\u2_Display/n2675 ),
    .b(\u2_Display/n2700 [22]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2710 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u668 (
    .a(\u2_Display/n2674 ),
    .b(\u2_Display/n2700 [23]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2709 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u669 (
    .a(\u2_Display/n2673 ),
    .b(\u2_Display/n2700 [24]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2708 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u670 (
    .a(\u2_Display/n2672 ),
    .b(\u2_Display/n2700 [25]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2707 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u671 (
    .a(\u2_Display/n2671 ),
    .b(\u2_Display/n2700 [26]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2706 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u672 (
    .a(\u2_Display/n2670 ),
    .b(\u2_Display/n2700 [27]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2705 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u673 (
    .a(\u2_Display/n2669 ),
    .b(\u2_Display/n2700 [28]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2704 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u674 (
    .a(\u2_Display/n2668 ),
    .b(\u2_Display/n2700 [29]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2703 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u675 (
    .a(\u2_Display/n2667 ),
    .b(\u2_Display/n2700 [30]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2702 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u676 (
    .a(\u2_Display/n2666 ),
    .b(\u2_Display/n2700 [31]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2701 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u677 (
    .a(\u2_Display/n3855 ),
    .b(\u2_Display/n3858 [0]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3890 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u678 (
    .a(\u2_Display/n3854 ),
    .b(\u2_Display/n3858 [1]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3889 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u679 (
    .a(\u2_Display/n3853 ),
    .b(\u2_Display/n3858 [2]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3888 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u680 (
    .a(\u2_Display/n3852 ),
    .b(\u2_Display/n3858 [3]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3887 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u681 (
    .a(\u2_Display/n3851 ),
    .b(\u2_Display/n3858 [4]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3886 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u682 (
    .a(\u2_Display/n3850 ),
    .b(\u2_Display/n3858 [5]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3885 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u683 (
    .a(\u2_Display/n3849 ),
    .b(\u2_Display/n3858 [6]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3884 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u684 (
    .a(\u2_Display/n3848 ),
    .b(\u2_Display/n3858 [7]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3883 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u685 (
    .a(\u2_Display/n3847 ),
    .b(\u2_Display/n3858 [8]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3882 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u686 (
    .a(\u2_Display/n3846 ),
    .b(\u2_Display/n3858 [9]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3881 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u687 (
    .a(\u2_Display/n3845 ),
    .b(\u2_Display/n3858 [10]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3880 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u688 (
    .a(\u2_Display/n3844 ),
    .b(\u2_Display/n3858 [11]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3879 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u689 (
    .a(\u2_Display/n3843 ),
    .b(\u2_Display/n3858 [12]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3878 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u690 (
    .a(\u2_Display/n3842 ),
    .b(\u2_Display/n3858 [13]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3877 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u691 (
    .a(\u2_Display/n3841 ),
    .b(\u2_Display/n3858 [14]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3876 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u692 (
    .a(\u2_Display/n3840 ),
    .b(\u2_Display/n3858 [15]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3875 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u693 (
    .a(\u2_Display/n3839 ),
    .b(\u2_Display/n3858 [16]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3874 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u694 (
    .a(\u2_Display/n3838 ),
    .b(\u2_Display/n3858 [17]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3873 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u695 (
    .a(\u2_Display/n3837 ),
    .b(\u2_Display/n3858 [18]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3872 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u696 (
    .a(\u2_Display/n3836 ),
    .b(\u2_Display/n3858 [19]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3871 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u697 (
    .a(\u2_Display/n3835 ),
    .b(\u2_Display/n3858 [20]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3870 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u698 (
    .a(\u2_Display/n3834 ),
    .b(\u2_Display/n3858 [21]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3869 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u699 (
    .a(\u2_Display/n3833 ),
    .b(\u2_Display/n3858 [22]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3868 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u700 (
    .a(\u2_Display/n3832 ),
    .b(\u2_Display/n3858 [23]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3867 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u701 (
    .a(\u2_Display/n3831 ),
    .b(\u2_Display/n3858 [24]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3866 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u702 (
    .a(\u2_Display/n3830 ),
    .b(\u2_Display/n3858 [25]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3865 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u703 (
    .a(\u2_Display/n3829 ),
    .b(\u2_Display/n3858 [26]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3864 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u704 (
    .a(\u2_Display/n3828 ),
    .b(\u2_Display/n3858 [27]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3863 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u705 (
    .a(\u2_Display/n3827 ),
    .b(\u2_Display/n3858 [28]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3862 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u706 (
    .a(\u2_Display/n3826 ),
    .b(\u2_Display/n3858 [29]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3861 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u707 (
    .a(\u2_Display/n3825 ),
    .b(\u2_Display/n3858 [30]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3860 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u708 (
    .a(\u2_Display/n3824 ),
    .b(\u2_Display/n3858 [31]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3859 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u709 (
    .a(\u2_Display/n6136 ),
    .b(\u2_Display/n4981 [0]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6171 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u710 (
    .a(\u2_Display/n6135 ),
    .b(\u2_Display/n4981 [1]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6170 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u711 (
    .a(\u2_Display/n6134 ),
    .b(\u2_Display/n4981 [2]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6169 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u712 (
    .a(\u2_Display/n6133 ),
    .b(\u2_Display/n4981 [3]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6168 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u713 (
    .a(\u2_Display/n6132 ),
    .b(\u2_Display/n4981 [4]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6167 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u714 (
    .a(\u2_Display/n6131 ),
    .b(\u2_Display/n4981 [5]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6166 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u715 (
    .a(\u2_Display/n6130 ),
    .b(\u2_Display/n4981 [6]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6165 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u716 (
    .a(\u2_Display/n6129 ),
    .b(\u2_Display/n4981 [7]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6164 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u717 (
    .a(\u2_Display/n6128 ),
    .b(\u2_Display/n4981 [8]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6163 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u718 (
    .a(\u2_Display/n6127 ),
    .b(\u2_Display/n4981 [9]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6162 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u719 (
    .a(\u2_Display/n6126 ),
    .b(\u2_Display/n4981 [10]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6161 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u720 (
    .a(\u2_Display/n6125 ),
    .b(\u2_Display/n4981 [11]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6160 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u721 (
    .a(\u2_Display/n6124 ),
    .b(\u2_Display/n4981 [12]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6159 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u722 (
    .a(\u2_Display/n6123 ),
    .b(\u2_Display/n4981 [13]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6158 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u723 (
    .a(\u2_Display/n6122 ),
    .b(\u2_Display/n4981 [14]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6157 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u724 (
    .a(\u2_Display/n6121 ),
    .b(\u2_Display/n4981 [15]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6156 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u725 (
    .a(\u2_Display/n6120 ),
    .b(\u2_Display/n4981 [16]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6155 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u726 (
    .a(\u2_Display/n6119 ),
    .b(\u2_Display/n4981 [17]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6154 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u727 (
    .a(\u2_Display/n6118 ),
    .b(\u2_Display/n4981 [18]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6153 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u728 (
    .a(\u2_Display/n6117 ),
    .b(\u2_Display/n4981 [19]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6152 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u729 (
    .a(\u2_Display/n6116 ),
    .b(\u2_Display/n4981 [20]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6151 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u730 (
    .a(\u2_Display/n6115 ),
    .b(\u2_Display/n4981 [21]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6150 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u731 (
    .a(\u2_Display/n6114 ),
    .b(\u2_Display/n4981 [22]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6149 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u732 (
    .a(\u2_Display/n6113 ),
    .b(\u2_Display/n4981 [23]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6148 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u733 (
    .a(\u2_Display/n6112 ),
    .b(\u2_Display/n4981 [24]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6147 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u734 (
    .a(\u2_Display/n6111 ),
    .b(\u2_Display/n4981 [25]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6146 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u735 (
    .a(\u2_Display/n6110 ),
    .b(\u2_Display/n4981 [26]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6145 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u736 (
    .a(\u2_Display/n6109 ),
    .b(\u2_Display/n4981 [27]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6144 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u737 (
    .a(\u2_Display/n6108 ),
    .b(\u2_Display/n4981 [28]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6143 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u738 (
    .a(\u2_Display/n6107 ),
    .b(\u2_Display/n4981 [29]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6142 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u739 (
    .a(\u2_Display/n6106 ),
    .b(\u2_Display/n4981 [30]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6141 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u740 (
    .a(\u2_Display/n6105 ),
    .b(\u2_Display/n4981 [31]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6140 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u741 (
    .a(\u2_Display/n486 ),
    .b(\u2_Display/n489 [0]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n521 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u742 (
    .a(\u2_Display/n485 ),
    .b(\u2_Display/n489 [1]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n520 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u743 (
    .a(\u2_Display/n484 ),
    .b(\u2_Display/n489 [2]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n519 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u744 (
    .a(\u2_Display/n483 ),
    .b(\u2_Display/n489 [3]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n518 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u745 (
    .a(\u2_Display/n482 ),
    .b(\u2_Display/n489 [4]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n517 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u746 (
    .a(\u2_Display/n481 ),
    .b(\u2_Display/n489 [5]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n516 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u747 (
    .a(\u2_Display/n480 ),
    .b(\u2_Display/n489 [6]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n515 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u748 (
    .a(\u2_Display/n479 ),
    .b(\u2_Display/n489 [7]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n514 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u749 (
    .a(\u2_Display/n478 ),
    .b(\u2_Display/n489 [8]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n513 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u750 (
    .a(\u2_Display/n477 ),
    .b(\u2_Display/n489 [9]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n512 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u751 (
    .a(\u2_Display/n476 ),
    .b(\u2_Display/n489 [10]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n511 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u752 (
    .a(\u2_Display/n475 ),
    .b(\u2_Display/n489 [11]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n510 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u753 (
    .a(\u2_Display/n474 ),
    .b(\u2_Display/n489 [12]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n509 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u754 (
    .a(\u2_Display/n473 ),
    .b(\u2_Display/n489 [13]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n508 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u755 (
    .a(\u2_Display/n472 ),
    .b(\u2_Display/n489 [14]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n507 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u756 (
    .a(\u2_Display/n471 ),
    .b(\u2_Display/n489 [15]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n506 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u757 (
    .a(\u2_Display/n470 ),
    .b(\u2_Display/n489 [16]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n505 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u758 (
    .a(\u2_Display/n469 ),
    .b(\u2_Display/n489 [17]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n504 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u759 (
    .a(\u2_Display/n468 ),
    .b(\u2_Display/n489 [18]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n503 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u760 (
    .a(\u2_Display/n467 ),
    .b(\u2_Display/n489 [19]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n502 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u761 (
    .a(\u2_Display/n466 ),
    .b(\u2_Display/n489 [20]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n501 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u762 (
    .a(\u2_Display/n465 ),
    .b(\u2_Display/n489 [21]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n500 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u763 (
    .a(\u2_Display/n464 ),
    .b(\u2_Display/n489 [22]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n499 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u764 (
    .a(\u2_Display/n463 ),
    .b(\u2_Display/n489 [23]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n498 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u765 (
    .a(\u2_Display/n462 ),
    .b(\u2_Display/n489 [24]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n497 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u766 (
    .a(\u2_Display/n461 ),
    .b(\u2_Display/n489 [25]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n496 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u767 (
    .a(\u2_Display/n460 ),
    .b(\u2_Display/n489 [26]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n495 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u768 (
    .a(\u2_Display/n459 ),
    .b(\u2_Display/n489 [27]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n494 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u769 (
    .a(\u2_Display/n458 ),
    .b(\u2_Display/n489 [28]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n493 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u770 (
    .a(\u2_Display/n457 ),
    .b(\u2_Display/n489 [29]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n492 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u771 (
    .a(\u2_Display/n456 ),
    .b(\u2_Display/n489 [30]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n491 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u772 (
    .a(\u2_Display/n455 ),
    .b(\u2_Display/n489 [31]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n490 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u773 (
    .a(\u2_Display/n1609 ),
    .b(\u2_Display/n1612 [0]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1644 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u774 (
    .a(\u2_Display/n1608 ),
    .b(\u2_Display/n1612 [1]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1643 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u775 (
    .a(\u2_Display/n1607 ),
    .b(\u2_Display/n1612 [2]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1642 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u776 (
    .a(\u2_Display/n1606 ),
    .b(\u2_Display/n1612 [3]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1641 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u777 (
    .a(\u2_Display/n1605 ),
    .b(\u2_Display/n1612 [4]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1640 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u778 (
    .a(\u2_Display/n1604 ),
    .b(\u2_Display/n1612 [5]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1639 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u779 (
    .a(\u2_Display/n1603 ),
    .b(\u2_Display/n1612 [6]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1638 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u780 (
    .a(\u2_Display/n1602 ),
    .b(\u2_Display/n1612 [7]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1637 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u781 (
    .a(\u2_Display/n1601 ),
    .b(\u2_Display/n1612 [8]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1636 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u782 (
    .a(\u2_Display/n1600 ),
    .b(\u2_Display/n1612 [9]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1635 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u783 (
    .a(\u2_Display/n1599 ),
    .b(\u2_Display/n1612 [10]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1634 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u784 (
    .a(\u2_Display/n1598 ),
    .b(\u2_Display/n1612 [11]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1633 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u785 (
    .a(\u2_Display/n1597 ),
    .b(\u2_Display/n1612 [12]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1632 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u786 (
    .a(\u2_Display/n1596 ),
    .b(\u2_Display/n1612 [13]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1631 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u787 (
    .a(\u2_Display/n1595 ),
    .b(\u2_Display/n1612 [14]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1630 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u788 (
    .a(\u2_Display/n1594 ),
    .b(\u2_Display/n1612 [15]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1629 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u789 (
    .a(\u2_Display/n1593 ),
    .b(\u2_Display/n1612 [16]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1628 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u790 (
    .a(\u2_Display/n1592 ),
    .b(\u2_Display/n1612 [17]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1627 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u791 (
    .a(\u2_Display/n1591 ),
    .b(\u2_Display/n1612 [18]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1626 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u792 (
    .a(\u2_Display/n1590 ),
    .b(\u2_Display/n1612 [19]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1625 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u793 (
    .a(\u2_Display/n1589 ),
    .b(\u2_Display/n1612 [20]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1624 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u794 (
    .a(\u2_Display/n1588 ),
    .b(\u2_Display/n1612 [21]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1623 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u795 (
    .a(\u2_Display/n1587 ),
    .b(\u2_Display/n1612 [22]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1622 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u796 (
    .a(\u2_Display/n1586 ),
    .b(\u2_Display/n1612 [23]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1621 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u797 (
    .a(\u2_Display/n1585 ),
    .b(\u2_Display/n1612 [24]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1620 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u798 (
    .a(\u2_Display/n1584 ),
    .b(\u2_Display/n1612 [25]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1619 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u799 (
    .a(\u2_Display/n1583 ),
    .b(\u2_Display/n1612 [26]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1618 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u800 (
    .a(\u2_Display/n1582 ),
    .b(\u2_Display/n1612 [27]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1617 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u801 (
    .a(\u2_Display/n1581 ),
    .b(\u2_Display/n1612 [28]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1616 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u802 (
    .a(\u2_Display/n1580 ),
    .b(\u2_Display/n1612 [29]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1615 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u803 (
    .a(\u2_Display/n1579 ),
    .b(\u2_Display/n1612 [30]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1614 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u804 (
    .a(\u2_Display/n1578 ),
    .b(\u2_Display/n1612 [31]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1613 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u805 (
    .a(\u2_Display/n2732 ),
    .b(\u2_Display/n2735 [0]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2767 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u806 (
    .a(\u2_Display/n2731 ),
    .b(\u2_Display/n2735 [1]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2766 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u807 (
    .a(\u2_Display/n2730 ),
    .b(\u2_Display/n2735 [2]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2765 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u808 (
    .a(\u2_Display/n2729 ),
    .b(\u2_Display/n2735 [3]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2764 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u809 (
    .a(\u2_Display/n2728 ),
    .b(\u2_Display/n2735 [4]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2763 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u810 (
    .a(\u2_Display/n2727 ),
    .b(\u2_Display/n2735 [5]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2762 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u811 (
    .a(\u2_Display/n2726 ),
    .b(\u2_Display/n2735 [6]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2761 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u812 (
    .a(\u2_Display/n2725 ),
    .b(\u2_Display/n2735 [7]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2760 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u813 (
    .a(\u2_Display/n2724 ),
    .b(\u2_Display/n2735 [8]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2759 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u814 (
    .a(\u2_Display/n2723 ),
    .b(\u2_Display/n2735 [9]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2758 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u815 (
    .a(\u2_Display/n2722 ),
    .b(\u2_Display/n2735 [10]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2757 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u816 (
    .a(\u2_Display/n2721 ),
    .b(\u2_Display/n2735 [11]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2756 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u817 (
    .a(\u2_Display/n2720 ),
    .b(\u2_Display/n2735 [12]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2755 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u818 (
    .a(\u2_Display/n2719 ),
    .b(\u2_Display/n2735 [13]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2754 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u819 (
    .a(\u2_Display/n2718 ),
    .b(\u2_Display/n2735 [14]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2753 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u820 (
    .a(\u2_Display/n2717 ),
    .b(\u2_Display/n2735 [15]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2752 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u821 (
    .a(\u2_Display/n2716 ),
    .b(\u2_Display/n2735 [16]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2751 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u822 (
    .a(\u2_Display/n2715 ),
    .b(\u2_Display/n2735 [17]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2750 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u823 (
    .a(\u2_Display/n2714 ),
    .b(\u2_Display/n2735 [18]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2749 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u824 (
    .a(\u2_Display/n2713 ),
    .b(\u2_Display/n2735 [19]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2748 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u825 (
    .a(\u2_Display/n2712 ),
    .b(\u2_Display/n2735 [20]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2747 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u826 (
    .a(\u2_Display/n2711 ),
    .b(\u2_Display/n2735 [21]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2746 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u827 (
    .a(\u2_Display/n2710 ),
    .b(\u2_Display/n2735 [22]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2745 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u828 (
    .a(\u2_Display/n2709 ),
    .b(\u2_Display/n2735 [23]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2744 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u829 (
    .a(\u2_Display/n2708 ),
    .b(\u2_Display/n2735 [24]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2743 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u830 (
    .a(\u2_Display/n2707 ),
    .b(\u2_Display/n2735 [25]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2742 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u831 (
    .a(\u2_Display/n2706 ),
    .b(\u2_Display/n2735 [26]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2741 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u832 (
    .a(\u2_Display/n2705 ),
    .b(\u2_Display/n2735 [27]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2740 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u833 (
    .a(\u2_Display/n2704 ),
    .b(\u2_Display/n2735 [28]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2739 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u834 (
    .a(\u2_Display/n2703 ),
    .b(\u2_Display/n2735 [29]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2738 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u835 (
    .a(\u2_Display/n2702 ),
    .b(\u2_Display/n2735 [30]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2737 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u836 (
    .a(\u2_Display/n2701 ),
    .b(\u2_Display/n2735 [31]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2736 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u837 (
    .a(\u2_Display/n3890 ),
    .b(\u2_Display/n3893 [0]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3925 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u838 (
    .a(\u2_Display/n3889 ),
    .b(\u2_Display/n3893 [1]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3924 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u839 (
    .a(\u2_Display/n3888 ),
    .b(\u2_Display/n3893 [2]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3923 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u840 (
    .a(\u2_Display/n3887 ),
    .b(\u2_Display/n3893 [3]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3922 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u841 (
    .a(\u2_Display/n3886 ),
    .b(\u2_Display/n3893 [4]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3921 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u842 (
    .a(\u2_Display/n3885 ),
    .b(\u2_Display/n3893 [5]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3920 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u843 (
    .a(\u2_Display/n3884 ),
    .b(\u2_Display/n3893 [6]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3919 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u844 (
    .a(\u2_Display/n3883 ),
    .b(\u2_Display/n3893 [7]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3918 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u845 (
    .a(\u2_Display/n3882 ),
    .b(\u2_Display/n3893 [8]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3917 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u846 (
    .a(\u2_Display/n3881 ),
    .b(\u2_Display/n3893 [9]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3916 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u847 (
    .a(\u2_Display/n3880 ),
    .b(\u2_Display/n3893 [10]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3915 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u848 (
    .a(\u2_Display/n3879 ),
    .b(\u2_Display/n3893 [11]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3914 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u849 (
    .a(\u2_Display/n3878 ),
    .b(\u2_Display/n3893 [12]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3913 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u850 (
    .a(\u2_Display/n3877 ),
    .b(\u2_Display/n3893 [13]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3912 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u851 (
    .a(\u2_Display/n3876 ),
    .b(\u2_Display/n3893 [14]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3911 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u852 (
    .a(\u2_Display/n3875 ),
    .b(\u2_Display/n3893 [15]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3910 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u853 (
    .a(\u2_Display/n3874 ),
    .b(\u2_Display/n3893 [16]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3909 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u854 (
    .a(\u2_Display/n3873 ),
    .b(\u2_Display/n3893 [17]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3908 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u855 (
    .a(\u2_Display/n3872 ),
    .b(\u2_Display/n3893 [18]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3907 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u856 (
    .a(\u2_Display/n3871 ),
    .b(\u2_Display/n3893 [19]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3906 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u857 (
    .a(\u2_Display/n3870 ),
    .b(\u2_Display/n3893 [20]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3905 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u858 (
    .a(\u2_Display/n3869 ),
    .b(\u2_Display/n3893 [21]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3904 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u859 (
    .a(\u2_Display/n3868 ),
    .b(\u2_Display/n3893 [22]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3903 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u860 (
    .a(\u2_Display/n3867 ),
    .b(\u2_Display/n3893 [23]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3902 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u861 (
    .a(\u2_Display/n3866 ),
    .b(\u2_Display/n3893 [24]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3901 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u862 (
    .a(\u2_Display/n3865 ),
    .b(\u2_Display/n3893 [25]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3900 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u863 (
    .a(\u2_Display/n3864 ),
    .b(\u2_Display/n3893 [26]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3899 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u864 (
    .a(\u2_Display/n3863 ),
    .b(\u2_Display/n3893 [27]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3898 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u865 (
    .a(\u2_Display/n3862 ),
    .b(\u2_Display/n3893 [28]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3897 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u866 (
    .a(\u2_Display/n3861 ),
    .b(\u2_Display/n3893 [29]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3896 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u867 (
    .a(\u2_Display/n3860 ),
    .b(\u2_Display/n3893 [30]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3895 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u868 (
    .a(\u2_Display/n3859 ),
    .b(\u2_Display/n3893 [31]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3894 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u869 (
    .a(\u2_Display/n6171 ),
    .b(\u2_Display/n5016 [0]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6206 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u870 (
    .a(\u2_Display/n6170 ),
    .b(\u2_Display/n5016 [1]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6205 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u871 (
    .a(\u2_Display/n6169 ),
    .b(\u2_Display/n5016 [2]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6204 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u872 (
    .a(\u2_Display/n6168 ),
    .b(\u2_Display/n5016 [3]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6203 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u873 (
    .a(\u2_Display/n6167 ),
    .b(\u2_Display/n5016 [4]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6202 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u874 (
    .a(\u2_Display/n6166 ),
    .b(\u2_Display/n5016 [5]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6201 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u875 (
    .a(\u2_Display/n6165 ),
    .b(\u2_Display/n5016 [6]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6200 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u876 (
    .a(\u2_Display/n6164 ),
    .b(\u2_Display/n5016 [7]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6199 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u877 (
    .a(\u2_Display/n6163 ),
    .b(\u2_Display/n5016 [8]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6198 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u878 (
    .a(\u2_Display/n6162 ),
    .b(\u2_Display/n5016 [9]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6197 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u879 (
    .a(\u2_Display/n6161 ),
    .b(\u2_Display/n5016 [10]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6196 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u880 (
    .a(\u2_Display/n6160 ),
    .b(\u2_Display/n5016 [11]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6195 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u881 (
    .a(\u2_Display/n6159 ),
    .b(\u2_Display/n5016 [12]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6194 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u882 (
    .a(\u2_Display/n6158 ),
    .b(\u2_Display/n5016 [13]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6193 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u883 (
    .a(\u2_Display/n6157 ),
    .b(\u2_Display/n5016 [14]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6192 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u884 (
    .a(\u2_Display/n6156 ),
    .b(\u2_Display/n5016 [15]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6191 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u885 (
    .a(\u2_Display/n6155 ),
    .b(\u2_Display/n5016 [16]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6190 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u886 (
    .a(\u2_Display/n6154 ),
    .b(\u2_Display/n5016 [17]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6189 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u887 (
    .a(\u2_Display/n6153 ),
    .b(\u2_Display/n5016 [18]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6188 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u888 (
    .a(\u2_Display/n6152 ),
    .b(\u2_Display/n5016 [19]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6187 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u889 (
    .a(\u2_Display/n6151 ),
    .b(\u2_Display/n5016 [20]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6186 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u890 (
    .a(\u2_Display/n6150 ),
    .b(\u2_Display/n5016 [21]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6185 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u891 (
    .a(\u2_Display/n6149 ),
    .b(\u2_Display/n5016 [22]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6184 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u892 (
    .a(\u2_Display/n6148 ),
    .b(\u2_Display/n5016 [23]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6183 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u893 (
    .a(\u2_Display/n6147 ),
    .b(\u2_Display/n5016 [24]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6182 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u894 (
    .a(\u2_Display/n6146 ),
    .b(\u2_Display/n5016 [25]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6181 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u895 (
    .a(\u2_Display/n6145 ),
    .b(\u2_Display/n5016 [26]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6180 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u896 (
    .a(\u2_Display/n6144 ),
    .b(\u2_Display/n5016 [27]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6179 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u897 (
    .a(\u2_Display/n6143 ),
    .b(\u2_Display/n5016 [28]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6178 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u898 (
    .a(\u2_Display/n6142 ),
    .b(\u2_Display/n5016 [29]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6177 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u899 (
    .a(\u2_Display/n6141 ),
    .b(\u2_Display/n5016 [30]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6176 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u900 (
    .a(\u2_Display/n6140 ),
    .b(\u2_Display/n5016 [31]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6175 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u901 (
    .a(\u2_Display/n521 ),
    .b(\u2_Display/n524 [0]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n556 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u902 (
    .a(\u2_Display/n520 ),
    .b(\u2_Display/n524 [1]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n555 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u903 (
    .a(\u2_Display/n519 ),
    .b(\u2_Display/n524 [2]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n554 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u904 (
    .a(\u2_Display/n518 ),
    .b(\u2_Display/n524 [3]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n553 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u905 (
    .a(\u2_Display/n517 ),
    .b(\u2_Display/n524 [4]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n552 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u906 (
    .a(\u2_Display/n516 ),
    .b(\u2_Display/n524 [5]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n551 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u907 (
    .a(\u2_Display/n515 ),
    .b(\u2_Display/n524 [6]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n550 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u908 (
    .a(\u2_Display/n514 ),
    .b(\u2_Display/n524 [7]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n549 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u909 (
    .a(\u2_Display/n513 ),
    .b(\u2_Display/n524 [8]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n548 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u910 (
    .a(\u2_Display/n512 ),
    .b(\u2_Display/n524 [9]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n547 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u911 (
    .a(\u2_Display/n511 ),
    .b(\u2_Display/n524 [10]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n546 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u912 (
    .a(\u2_Display/n510 ),
    .b(\u2_Display/n524 [11]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n545 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u913 (
    .a(\u2_Display/n509 ),
    .b(\u2_Display/n524 [12]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n544 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u914 (
    .a(\u2_Display/n508 ),
    .b(\u2_Display/n524 [13]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n543 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u915 (
    .a(\u2_Display/n507 ),
    .b(\u2_Display/n524 [14]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n542 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u916 (
    .a(\u2_Display/n506 ),
    .b(\u2_Display/n524 [15]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n541 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u917 (
    .a(\u2_Display/n505 ),
    .b(\u2_Display/n524 [16]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n540 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u918 (
    .a(\u2_Display/n504 ),
    .b(\u2_Display/n524 [17]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n539 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u919 (
    .a(\u2_Display/n503 ),
    .b(\u2_Display/n524 [18]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n538 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u920 (
    .a(\u2_Display/n502 ),
    .b(\u2_Display/n524 [19]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n537 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u921 (
    .a(\u2_Display/n501 ),
    .b(\u2_Display/n524 [20]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n536 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u922 (
    .a(\u2_Display/n500 ),
    .b(\u2_Display/n524 [21]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n535 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u923 (
    .a(\u2_Display/n499 ),
    .b(\u2_Display/n524 [22]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n534 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u924 (
    .a(\u2_Display/n498 ),
    .b(\u2_Display/n524 [23]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n533 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u925 (
    .a(\u2_Display/n497 ),
    .b(\u2_Display/n524 [24]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n532 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u926 (
    .a(\u2_Display/n496 ),
    .b(\u2_Display/n524 [25]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n531 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u927 (
    .a(\u2_Display/n495 ),
    .b(\u2_Display/n524 [26]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n530 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u928 (
    .a(\u2_Display/n494 ),
    .b(\u2_Display/n524 [27]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n529 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u929 (
    .a(\u2_Display/n493 ),
    .b(\u2_Display/n524 [28]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n528 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u930 (
    .a(\u2_Display/n492 ),
    .b(\u2_Display/n524 [29]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n527 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u931 (
    .a(\u2_Display/n491 ),
    .b(\u2_Display/n524 [30]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n526 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u932 (
    .a(\u2_Display/n490 ),
    .b(\u2_Display/n524 [31]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n525 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u933 (
    .a(\u2_Display/n1644 ),
    .b(\u2_Display/n1647 [0]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1679 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u934 (
    .a(\u2_Display/n1643 ),
    .b(\u2_Display/n1647 [1]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1678 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u935 (
    .a(\u2_Display/n1642 ),
    .b(\u2_Display/n1647 [2]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1677 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u936 (
    .a(\u2_Display/n1641 ),
    .b(\u2_Display/n1647 [3]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1676 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u937 (
    .a(\u2_Display/n1640 ),
    .b(\u2_Display/n1647 [4]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1675 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u938 (
    .a(\u2_Display/n1639 ),
    .b(\u2_Display/n1647 [5]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1674 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u939 (
    .a(\u2_Display/n1638 ),
    .b(\u2_Display/n1647 [6]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1673 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u940 (
    .a(\u2_Display/n1637 ),
    .b(\u2_Display/n1647 [7]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1672 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u941 (
    .a(\u2_Display/n1636 ),
    .b(\u2_Display/n1647 [8]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1671 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u942 (
    .a(\u2_Display/n1635 ),
    .b(\u2_Display/n1647 [9]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1670 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u943 (
    .a(\u2_Display/n1634 ),
    .b(\u2_Display/n1647 [10]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1669 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u944 (
    .a(\u2_Display/n1633 ),
    .b(\u2_Display/n1647 [11]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1668 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u945 (
    .a(\u2_Display/n1632 ),
    .b(\u2_Display/n1647 [12]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1667 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u946 (
    .a(\u2_Display/n1631 ),
    .b(\u2_Display/n1647 [13]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1666 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u947 (
    .a(\u2_Display/n1630 ),
    .b(\u2_Display/n1647 [14]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1665 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u948 (
    .a(\u2_Display/n1629 ),
    .b(\u2_Display/n1647 [15]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1664 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u949 (
    .a(\u2_Display/n1628 ),
    .b(\u2_Display/n1647 [16]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1663 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u950 (
    .a(\u2_Display/n1627 ),
    .b(\u2_Display/n1647 [17]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1662 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u951 (
    .a(\u2_Display/n1626 ),
    .b(\u2_Display/n1647 [18]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1661 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u952 (
    .a(\u2_Display/n1625 ),
    .b(\u2_Display/n1647 [19]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1660 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u953 (
    .a(\u2_Display/n1624 ),
    .b(\u2_Display/n1647 [20]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1659 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u954 (
    .a(\u2_Display/n1623 ),
    .b(\u2_Display/n1647 [21]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1658 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u955 (
    .a(\u2_Display/n1622 ),
    .b(\u2_Display/n1647 [22]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1657 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u956 (
    .a(\u2_Display/n1621 ),
    .b(\u2_Display/n1647 [23]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1656 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u957 (
    .a(\u2_Display/n1620 ),
    .b(\u2_Display/n1647 [24]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1655 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u958 (
    .a(\u2_Display/n1619 ),
    .b(\u2_Display/n1647 [25]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1654 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u959 (
    .a(\u2_Display/n1618 ),
    .b(\u2_Display/n1647 [26]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1653 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u960 (
    .a(\u2_Display/n1617 ),
    .b(\u2_Display/n1647 [27]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1652 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u961 (
    .a(\u2_Display/n1616 ),
    .b(\u2_Display/n1647 [28]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1651 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u962 (
    .a(\u2_Display/n1615 ),
    .b(\u2_Display/n1647 [29]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1650 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u963 (
    .a(\u2_Display/n1614 ),
    .b(\u2_Display/n1647 [30]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1649 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u964 (
    .a(\u2_Display/n1613 ),
    .b(\u2_Display/n1647 [31]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1648 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u965 (
    .a(\u2_Display/n2767 ),
    .b(\u2_Display/n2770 [0]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2802 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u966 (
    .a(\u2_Display/n2766 ),
    .b(\u2_Display/n2770 [1]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2801 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u967 (
    .a(\u2_Display/n2765 ),
    .b(\u2_Display/n2770 [2]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2800 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u968 (
    .a(\u2_Display/n2764 ),
    .b(\u2_Display/n2770 [3]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2799 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u969 (
    .a(\u2_Display/n2763 ),
    .b(\u2_Display/n2770 [4]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2798 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u970 (
    .a(\u2_Display/n2762 ),
    .b(\u2_Display/n2770 [5]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2797 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u971 (
    .a(\u2_Display/n2761 ),
    .b(\u2_Display/n2770 [6]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2796 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u972 (
    .a(\u2_Display/n2760 ),
    .b(\u2_Display/n2770 [7]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2795 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u973 (
    .a(\u2_Display/n2759 ),
    .b(\u2_Display/n2770 [8]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2794 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u974 (
    .a(\u2_Display/n2758 ),
    .b(\u2_Display/n2770 [9]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2793 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u975 (
    .a(\u2_Display/n2757 ),
    .b(\u2_Display/n2770 [10]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2792 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u976 (
    .a(\u2_Display/n2756 ),
    .b(\u2_Display/n2770 [11]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2791 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u977 (
    .a(\u2_Display/n2755 ),
    .b(\u2_Display/n2770 [12]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2790 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u978 (
    .a(\u2_Display/n2754 ),
    .b(\u2_Display/n2770 [13]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2789 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u979 (
    .a(\u2_Display/n2753 ),
    .b(\u2_Display/n2770 [14]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2788 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u980 (
    .a(\u2_Display/n2752 ),
    .b(\u2_Display/n2770 [15]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2787 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u981 (
    .a(\u2_Display/n2751 ),
    .b(\u2_Display/n2770 [16]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2786 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u982 (
    .a(\u2_Display/n2750 ),
    .b(\u2_Display/n2770 [17]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2785 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u983 (
    .a(\u2_Display/n2749 ),
    .b(\u2_Display/n2770 [18]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2784 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u984 (
    .a(\u2_Display/n2748 ),
    .b(\u2_Display/n2770 [19]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2783 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u985 (
    .a(\u2_Display/n2747 ),
    .b(\u2_Display/n2770 [20]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2782 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u986 (
    .a(\u2_Display/n2746 ),
    .b(\u2_Display/n2770 [21]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2781 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u987 (
    .a(\u2_Display/n2745 ),
    .b(\u2_Display/n2770 [22]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2780 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u988 (
    .a(\u2_Display/n2744 ),
    .b(\u2_Display/n2770 [23]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2779 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u989 (
    .a(\u2_Display/n2743 ),
    .b(\u2_Display/n2770 [24]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2778 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u990 (
    .a(\u2_Display/n2742 ),
    .b(\u2_Display/n2770 [25]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2777 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u991 (
    .a(\u2_Display/n2741 ),
    .b(\u2_Display/n2770 [26]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2776 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u992 (
    .a(\u2_Display/n2740 ),
    .b(\u2_Display/n2770 [27]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2775 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u993 (
    .a(\u2_Display/n2739 ),
    .b(\u2_Display/n2770 [28]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2774 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u994 (
    .a(\u2_Display/n2738 ),
    .b(\u2_Display/n2770 [29]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2773 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u995 (
    .a(\u2_Display/n2737 ),
    .b(\u2_Display/n2770 [30]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2772 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u996 (
    .a(\u2_Display/n2736 ),
    .b(\u2_Display/n2770 [31]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2771 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u997 (
    .a(\u1_Driver/hcnt [0]),
    .b(\u1_Driver/hcnt [1]),
    .c(\u1_Driver/hcnt [10]),
    .d(\u1_Driver/hcnt [11]),
    .o(_al_u997_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    _al_u998 (
    .a(_al_u997_o),
    .b(\u1_Driver/hcnt [2]),
    .c(\u1_Driver/hcnt [3]),
    .d(\u1_Driver/hcnt [4]),
    .e(\u1_Driver/hcnt [5]),
    .o(_al_u998_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*A)"),
    .INIT(32'h00200000))
    _al_u999 (
    .a(_al_u998_o),
    .b(\u1_Driver/hcnt [6]),
    .c(\u1_Driver/hcnt [7]),
    .d(\u1_Driver/hcnt [8]),
    .e(\u1_Driver/hcnt [9]),
    .o(\u1_Driver/n5 ));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  EG_PHY_GCLK \u0_PLL/uut/bufg_feedback  (
    .clki(\u0_PLL/uut/clk0_buf ),
    .clko(clk_vga));  // al_ip/PLL.v(34)
  EG_PHY_PLL #(
    .CLKC0_CPHASE(8),
    .CLKC0_DIV(9),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(1),
    .CLKC1_DIV(1),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_ENABLE("DISABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(1),
    .CLKC2_DIV(1),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("DISABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(1),
    .CLKC3_DIV(1),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("DISABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(9),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("24.000"),
    .FREQ_LOCK_ACCURACY(2),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .REFCLK_DIV(2),
    .REFCLK_SEL("INTERNAL"),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \u0_PLL/uut/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dwe(1'b0),
    .fbclk(clk_vga),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(clk_24m_pad),
    .reset(\u0_PLL/n0 ),
    .stdby(1'b0),
    .clkc({open_n697,open_n698,open_n699,open_n700,\u0_PLL/uut/clk0_buf }));  // al_ip/PLL.v(57)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add0/u0  (
    .a(\u1_Driver/hcnt [0]),
    .b(1'b1),
    .c(\u1_Driver/add0/c0 ),
    .o({\u1_Driver/add0/c1 ,\u1_Driver/n2 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add0/u1  (
    .a(\u1_Driver/hcnt [1]),
    .b(1'b0),
    .c(\u1_Driver/add0/c1 ),
    .o({\u1_Driver/add0/c2 ,\u1_Driver/n2 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add0/u10  (
    .a(\u1_Driver/hcnt [10]),
    .b(1'b0),
    .c(\u1_Driver/add0/c10 ),
    .o({\u1_Driver/add0/c11 ,\u1_Driver/n2 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add0/u11  (
    .a(\u1_Driver/hcnt [11]),
    .b(1'b0),
    .c(\u1_Driver/add0/c11 ),
    .o({open_n711,\u1_Driver/n2 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add0/u2  (
    .a(\u1_Driver/hcnt [2]),
    .b(1'b0),
    .c(\u1_Driver/add0/c2 ),
    .o({\u1_Driver/add0/c3 ,\u1_Driver/n2 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add0/u3  (
    .a(\u1_Driver/hcnt [3]),
    .b(1'b0),
    .c(\u1_Driver/add0/c3 ),
    .o({\u1_Driver/add0/c4 ,\u1_Driver/n2 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add0/u4  (
    .a(\u1_Driver/hcnt [4]),
    .b(1'b0),
    .c(\u1_Driver/add0/c4 ),
    .o({\u1_Driver/add0/c5 ,\u1_Driver/n2 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add0/u5  (
    .a(\u1_Driver/hcnt [5]),
    .b(1'b0),
    .c(\u1_Driver/add0/c5 ),
    .o({\u1_Driver/add0/c6 ,\u1_Driver/n2 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add0/u6  (
    .a(\u1_Driver/hcnt [6]),
    .b(1'b0),
    .c(\u1_Driver/add0/c6 ),
    .o({\u1_Driver/add0/c7 ,\u1_Driver/n2 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add0/u7  (
    .a(\u1_Driver/hcnt [7]),
    .b(1'b0),
    .c(\u1_Driver/add0/c7 ),
    .o({\u1_Driver/add0/c8 ,\u1_Driver/n2 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add0/u8  (
    .a(\u1_Driver/hcnt [8]),
    .b(1'b0),
    .c(\u1_Driver/add0/c8 ),
    .o({\u1_Driver/add0/c9 ,\u1_Driver/n2 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add0/u9  (
    .a(\u1_Driver/hcnt [9]),
    .b(1'b0),
    .c(\u1_Driver/add0/c9 ),
    .o({\u1_Driver/add0/c10 ,\u1_Driver/n2 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u1_Driver/add0/ucin  (
    .a(1'b0),
    .o({\u1_Driver/add0/c0 ,open_n714}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add1/u0  (
    .a(\u1_Driver/vcnt [0]),
    .b(1'b1),
    .c(\u1_Driver/add1/c0 ),
    .o({\u1_Driver/add1/c1 ,\u1_Driver/n7 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add1/u1  (
    .a(\u1_Driver/vcnt [1]),
    .b(1'b0),
    .c(\u1_Driver/add1/c1 ),
    .o({\u1_Driver/add1/c2 ,\u1_Driver/n7 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add1/u10  (
    .a(\u1_Driver/vcnt [10]),
    .b(1'b0),
    .c(\u1_Driver/add1/c10 ),
    .o({\u1_Driver/add1/c11 ,\u1_Driver/n7 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add1/u11  (
    .a(\u1_Driver/vcnt [11]),
    .b(1'b0),
    .c(\u1_Driver/add1/c11 ),
    .o({open_n715,\u1_Driver/n7 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add1/u2  (
    .a(\u1_Driver/vcnt [2]),
    .b(1'b0),
    .c(\u1_Driver/add1/c2 ),
    .o({\u1_Driver/add1/c3 ,\u1_Driver/n7 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add1/u3  (
    .a(\u1_Driver/vcnt [3]),
    .b(1'b0),
    .c(\u1_Driver/add1/c3 ),
    .o({\u1_Driver/add1/c4 ,\u1_Driver/n7 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add1/u4  (
    .a(\u1_Driver/vcnt [4]),
    .b(1'b0),
    .c(\u1_Driver/add1/c4 ),
    .o({\u1_Driver/add1/c5 ,\u1_Driver/n7 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add1/u5  (
    .a(\u1_Driver/vcnt [5]),
    .b(1'b0),
    .c(\u1_Driver/add1/c5 ),
    .o({\u1_Driver/add1/c6 ,\u1_Driver/n7 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add1/u6  (
    .a(\u1_Driver/vcnt [6]),
    .b(1'b0),
    .c(\u1_Driver/add1/c6 ),
    .o({\u1_Driver/add1/c7 ,\u1_Driver/n7 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add1/u7  (
    .a(\u1_Driver/vcnt [7]),
    .b(1'b0),
    .c(\u1_Driver/add1/c7 ),
    .o({\u1_Driver/add1/c8 ,\u1_Driver/n7 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add1/u8  (
    .a(\u1_Driver/vcnt [8]),
    .b(1'b0),
    .c(\u1_Driver/add1/c8 ),
    .o({\u1_Driver/add1/c9 ,\u1_Driver/n7 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u1_Driver/add1/u9  (
    .a(\u1_Driver/vcnt [9]),
    .b(1'b0),
    .c(\u1_Driver/add1/c9 ),
    .o({\u1_Driver/add1/c10 ,\u1_Driver/n7 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u1_Driver/add1/ucin  (
    .a(1'b0),
    .o({\u1_Driver/add1/c0 ,open_n718}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt0_0  (
    .a(\u1_Driver/hcnt [0]),
    .b(1'b1),
    .c(\u1_Driver/lt0_c0 ),
    .o({\u1_Driver/lt0_c1 ,open_n719}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt0_1  (
    .a(\u1_Driver/hcnt [1]),
    .b(1'b1),
    .c(\u1_Driver/lt0_c1 ),
    .o({\u1_Driver/lt0_c2 ,open_n720}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt0_10  (
    .a(\u1_Driver/hcnt [10]),
    .b(1'b1),
    .c(\u1_Driver/lt0_c10 ),
    .o({\u1_Driver/lt0_c11 ,open_n721}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt0_11  (
    .a(\u1_Driver/hcnt [11]),
    .b(1'b0),
    .c(\u1_Driver/lt0_c11 ),
    .o({\u1_Driver/lt0_c12 ,open_n722}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt0_2  (
    .a(\u1_Driver/hcnt [2]),
    .b(1'b1),
    .c(\u1_Driver/lt0_c2 ),
    .o({\u1_Driver/lt0_c3 ,open_n723}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt0_3  (
    .a(\u1_Driver/hcnt [3]),
    .b(1'b0),
    .c(\u1_Driver/lt0_c3 ),
    .o({\u1_Driver/lt0_c4 ,open_n724}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt0_4  (
    .a(\u1_Driver/hcnt [4]),
    .b(1'b1),
    .c(\u1_Driver/lt0_c4 ),
    .o({\u1_Driver/lt0_c5 ,open_n725}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt0_5  (
    .a(\u1_Driver/hcnt [5]),
    .b(1'b0),
    .c(\u1_Driver/lt0_c5 ),
    .o({\u1_Driver/lt0_c6 ,open_n726}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt0_6  (
    .a(\u1_Driver/hcnt [6]),
    .b(1'b0),
    .c(\u1_Driver/lt0_c6 ),
    .o({\u1_Driver/lt0_c7 ,open_n727}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt0_7  (
    .a(\u1_Driver/hcnt [7]),
    .b(1'b1),
    .c(\u1_Driver/lt0_c7 ),
    .o({\u1_Driver/lt0_c8 ,open_n728}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt0_8  (
    .a(\u1_Driver/hcnt [8]),
    .b(1'b0),
    .c(\u1_Driver/lt0_c8 ),
    .o({\u1_Driver/lt0_c9 ,open_n729}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt0_9  (
    .a(\u1_Driver/hcnt [9]),
    .b(1'b1),
    .c(\u1_Driver/lt0_c9 ),
    .o({\u1_Driver/lt0_c10 ,open_n730}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u1_Driver/lt0_cin  (
    .a(1'b0),
    .o({\u1_Driver/lt0_c0 ,open_n733}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt0_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u1_Driver/lt0_c12 ),
    .o({open_n734,\u1_Driver/n1 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt1_0  (
    .a(\u1_Driver/hcnt [0]),
    .b(1'b1),
    .c(\u1_Driver/lt1_c0 ),
    .o({\u1_Driver/lt1_c1 ,open_n735}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt1_1  (
    .a(\u1_Driver/hcnt [1]),
    .b(1'b1),
    .c(\u1_Driver/lt1_c1 ),
    .o({\u1_Driver/lt1_c2 ,open_n736}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt1_10  (
    .a(\u1_Driver/hcnt [10]),
    .b(1'b0),
    .c(\u1_Driver/lt1_c10 ),
    .o({\u1_Driver/lt1_c11 ,open_n737}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt1_11  (
    .a(\u1_Driver/hcnt [11]),
    .b(1'b0),
    .c(\u1_Driver/lt1_c11 ),
    .o({\u1_Driver/lt1_c12 ,open_n738}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt1_2  (
    .a(\u1_Driver/hcnt [2]),
    .b(1'b1),
    .c(\u1_Driver/lt1_c2 ),
    .o({\u1_Driver/lt1_c3 ,open_n739}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt1_3  (
    .a(\u1_Driver/hcnt [3]),
    .b(1'b1),
    .c(\u1_Driver/lt1_c3 ),
    .o({\u1_Driver/lt1_c4 ,open_n740}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt1_4  (
    .a(\u1_Driver/hcnt [4]),
    .b(1'b0),
    .c(\u1_Driver/lt1_c4 ),
    .o({\u1_Driver/lt1_c5 ,open_n741}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt1_5  (
    .a(\u1_Driver/hcnt [5]),
    .b(1'b1),
    .c(\u1_Driver/lt1_c5 ),
    .o({\u1_Driver/lt1_c6 ,open_n742}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt1_6  (
    .a(\u1_Driver/hcnt [6]),
    .b(1'b1),
    .c(\u1_Driver/lt1_c6 ),
    .o({\u1_Driver/lt1_c7 ,open_n743}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt1_7  (
    .a(\u1_Driver/hcnt [7]),
    .b(1'b0),
    .c(\u1_Driver/lt1_c7 ),
    .o({\u1_Driver/lt1_c8 ,open_n744}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt1_8  (
    .a(\u1_Driver/hcnt [8]),
    .b(1'b0),
    .c(\u1_Driver/lt1_c8 ),
    .o({\u1_Driver/lt1_c9 ,open_n745}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt1_9  (
    .a(\u1_Driver/hcnt [9]),
    .b(1'b0),
    .c(\u1_Driver/lt1_c9 ),
    .o({\u1_Driver/lt1_c10 ,open_n746}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u1_Driver/lt1_cin  (
    .a(1'b1),
    .o({\u1_Driver/lt1_c0 ,open_n749}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt1_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u1_Driver/lt1_c12 ),
    .o({open_n750,\u1_Driver/n4 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt2_0  (
    .a(\u1_Driver/vcnt [0]),
    .b(1'b0),
    .c(\u1_Driver/lt2_c0 ),
    .o({\u1_Driver/lt2_c1 ,open_n751}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt2_1  (
    .a(\u1_Driver/vcnt [1]),
    .b(1'b1),
    .c(\u1_Driver/lt2_c1 ),
    .o({\u1_Driver/lt2_c2 ,open_n752}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt2_10  (
    .a(\u1_Driver/vcnt [10]),
    .b(1'b0),
    .c(\u1_Driver/lt2_c10 ),
    .o({\u1_Driver/lt2_c11 ,open_n753}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt2_11  (
    .a(\u1_Driver/vcnt [11]),
    .b(1'b0),
    .c(\u1_Driver/lt2_c11 ),
    .o({\u1_Driver/lt2_c12 ,open_n754}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt2_2  (
    .a(\u1_Driver/vcnt [2]),
    .b(1'b0),
    .c(\u1_Driver/lt2_c2 ),
    .o({\u1_Driver/lt2_c3 ,open_n755}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt2_3  (
    .a(\u1_Driver/vcnt [3]),
    .b(1'b0),
    .c(\u1_Driver/lt2_c3 ),
    .o({\u1_Driver/lt2_c4 ,open_n756}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt2_4  (
    .a(\u1_Driver/vcnt [4]),
    .b(1'b0),
    .c(\u1_Driver/lt2_c4 ),
    .o({\u1_Driver/lt2_c5 ,open_n757}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt2_5  (
    .a(\u1_Driver/vcnt [5]),
    .b(1'b0),
    .c(\u1_Driver/lt2_c5 ),
    .o({\u1_Driver/lt2_c6 ,open_n758}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt2_6  (
    .a(\u1_Driver/vcnt [6]),
    .b(1'b0),
    .c(\u1_Driver/lt2_c6 ),
    .o({\u1_Driver/lt2_c7 ,open_n759}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt2_7  (
    .a(\u1_Driver/vcnt [7]),
    .b(1'b0),
    .c(\u1_Driver/lt2_c7 ),
    .o({\u1_Driver/lt2_c8 ,open_n760}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt2_8  (
    .a(\u1_Driver/vcnt [8]),
    .b(1'b0),
    .c(\u1_Driver/lt2_c8 ),
    .o({\u1_Driver/lt2_c9 ,open_n761}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt2_9  (
    .a(\u1_Driver/vcnt [9]),
    .b(1'b0),
    .c(\u1_Driver/lt2_c9 ),
    .o({\u1_Driver/lt2_c10 ,open_n762}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u1_Driver/lt2_cin  (
    .a(1'b1),
    .o({\u1_Driver/lt2_c0 ,open_n765}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt2_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u1_Driver/lt2_c12 ),
    .o({open_n766,\u1_Driver/n10 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt3_0  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [0]),
    .c(\u1_Driver/lt3_c0 ),
    .o({\u1_Driver/lt3_c1 ,open_n767}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt3_1  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [1]),
    .c(\u1_Driver/lt3_c1 ),
    .o({\u1_Driver/lt3_c2 ,open_n768}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt3_10  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [10]),
    .c(\u1_Driver/lt3_c10 ),
    .o({\u1_Driver/lt3_c11 ,open_n769}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt3_11  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [11]),
    .c(\u1_Driver/lt3_c11 ),
    .o({\u1_Driver/lt3_c12 ,open_n770}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt3_2  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [2]),
    .c(\u1_Driver/lt3_c2 ),
    .o({\u1_Driver/lt3_c3 ,open_n771}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt3_3  (
    .a(1'b1),
    .b(\u1_Driver/hcnt [3]),
    .c(\u1_Driver/lt3_c3 ),
    .o({\u1_Driver/lt3_c4 ,open_n772}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt3_4  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [4]),
    .c(\u1_Driver/lt3_c4 ),
    .o({\u1_Driver/lt3_c5 ,open_n773}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt3_5  (
    .a(1'b1),
    .b(\u1_Driver/hcnt [5]),
    .c(\u1_Driver/lt3_c5 ),
    .o({\u1_Driver/lt3_c6 ,open_n774}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt3_6  (
    .a(1'b1),
    .b(\u1_Driver/hcnt [6]),
    .c(\u1_Driver/lt3_c6 ),
    .o({\u1_Driver/lt3_c7 ,open_n775}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt3_7  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [7]),
    .c(\u1_Driver/lt3_c7 ),
    .o({\u1_Driver/lt3_c8 ,open_n776}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt3_8  (
    .a(1'b1),
    .b(\u1_Driver/hcnt [8]),
    .c(\u1_Driver/lt3_c8 ),
    .o({\u1_Driver/lt3_c9 ,open_n777}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt3_9  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [9]),
    .c(\u1_Driver/lt3_c9 ),
    .o({\u1_Driver/lt3_c10 ,open_n778}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u1_Driver/lt3_cin  (
    .a(1'b1),
    .o({\u1_Driver/lt3_c0 ,open_n781}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt3_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u1_Driver/lt3_c12 ),
    .o({open_n782,\u1_Driver/n11 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt4_0  (
    .a(\u1_Driver/hcnt [0]),
    .b(1'b0),
    .c(\u1_Driver/lt4_c0 ),
    .o({\u1_Driver/lt4_c1 ,open_n783}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt4_1  (
    .a(\u1_Driver/hcnt [1]),
    .b(1'b0),
    .c(\u1_Driver/lt4_c1 ),
    .o({\u1_Driver/lt4_c2 ,open_n784}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt4_10  (
    .a(\u1_Driver/hcnt [10]),
    .b(1'b1),
    .c(\u1_Driver/lt4_c10 ),
    .o({\u1_Driver/lt4_c11 ,open_n785}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt4_11  (
    .a(\u1_Driver/hcnt [11]),
    .b(1'b0),
    .c(\u1_Driver/lt4_c11 ),
    .o({\u1_Driver/lt4_c12 ,open_n786}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt4_2  (
    .a(\u1_Driver/hcnt [2]),
    .b(1'b0),
    .c(\u1_Driver/lt4_c2 ),
    .o({\u1_Driver/lt4_c3 ,open_n787}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt4_3  (
    .a(\u1_Driver/hcnt [3]),
    .b(1'b1),
    .c(\u1_Driver/lt4_c3 ),
    .o({\u1_Driver/lt4_c4 ,open_n788}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt4_4  (
    .a(\u1_Driver/hcnt [4]),
    .b(1'b0),
    .c(\u1_Driver/lt4_c4 ),
    .o({\u1_Driver/lt4_c5 ,open_n789}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt4_5  (
    .a(\u1_Driver/hcnt [5]),
    .b(1'b1),
    .c(\u1_Driver/lt4_c5 ),
    .o({\u1_Driver/lt4_c6 ,open_n790}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt4_6  (
    .a(\u1_Driver/hcnt [6]),
    .b(1'b1),
    .c(\u1_Driver/lt4_c6 ),
    .o({\u1_Driver/lt4_c7 ,open_n791}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt4_7  (
    .a(\u1_Driver/hcnt [7]),
    .b(1'b0),
    .c(\u1_Driver/lt4_c7 ),
    .o({\u1_Driver/lt4_c8 ,open_n792}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt4_8  (
    .a(\u1_Driver/hcnt [8]),
    .b(1'b0),
    .c(\u1_Driver/lt4_c8 ),
    .o({\u1_Driver/lt4_c9 ,open_n793}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt4_9  (
    .a(\u1_Driver/hcnt [9]),
    .b(1'b1),
    .c(\u1_Driver/lt4_c9 ),
    .o({\u1_Driver/lt4_c10 ,open_n794}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u1_Driver/lt4_cin  (
    .a(1'b0),
    .o({\u1_Driver/lt4_c0 ,open_n797}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt4_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u1_Driver/lt4_c12 ),
    .o({open_n798,\u1_Driver/n12 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt5_0  (
    .a(1'b1),
    .b(\u1_Driver/vcnt [0]),
    .c(\u1_Driver/lt5_c0 ),
    .o({\u1_Driver/lt5_c1 ,open_n799}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt5_1  (
    .a(1'b0),
    .b(\u1_Driver/vcnt [1]),
    .c(\u1_Driver/lt5_c1 ),
    .o({\u1_Driver/lt5_c2 ,open_n800}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt5_10  (
    .a(1'b0),
    .b(\u1_Driver/vcnt [10]),
    .c(\u1_Driver/lt5_c10 ),
    .o({\u1_Driver/lt5_c11 ,open_n801}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt5_11  (
    .a(1'b0),
    .b(\u1_Driver/vcnt [11]),
    .c(\u1_Driver/lt5_c11 ),
    .o({\u1_Driver/lt5_c12 ,open_n802}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt5_2  (
    .a(1'b0),
    .b(\u1_Driver/vcnt [2]),
    .c(\u1_Driver/lt5_c2 ),
    .o({\u1_Driver/lt5_c3 ,open_n803}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt5_3  (
    .a(1'b1),
    .b(\u1_Driver/vcnt [3]),
    .c(\u1_Driver/lt5_c3 ),
    .o({\u1_Driver/lt5_c4 ,open_n804}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt5_4  (
    .a(1'b0),
    .b(\u1_Driver/vcnt [4]),
    .c(\u1_Driver/lt5_c4 ),
    .o({\u1_Driver/lt5_c5 ,open_n805}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt5_5  (
    .a(1'b1),
    .b(\u1_Driver/vcnt [5]),
    .c(\u1_Driver/lt5_c5 ),
    .o({\u1_Driver/lt5_c6 ,open_n806}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt5_6  (
    .a(1'b0),
    .b(\u1_Driver/vcnt [6]),
    .c(\u1_Driver/lt5_c6 ),
    .o({\u1_Driver/lt5_c7 ,open_n807}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt5_7  (
    .a(1'b0),
    .b(\u1_Driver/vcnt [7]),
    .c(\u1_Driver/lt5_c7 ),
    .o({\u1_Driver/lt5_c8 ,open_n808}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt5_8  (
    .a(1'b0),
    .b(\u1_Driver/vcnt [8]),
    .c(\u1_Driver/lt5_c8 ),
    .o({\u1_Driver/lt5_c9 ,open_n809}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt5_9  (
    .a(1'b0),
    .b(\u1_Driver/vcnt [9]),
    .c(\u1_Driver/lt5_c9 ),
    .o({\u1_Driver/lt5_c10 ,open_n810}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u1_Driver/lt5_cin  (
    .a(1'b1),
    .o({\u1_Driver/lt5_c0 ,open_n813}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt5_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u1_Driver/lt5_c12 ),
    .o({open_n814,\u1_Driver/n14 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt6_0  (
    .a(\u1_Driver/vcnt [0]),
    .b(1'b1),
    .c(\u1_Driver/lt6_c0 ),
    .o({\u1_Driver/lt6_c1 ,open_n815}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt6_1  (
    .a(\u1_Driver/vcnt [1]),
    .b(1'b0),
    .c(\u1_Driver/lt6_c1 ),
    .o({\u1_Driver/lt6_c2 ,open_n816}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt6_10  (
    .a(\u1_Driver/vcnt [10]),
    .b(1'b1),
    .c(\u1_Driver/lt6_c10 ),
    .o({\u1_Driver/lt6_c11 ,open_n817}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt6_11  (
    .a(\u1_Driver/vcnt [11]),
    .b(1'b0),
    .c(\u1_Driver/lt6_c11 ),
    .o({\u1_Driver/lt6_c12 ,open_n818}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt6_2  (
    .a(\u1_Driver/vcnt [2]),
    .b(1'b0),
    .c(\u1_Driver/lt6_c2 ),
    .o({\u1_Driver/lt6_c3 ,open_n819}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt6_3  (
    .a(\u1_Driver/vcnt [3]),
    .b(1'b1),
    .c(\u1_Driver/lt6_c3 ),
    .o({\u1_Driver/lt6_c4 ,open_n820}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt6_4  (
    .a(\u1_Driver/vcnt [4]),
    .b(1'b0),
    .c(\u1_Driver/lt6_c4 ),
    .o({\u1_Driver/lt6_c5 ,open_n821}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt6_5  (
    .a(\u1_Driver/vcnt [5]),
    .b(1'b1),
    .c(\u1_Driver/lt6_c5 ),
    .o({\u1_Driver/lt6_c6 ,open_n822}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt6_6  (
    .a(\u1_Driver/vcnt [6]),
    .b(1'b0),
    .c(\u1_Driver/lt6_c6 ),
    .o({\u1_Driver/lt6_c7 ,open_n823}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt6_7  (
    .a(\u1_Driver/vcnt [7]),
    .b(1'b0),
    .c(\u1_Driver/lt6_c7 ),
    .o({\u1_Driver/lt6_c8 ,open_n824}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt6_8  (
    .a(\u1_Driver/vcnt [8]),
    .b(1'b0),
    .c(\u1_Driver/lt6_c8 ),
    .o({\u1_Driver/lt6_c9 ,open_n825}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt6_9  (
    .a(\u1_Driver/vcnt [9]),
    .b(1'b0),
    .c(\u1_Driver/lt6_c9 ),
    .o({\u1_Driver/lt6_c10 ,open_n826}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u1_Driver/lt6_cin  (
    .a(1'b0),
    .o({\u1_Driver/lt6_c0 ,open_n829}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt6_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u1_Driver/lt6_c12 ),
    .o({open_n830,\u1_Driver/n15 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt7_0  (
    .a(1'b1),
    .b(\u1_Driver/hcnt [0]),
    .c(\u1_Driver/lt7_c0 ),
    .o({\u1_Driver/lt7_c1 ,open_n831}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt7_1  (
    .a(1'b1),
    .b(\u1_Driver/hcnt [1]),
    .c(\u1_Driver/lt7_c1 ),
    .o({\u1_Driver/lt7_c2 ,open_n832}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt7_10  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [10]),
    .c(\u1_Driver/lt7_c10 ),
    .o({\u1_Driver/lt7_c11 ,open_n833}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt7_11  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [11]),
    .c(\u1_Driver/lt7_c11 ),
    .o({\u1_Driver/lt7_c12 ,open_n834}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt7_2  (
    .a(1'b1),
    .b(\u1_Driver/hcnt [2]),
    .c(\u1_Driver/lt7_c2 ),
    .o({\u1_Driver/lt7_c3 ,open_n835}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt7_3  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [3]),
    .c(\u1_Driver/lt7_c3 ),
    .o({\u1_Driver/lt7_c4 ,open_n836}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt7_4  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [4]),
    .c(\u1_Driver/lt7_c4 ),
    .o({\u1_Driver/lt7_c5 ,open_n837}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt7_5  (
    .a(1'b1),
    .b(\u1_Driver/hcnt [5]),
    .c(\u1_Driver/lt7_c5 ),
    .o({\u1_Driver/lt7_c6 ,open_n838}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt7_6  (
    .a(1'b1),
    .b(\u1_Driver/hcnt [6]),
    .c(\u1_Driver/lt7_c6 ),
    .o({\u1_Driver/lt7_c7 ,open_n839}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt7_7  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [7]),
    .c(\u1_Driver/lt7_c7 ),
    .o({\u1_Driver/lt7_c8 ,open_n840}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt7_8  (
    .a(1'b1),
    .b(\u1_Driver/hcnt [8]),
    .c(\u1_Driver/lt7_c8 ),
    .o({\u1_Driver/lt7_c9 ,open_n841}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt7_9  (
    .a(1'b0),
    .b(\u1_Driver/hcnt [9]),
    .c(\u1_Driver/lt7_c9 ),
    .o({\u1_Driver/lt7_c10 ,open_n842}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u1_Driver/lt7_cin  (
    .a(1'b1),
    .o({\u1_Driver/lt7_c0 ,open_n845}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt7_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u1_Driver/lt7_c12 ),
    .o({open_n846,\u1_Driver/n17 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt8_0  (
    .a(\u1_Driver/hcnt [0]),
    .b(1'b1),
    .c(\u1_Driver/lt8_c0 ),
    .o({\u1_Driver/lt8_c1 ,open_n847}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt8_1  (
    .a(\u1_Driver/hcnt [1]),
    .b(1'b1),
    .c(\u1_Driver/lt8_c1 ),
    .o({\u1_Driver/lt8_c2 ,open_n848}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt8_10  (
    .a(\u1_Driver/hcnt [10]),
    .b(1'b1),
    .c(\u1_Driver/lt8_c10 ),
    .o({\u1_Driver/lt8_c11 ,open_n849}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt8_11  (
    .a(\u1_Driver/hcnt [11]),
    .b(1'b0),
    .c(\u1_Driver/lt8_c11 ),
    .o({\u1_Driver/lt8_c12 ,open_n850}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt8_2  (
    .a(\u1_Driver/hcnt [2]),
    .b(1'b1),
    .c(\u1_Driver/lt8_c2 ),
    .o({\u1_Driver/lt8_c3 ,open_n851}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt8_3  (
    .a(\u1_Driver/hcnt [3]),
    .b(1'b0),
    .c(\u1_Driver/lt8_c3 ),
    .o({\u1_Driver/lt8_c4 ,open_n852}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt8_4  (
    .a(\u1_Driver/hcnt [4]),
    .b(1'b0),
    .c(\u1_Driver/lt8_c4 ),
    .o({\u1_Driver/lt8_c5 ,open_n853}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt8_5  (
    .a(\u1_Driver/hcnt [5]),
    .b(1'b1),
    .c(\u1_Driver/lt8_c5 ),
    .o({\u1_Driver/lt8_c6 ,open_n854}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt8_6  (
    .a(\u1_Driver/hcnt [6]),
    .b(1'b1),
    .c(\u1_Driver/lt8_c6 ),
    .o({\u1_Driver/lt8_c7 ,open_n855}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt8_7  (
    .a(\u1_Driver/hcnt [7]),
    .b(1'b0),
    .c(\u1_Driver/lt8_c7 ),
    .o({\u1_Driver/lt8_c8 ,open_n856}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt8_8  (
    .a(\u1_Driver/hcnt [8]),
    .b(1'b0),
    .c(\u1_Driver/lt8_c8 ),
    .o({\u1_Driver/lt8_c9 ,open_n857}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt8_9  (
    .a(\u1_Driver/hcnt [9]),
    .b(1'b1),
    .c(\u1_Driver/lt8_c9 ),
    .o({\u1_Driver/lt8_c10 ,open_n858}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u1_Driver/lt8_cin  (
    .a(1'b0),
    .o({\u1_Driver/lt8_c0 ,open_n861}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u1_Driver/lt8_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u1_Driver/lt8_c12 ),
    .o({open_n862,\u1_Driver/n18 }));
  reg_ar_as_w1 \u1_Driver/reg0_b0  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [0]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/vcnt [0]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b1  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [1]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/vcnt [1]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b10  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [10]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/vcnt [10]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b11  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [11]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/vcnt [11]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b2  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [2]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/vcnt [2]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b3  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [3]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/vcnt [3]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b4  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [4]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/vcnt [4]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b5  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [5]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/vcnt [5]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b6  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [6]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/vcnt [6]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b7  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [7]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/vcnt [7]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b8  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [8]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/vcnt [8]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg0_b9  (
    .clk(clk_vga),
    .d(\u1_Driver/n8 [9]),
    .en(\u1_Driver/n5 ),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/vcnt [9]));  // source/rtl/Driver.v(78)
  reg_ar_as_w1 \u1_Driver/reg1_b0  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [0]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/hcnt [0]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b1  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [1]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/hcnt [1]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b10  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [10]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/hcnt [10]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b11  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [11]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/hcnt [11]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b2  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [2]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/hcnt [2]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b3  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [3]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/hcnt [3]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b4  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [4]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/hcnt [4]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b5  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [5]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/hcnt [5]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b6  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [6]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/hcnt [6]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b7  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [7]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/hcnt [7]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b8  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [8]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/hcnt [8]));  // source/rtl/Driver.v(62)
  reg_ar_as_w1 \u1_Driver/reg1_b9  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [9]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(\u1_Driver/hcnt [9]));  // source/rtl/Driver.v(62)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub0/u0  (
    .a(\u1_Driver/hcnt [0]),
    .b(1'b1),
    .c(\u1_Driver/sub0/c0 ),
    .o({\u1_Driver/sub0/c1 ,\u1_Driver/n20 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub0/u1  (
    .a(\u1_Driver/hcnt [1]),
    .b(1'b1),
    .c(\u1_Driver/sub0/c1 ),
    .o({\u1_Driver/sub0/c2 ,\u1_Driver/n20 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub0/u10  (
    .a(\u1_Driver/hcnt [10]),
    .b(1'b0),
    .c(\u1_Driver/sub0/c10 ),
    .o({\u1_Driver/sub0/c11 ,\u1_Driver/n20 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub0/u11  (
    .a(\u1_Driver/hcnt [11]),
    .b(1'b0),
    .c(\u1_Driver/sub0/c11 ),
    .o({open_n863,\u1_Driver/n20 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub0/u2  (
    .a(\u1_Driver/hcnt [2]),
    .b(1'b1),
    .c(\u1_Driver/sub0/c2 ),
    .o({\u1_Driver/sub0/c3 ,\u1_Driver/n20 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub0/u3  (
    .a(\u1_Driver/hcnt [3]),
    .b(1'b0),
    .c(\u1_Driver/sub0/c3 ),
    .o({\u1_Driver/sub0/c4 ,\u1_Driver/n20 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub0/u4  (
    .a(\u1_Driver/hcnt [4]),
    .b(1'b0),
    .c(\u1_Driver/sub0/c4 ),
    .o({\u1_Driver/sub0/c5 ,\u1_Driver/n20 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub0/u5  (
    .a(\u1_Driver/hcnt [5]),
    .b(1'b1),
    .c(\u1_Driver/sub0/c5 ),
    .o({\u1_Driver/sub0/c6 ,\u1_Driver/n20 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub0/u6  (
    .a(\u1_Driver/hcnt [6]),
    .b(1'b1),
    .c(\u1_Driver/sub0/c6 ),
    .o({\u1_Driver/sub0/c7 ,\u1_Driver/n20 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub0/u7  (
    .a(\u1_Driver/hcnt [7]),
    .b(1'b0),
    .c(\u1_Driver/sub0/c7 ),
    .o({\u1_Driver/sub0/c8 ,\u1_Driver/n20 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub0/u8  (
    .a(\u1_Driver/hcnt [8]),
    .b(1'b1),
    .c(\u1_Driver/sub0/c8 ),
    .o({\u1_Driver/sub0/c9 ,\u1_Driver/n20 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub0/u9  (
    .a(\u1_Driver/hcnt [9]),
    .b(1'b0),
    .c(\u1_Driver/sub0/c9 ),
    .o({\u1_Driver/sub0/c10 ,\u1_Driver/n20 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u1_Driver/sub0/ucin  (
    .a(1'b0),
    .o({\u1_Driver/sub0/c0 ,open_n866}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub1/u0  (
    .a(\u1_Driver/vcnt [0]),
    .b(1'b1),
    .c(\u1_Driver/sub1/c0 ),
    .o({\u1_Driver/sub1/c1 ,\u1_Driver/n21 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub1/u1  (
    .a(\u1_Driver/vcnt [1]),
    .b(1'b0),
    .c(\u1_Driver/sub1/c1 ),
    .o({\u1_Driver/sub1/c2 ,\u1_Driver/n21 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub1/u10  (
    .a(\u1_Driver/vcnt [10]),
    .b(1'b0),
    .c(\u1_Driver/sub1/c10 ),
    .o({\u1_Driver/sub1/c11 ,\u1_Driver/n21 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub1/u11  (
    .a(\u1_Driver/vcnt [11]),
    .b(1'b0),
    .c(\u1_Driver/sub1/c11 ),
    .o({open_n867,\u1_Driver/n21 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub1/u2  (
    .a(\u1_Driver/vcnt [2]),
    .b(1'b0),
    .c(\u1_Driver/sub1/c2 ),
    .o({\u1_Driver/sub1/c3 ,\u1_Driver/n21 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub1/u3  (
    .a(\u1_Driver/vcnt [3]),
    .b(1'b1),
    .c(\u1_Driver/sub1/c3 ),
    .o({\u1_Driver/sub1/c4 ,\u1_Driver/n21 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub1/u4  (
    .a(\u1_Driver/vcnt [4]),
    .b(1'b0),
    .c(\u1_Driver/sub1/c4 ),
    .o({\u1_Driver/sub1/c5 ,\u1_Driver/n21 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub1/u5  (
    .a(\u1_Driver/vcnt [5]),
    .b(1'b1),
    .c(\u1_Driver/sub1/c5 ),
    .o({\u1_Driver/sub1/c6 ,\u1_Driver/n21 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub1/u6  (
    .a(\u1_Driver/vcnt [6]),
    .b(1'b0),
    .c(\u1_Driver/sub1/c6 ),
    .o({\u1_Driver/sub1/c7 ,\u1_Driver/n21 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub1/u7  (
    .a(\u1_Driver/vcnt [7]),
    .b(1'b0),
    .c(\u1_Driver/sub1/c7 ),
    .o({\u1_Driver/sub1/c8 ,\u1_Driver/n21 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub1/u8  (
    .a(\u1_Driver/vcnt [8]),
    .b(1'b0),
    .c(\u1_Driver/sub1/c8 ),
    .o({\u1_Driver/sub1/c9 ,\u1_Driver/n21 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u1_Driver/sub1/u9  (
    .a(\u1_Driver/vcnt [9]),
    .b(1'b0),
    .c(\u1_Driver/sub1/c9 ),
    .o({\u1_Driver/sub1/c10 ,\u1_Driver/n21 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u1_Driver/sub1/ucin  (
    .a(1'b0),
    .o({\u1_Driver/sub1/c0 ,open_n870}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u0  (
    .a(\u2_Display/n [0]),
    .b(1'b1),
    .c(\u2_Display/add0/c0 ),
    .o({\u2_Display/add0/c1 ,\u2_Display/n37 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u1  (
    .a(\u2_Display/n [1]),
    .b(1'b0),
    .c(\u2_Display/add0/c1 ),
    .o({\u2_Display/add0/c2 ,\u2_Display/n37 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u10  (
    .a(\u2_Display/n [10]),
    .b(1'b0),
    .c(\u2_Display/add0/c10 ),
    .o({\u2_Display/add0/c11 ,\u2_Display/n37 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u11  (
    .a(\u2_Display/n [11]),
    .b(1'b0),
    .c(\u2_Display/add0/c11 ),
    .o({\u2_Display/add0/c12 ,\u2_Display/n37 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u12  (
    .a(\u2_Display/n [12]),
    .b(1'b0),
    .c(\u2_Display/add0/c12 ),
    .o({\u2_Display/add0/c13 ,\u2_Display/n37 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u13  (
    .a(\u2_Display/n [13]),
    .b(1'b0),
    .c(\u2_Display/add0/c13 ),
    .o({\u2_Display/add0/c14 ,\u2_Display/n37 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u14  (
    .a(\u2_Display/n [14]),
    .b(1'b0),
    .c(\u2_Display/add0/c14 ),
    .o({\u2_Display/add0/c15 ,\u2_Display/n37 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u15  (
    .a(\u2_Display/n [15]),
    .b(1'b0),
    .c(\u2_Display/add0/c15 ),
    .o({\u2_Display/add0/c16 ,\u2_Display/n37 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u16  (
    .a(\u2_Display/n [16]),
    .b(1'b0),
    .c(\u2_Display/add0/c16 ),
    .o({\u2_Display/add0/c17 ,\u2_Display/n37 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u17  (
    .a(\u2_Display/n [17]),
    .b(1'b0),
    .c(\u2_Display/add0/c17 ),
    .o({\u2_Display/add0/c18 ,\u2_Display/n37 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u18  (
    .a(\u2_Display/n [18]),
    .b(1'b0),
    .c(\u2_Display/add0/c18 ),
    .o({\u2_Display/add0/c19 ,\u2_Display/n37 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u19  (
    .a(\u2_Display/n [19]),
    .b(1'b0),
    .c(\u2_Display/add0/c19 ),
    .o({\u2_Display/add0/c20 ,\u2_Display/n37 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u2  (
    .a(\u2_Display/n [2]),
    .b(1'b0),
    .c(\u2_Display/add0/c2 ),
    .o({\u2_Display/add0/c3 ,\u2_Display/n37 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u20  (
    .a(\u2_Display/n [20]),
    .b(1'b0),
    .c(\u2_Display/add0/c20 ),
    .o({\u2_Display/add0/c21 ,\u2_Display/n37 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u21  (
    .a(\u2_Display/n [21]),
    .b(1'b0),
    .c(\u2_Display/add0/c21 ),
    .o({\u2_Display/add0/c22 ,\u2_Display/n37 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u22  (
    .a(\u2_Display/n [22]),
    .b(1'b0),
    .c(\u2_Display/add0/c22 ),
    .o({\u2_Display/add0/c23 ,\u2_Display/n37 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u23  (
    .a(\u2_Display/n [23]),
    .b(1'b0),
    .c(\u2_Display/add0/c23 ),
    .o({\u2_Display/add0/c24 ,\u2_Display/n37 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u24  (
    .a(\u2_Display/n [24]),
    .b(1'b0),
    .c(\u2_Display/add0/c24 ),
    .o({\u2_Display/add0/c25 ,\u2_Display/n37 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u25  (
    .a(\u2_Display/n [25]),
    .b(1'b0),
    .c(\u2_Display/add0/c25 ),
    .o({\u2_Display/add0/c26 ,\u2_Display/n37 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u26  (
    .a(\u2_Display/n [26]),
    .b(1'b0),
    .c(\u2_Display/add0/c26 ),
    .o({\u2_Display/add0/c27 ,\u2_Display/n37 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u27  (
    .a(\u2_Display/n [27]),
    .b(1'b0),
    .c(\u2_Display/add0/c27 ),
    .o({\u2_Display/add0/c28 ,\u2_Display/n37 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u28  (
    .a(\u2_Display/n [28]),
    .b(1'b0),
    .c(\u2_Display/add0/c28 ),
    .o({\u2_Display/add0/c29 ,\u2_Display/n37 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u29  (
    .a(\u2_Display/n [29]),
    .b(1'b0),
    .c(\u2_Display/add0/c29 ),
    .o({\u2_Display/add0/c30 ,\u2_Display/n37 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u3  (
    .a(\u2_Display/n [3]),
    .b(1'b0),
    .c(\u2_Display/add0/c3 ),
    .o({\u2_Display/add0/c4 ,\u2_Display/n37 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u30  (
    .a(\u2_Display/n [30]),
    .b(1'b0),
    .c(\u2_Display/add0/c30 ),
    .o({open_n871,\u2_Display/n37 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u4  (
    .a(\u2_Display/n [4]),
    .b(1'b0),
    .c(\u2_Display/add0/c4 ),
    .o({\u2_Display/add0/c5 ,\u2_Display/n37 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u5  (
    .a(\u2_Display/n [5]),
    .b(1'b0),
    .c(\u2_Display/add0/c5 ),
    .o({\u2_Display/add0/c6 ,\u2_Display/n37 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u6  (
    .a(\u2_Display/n [6]),
    .b(1'b0),
    .c(\u2_Display/add0/c6 ),
    .o({\u2_Display/add0/c7 ,\u2_Display/n37 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u7  (
    .a(\u2_Display/n [7]),
    .b(1'b0),
    .c(\u2_Display/add0/c7 ),
    .o({\u2_Display/add0/c8 ,\u2_Display/n37 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u8  (
    .a(\u2_Display/n [8]),
    .b(1'b0),
    .c(\u2_Display/add0/c8 ),
    .o({\u2_Display/add0/c9 ,\u2_Display/n37 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add0/u9  (
    .a(\u2_Display/n [9]),
    .b(1'b0),
    .c(\u2_Display/add0/c9 ),
    .o({\u2_Display/add0/c10 ,\u2_Display/n37 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add0/ucin  (
    .a(1'b0),
    .o({\u2_Display/add0/c0 ,open_n874}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u0  (
    .a(\u2_Display/counta [0]),
    .b(1'b1),
    .c(\u2_Display/add1/c0 ),
    .o({\u2_Display/add1/c1 ,\u2_Display/n41 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u1  (
    .a(\u2_Display/counta [1]),
    .b(1'b0),
    .c(\u2_Display/add1/c1 ),
    .o({\u2_Display/add1/c2 ,\u2_Display/n41 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u10  (
    .a(\u2_Display/counta [10]),
    .b(1'b0),
    .c(\u2_Display/add1/c10 ),
    .o({\u2_Display/add1/c11 ,\u2_Display/n41 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u11  (
    .a(\u2_Display/counta [11]),
    .b(1'b0),
    .c(\u2_Display/add1/c11 ),
    .o({\u2_Display/add1/c12 ,\u2_Display/n41 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u12  (
    .a(\u2_Display/counta [12]),
    .b(1'b0),
    .c(\u2_Display/add1/c12 ),
    .o({\u2_Display/add1/c13 ,\u2_Display/n41 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u13  (
    .a(\u2_Display/counta [13]),
    .b(1'b0),
    .c(\u2_Display/add1/c13 ),
    .o({\u2_Display/add1/c14 ,\u2_Display/n41 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u14  (
    .a(\u2_Display/counta [14]),
    .b(1'b0),
    .c(\u2_Display/add1/c14 ),
    .o({\u2_Display/add1/c15 ,\u2_Display/n41 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u15  (
    .a(\u2_Display/counta [15]),
    .b(1'b0),
    .c(\u2_Display/add1/c15 ),
    .o({\u2_Display/add1/c16 ,\u2_Display/n41 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u16  (
    .a(\u2_Display/counta [16]),
    .b(1'b0),
    .c(\u2_Display/add1/c16 ),
    .o({\u2_Display/add1/c17 ,\u2_Display/n41 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u17  (
    .a(\u2_Display/counta [17]),
    .b(1'b0),
    .c(\u2_Display/add1/c17 ),
    .o({\u2_Display/add1/c18 ,\u2_Display/n41 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u18  (
    .a(\u2_Display/counta [18]),
    .b(1'b0),
    .c(\u2_Display/add1/c18 ),
    .o({\u2_Display/add1/c19 ,\u2_Display/n41 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u19  (
    .a(\u2_Display/counta [19]),
    .b(1'b0),
    .c(\u2_Display/add1/c19 ),
    .o({\u2_Display/add1/c20 ,\u2_Display/n41 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u2  (
    .a(\u2_Display/counta [2]),
    .b(1'b0),
    .c(\u2_Display/add1/c2 ),
    .o({\u2_Display/add1/c3 ,\u2_Display/n41 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u20  (
    .a(\u2_Display/counta [20]),
    .b(1'b0),
    .c(\u2_Display/add1/c20 ),
    .o({\u2_Display/add1/c21 ,\u2_Display/n41 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u21  (
    .a(\u2_Display/counta [21]),
    .b(1'b0),
    .c(\u2_Display/add1/c21 ),
    .o({\u2_Display/add1/c22 ,\u2_Display/n41 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u22  (
    .a(\u2_Display/counta [22]),
    .b(1'b0),
    .c(\u2_Display/add1/c22 ),
    .o({\u2_Display/add1/c23 ,\u2_Display/n41 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u23  (
    .a(\u2_Display/counta [23]),
    .b(1'b0),
    .c(\u2_Display/add1/c23 ),
    .o({\u2_Display/add1/c24 ,\u2_Display/n41 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u24  (
    .a(\u2_Display/counta [24]),
    .b(1'b0),
    .c(\u2_Display/add1/c24 ),
    .o({\u2_Display/add1/c25 ,\u2_Display/n41 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u25  (
    .a(\u2_Display/counta [25]),
    .b(1'b0),
    .c(\u2_Display/add1/c25 ),
    .o({\u2_Display/add1/c26 ,\u2_Display/n41 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u26  (
    .a(\u2_Display/counta [26]),
    .b(1'b0),
    .c(\u2_Display/add1/c26 ),
    .o({\u2_Display/add1/c27 ,\u2_Display/n41 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u27  (
    .a(\u2_Display/counta [27]),
    .b(1'b0),
    .c(\u2_Display/add1/c27 ),
    .o({\u2_Display/add1/c28 ,\u2_Display/n41 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u28  (
    .a(\u2_Display/counta [28]),
    .b(1'b0),
    .c(\u2_Display/add1/c28 ),
    .o({\u2_Display/add1/c29 ,\u2_Display/n41 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u29  (
    .a(\u2_Display/counta [29]),
    .b(1'b0),
    .c(\u2_Display/add1/c29 ),
    .o({\u2_Display/add1/c30 ,\u2_Display/n41 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u3  (
    .a(\u2_Display/counta [3]),
    .b(1'b0),
    .c(\u2_Display/add1/c3 ),
    .o({\u2_Display/add1/c4 ,\u2_Display/n41 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u30  (
    .a(\u2_Display/counta [30]),
    .b(1'b0),
    .c(\u2_Display/add1/c30 ),
    .o({\u2_Display/add1/c31 ,\u2_Display/n41 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u31  (
    .a(\u2_Display/counta [31]),
    .b(1'b0),
    .c(\u2_Display/add1/c31 ),
    .o({open_n875,\u2_Display/n41 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u4  (
    .a(\u2_Display/counta [4]),
    .b(1'b0),
    .c(\u2_Display/add1/c4 ),
    .o({\u2_Display/add1/c5 ,\u2_Display/n41 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u5  (
    .a(\u2_Display/counta [5]),
    .b(1'b0),
    .c(\u2_Display/add1/c5 ),
    .o({\u2_Display/add1/c6 ,\u2_Display/n41 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u6  (
    .a(\u2_Display/counta [6]),
    .b(1'b0),
    .c(\u2_Display/add1/c6 ),
    .o({\u2_Display/add1/c7 ,\u2_Display/n41 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u7  (
    .a(\u2_Display/counta [7]),
    .b(1'b0),
    .c(\u2_Display/add1/c7 ),
    .o({\u2_Display/add1/c8 ,\u2_Display/n41 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u8  (
    .a(\u2_Display/counta [8]),
    .b(1'b0),
    .c(\u2_Display/add1/c8 ),
    .o({\u2_Display/add1/c9 ,\u2_Display/n41 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add1/u9  (
    .a(\u2_Display/counta [9]),
    .b(1'b0),
    .c(\u2_Display/add1/c9 ),
    .o({\u2_Display/add1/c10 ,\u2_Display/n41 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add1/ucin  (
    .a(1'b0),
    .o({\u2_Display/add1/c0 ,open_n878}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u0  (
    .a(\u2_Display/n3222 ),
    .b(1'b1),
    .c(\u2_Display/add100/c0 ),
    .o({\u2_Display/add100/c1 ,\u2_Display/n3225 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u1  (
    .a(\u2_Display/n3221 ),
    .b(1'b1),
    .c(\u2_Display/add100/c1 ),
    .o({\u2_Display/add100/c2 ,\u2_Display/n3225 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u10  (
    .a(\u2_Display/n3212 ),
    .b(1'b0),
    .c(\u2_Display/add100/c10 ),
    .o({\u2_Display/add100/c11 ,\u2_Display/n3225 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u11  (
    .a(\u2_Display/n3211 ),
    .b(1'b1),
    .c(\u2_Display/add100/c11 ),
    .o({\u2_Display/add100/c12 ,\u2_Display/n3225 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u12  (
    .a(\u2_Display/n3210 ),
    .b(1'b0),
    .c(\u2_Display/add100/c12 ),
    .o({\u2_Display/add100/c13 ,\u2_Display/n3225 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u13  (
    .a(\u2_Display/n3209 ),
    .b(1'b1),
    .c(\u2_Display/add100/c13 ),
    .o({\u2_Display/add100/c14 ,\u2_Display/n3225 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u14  (
    .a(\u2_Display/n3208 ),
    .b(1'b1),
    .c(\u2_Display/add100/c14 ),
    .o({\u2_Display/add100/c15 ,\u2_Display/n3225 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u15  (
    .a(\u2_Display/n3207 ),
    .b(1'b0),
    .c(\u2_Display/add100/c15 ),
    .o({\u2_Display/add100/c16 ,\u2_Display/n3225 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u16  (
    .a(\u2_Display/n3206 ),
    .b(1'b1),
    .c(\u2_Display/add100/c16 ),
    .o({\u2_Display/add100/c17 ,\u2_Display/n3225 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u17  (
    .a(\u2_Display/n3205 ),
    .b(1'b1),
    .c(\u2_Display/add100/c17 ),
    .o({\u2_Display/add100/c18 ,\u2_Display/n3225 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u18  (
    .a(\u2_Display/n3204 ),
    .b(1'b1),
    .c(\u2_Display/add100/c18 ),
    .o({\u2_Display/add100/c19 ,\u2_Display/n3225 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u19  (
    .a(\u2_Display/n3203 ),
    .b(1'b1),
    .c(\u2_Display/add100/c19 ),
    .o({\u2_Display/add100/c20 ,\u2_Display/n3225 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u2  (
    .a(\u2_Display/n3220 ),
    .b(1'b1),
    .c(\u2_Display/add100/c2 ),
    .o({\u2_Display/add100/c3 ,\u2_Display/n3225 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u20  (
    .a(\u2_Display/n3202 ),
    .b(1'b1),
    .c(\u2_Display/add100/c20 ),
    .o({\u2_Display/add100/c21 ,\u2_Display/n3225 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u21  (
    .a(\u2_Display/n3201 ),
    .b(1'b1),
    .c(\u2_Display/add100/c21 ),
    .o({\u2_Display/add100/c22 ,\u2_Display/n3225 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u22  (
    .a(\u2_Display/n3200 ),
    .b(1'b1),
    .c(\u2_Display/add100/c22 ),
    .o({\u2_Display/add100/c23 ,\u2_Display/n3225 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u23  (
    .a(\u2_Display/n3199 ),
    .b(1'b1),
    .c(\u2_Display/add100/c23 ),
    .o({\u2_Display/add100/c24 ,\u2_Display/n3225 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u24  (
    .a(\u2_Display/n3198 ),
    .b(1'b1),
    .c(\u2_Display/add100/c24 ),
    .o({\u2_Display/add100/c25 ,\u2_Display/n3225 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u25  (
    .a(\u2_Display/n3197 ),
    .b(1'b1),
    .c(\u2_Display/add100/c25 ),
    .o({\u2_Display/add100/c26 ,\u2_Display/n3225 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u26  (
    .a(\u2_Display/n3196 ),
    .b(1'b1),
    .c(\u2_Display/add100/c26 ),
    .o({\u2_Display/add100/c27 ,\u2_Display/n3225 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u27  (
    .a(\u2_Display/n3195 ),
    .b(1'b1),
    .c(\u2_Display/add100/c27 ),
    .o({\u2_Display/add100/c28 ,\u2_Display/n3225 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u28  (
    .a(\u2_Display/n3194 ),
    .b(1'b1),
    .c(\u2_Display/add100/c28 ),
    .o({\u2_Display/add100/c29 ,\u2_Display/n3225 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u29  (
    .a(\u2_Display/n3193 ),
    .b(1'b1),
    .c(\u2_Display/add100/c29 ),
    .o({\u2_Display/add100/c30 ,\u2_Display/n3225 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u3  (
    .a(\u2_Display/n3219 ),
    .b(1'b1),
    .c(\u2_Display/add100/c3 ),
    .o({\u2_Display/add100/c4 ,\u2_Display/n3225 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u30  (
    .a(\u2_Display/n3192 ),
    .b(1'b1),
    .c(\u2_Display/add100/c30 ),
    .o({\u2_Display/add100/c31 ,\u2_Display/n3225 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u31  (
    .a(\u2_Display/n3191 ),
    .b(1'b1),
    .c(\u2_Display/add100/c31 ),
    .o({open_n879,\u2_Display/n3225 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u4  (
    .a(\u2_Display/n3218 ),
    .b(1'b1),
    .c(\u2_Display/add100/c4 ),
    .o({\u2_Display/add100/c5 ,\u2_Display/n3225 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u5  (
    .a(\u2_Display/n3217 ),
    .b(1'b1),
    .c(\u2_Display/add100/c5 ),
    .o({\u2_Display/add100/c6 ,\u2_Display/n3225 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u6  (
    .a(\u2_Display/n3216 ),
    .b(1'b1),
    .c(\u2_Display/add100/c6 ),
    .o({\u2_Display/add100/c7 ,\u2_Display/n3225 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u7  (
    .a(\u2_Display/n3215 ),
    .b(1'b1),
    .c(\u2_Display/add100/c7 ),
    .o({\u2_Display/add100/c8 ,\u2_Display/n3225 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u8  (
    .a(\u2_Display/n3214 ),
    .b(1'b1),
    .c(\u2_Display/add100/c8 ),
    .o({\u2_Display/add100/c9 ,\u2_Display/n3225 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add100/u9  (
    .a(\u2_Display/n3213 ),
    .b(1'b0),
    .c(\u2_Display/add100/c9 ),
    .o({\u2_Display/add100/c10 ,\u2_Display/n3225 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add100/ucin  (
    .a(1'b1),
    .o({\u2_Display/add100/c0 ,open_n882}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u0  (
    .a(\u2_Display/n3257 ),
    .b(1'b1),
    .c(\u2_Display/add101/c0 ),
    .o({\u2_Display/add101/c1 ,\u2_Display/n3260 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u1  (
    .a(\u2_Display/n3256 ),
    .b(1'b1),
    .c(\u2_Display/add101/c1 ),
    .o({\u2_Display/add101/c2 ,\u2_Display/n3260 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u10  (
    .a(\u2_Display/n3247 ),
    .b(1'b1),
    .c(\u2_Display/add101/c10 ),
    .o({\u2_Display/add101/c11 ,\u2_Display/n3260 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u11  (
    .a(\u2_Display/n3246 ),
    .b(1'b0),
    .c(\u2_Display/add101/c11 ),
    .o({\u2_Display/add101/c12 ,\u2_Display/n3260 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u12  (
    .a(\u2_Display/n3245 ),
    .b(1'b1),
    .c(\u2_Display/add101/c12 ),
    .o({\u2_Display/add101/c13 ,\u2_Display/n3260 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u13  (
    .a(\u2_Display/n3244 ),
    .b(1'b1),
    .c(\u2_Display/add101/c13 ),
    .o({\u2_Display/add101/c14 ,\u2_Display/n3260 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u14  (
    .a(\u2_Display/n3243 ),
    .b(1'b0),
    .c(\u2_Display/add101/c14 ),
    .o({\u2_Display/add101/c15 ,\u2_Display/n3260 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u15  (
    .a(\u2_Display/n3242 ),
    .b(1'b1),
    .c(\u2_Display/add101/c15 ),
    .o({\u2_Display/add101/c16 ,\u2_Display/n3260 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u16  (
    .a(\u2_Display/n3241 ),
    .b(1'b1),
    .c(\u2_Display/add101/c16 ),
    .o({\u2_Display/add101/c17 ,\u2_Display/n3260 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u17  (
    .a(\u2_Display/n3240 ),
    .b(1'b1),
    .c(\u2_Display/add101/c17 ),
    .o({\u2_Display/add101/c18 ,\u2_Display/n3260 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u18  (
    .a(\u2_Display/n3239 ),
    .b(1'b1),
    .c(\u2_Display/add101/c18 ),
    .o({\u2_Display/add101/c19 ,\u2_Display/n3260 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u19  (
    .a(\u2_Display/n3238 ),
    .b(1'b1),
    .c(\u2_Display/add101/c19 ),
    .o({\u2_Display/add101/c20 ,\u2_Display/n3260 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u2  (
    .a(\u2_Display/n3255 ),
    .b(1'b1),
    .c(\u2_Display/add101/c2 ),
    .o({\u2_Display/add101/c3 ,\u2_Display/n3260 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u20  (
    .a(\u2_Display/n3237 ),
    .b(1'b1),
    .c(\u2_Display/add101/c20 ),
    .o({\u2_Display/add101/c21 ,\u2_Display/n3260 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u21  (
    .a(\u2_Display/n3236 ),
    .b(1'b1),
    .c(\u2_Display/add101/c21 ),
    .o({\u2_Display/add101/c22 ,\u2_Display/n3260 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u22  (
    .a(\u2_Display/n3235 ),
    .b(1'b1),
    .c(\u2_Display/add101/c22 ),
    .o({\u2_Display/add101/c23 ,\u2_Display/n3260 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u23  (
    .a(\u2_Display/n3234 ),
    .b(1'b1),
    .c(\u2_Display/add101/c23 ),
    .o({\u2_Display/add101/c24 ,\u2_Display/n3260 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u24  (
    .a(\u2_Display/n3233 ),
    .b(1'b1),
    .c(\u2_Display/add101/c24 ),
    .o({\u2_Display/add101/c25 ,\u2_Display/n3260 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u25  (
    .a(\u2_Display/n3232 ),
    .b(1'b1),
    .c(\u2_Display/add101/c25 ),
    .o({\u2_Display/add101/c26 ,\u2_Display/n3260 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u26  (
    .a(\u2_Display/n3231 ),
    .b(1'b1),
    .c(\u2_Display/add101/c26 ),
    .o({\u2_Display/add101/c27 ,\u2_Display/n3260 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u27  (
    .a(\u2_Display/n3230 ),
    .b(1'b1),
    .c(\u2_Display/add101/c27 ),
    .o({\u2_Display/add101/c28 ,\u2_Display/n3260 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u28  (
    .a(\u2_Display/n3229 ),
    .b(1'b1),
    .c(\u2_Display/add101/c28 ),
    .o({\u2_Display/add101/c29 ,\u2_Display/n3260 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u29  (
    .a(\u2_Display/n3228 ),
    .b(1'b1),
    .c(\u2_Display/add101/c29 ),
    .o({\u2_Display/add101/c30 ,\u2_Display/n3260 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u3  (
    .a(\u2_Display/n3254 ),
    .b(1'b1),
    .c(\u2_Display/add101/c3 ),
    .o({\u2_Display/add101/c4 ,\u2_Display/n3260 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u30  (
    .a(\u2_Display/n3227 ),
    .b(1'b1),
    .c(\u2_Display/add101/c30 ),
    .o({\u2_Display/add101/c31 ,\u2_Display/n3260 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u31  (
    .a(\u2_Display/n3226 ),
    .b(1'b1),
    .c(\u2_Display/add101/c31 ),
    .o({open_n883,\u2_Display/n3260 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u4  (
    .a(\u2_Display/n3253 ),
    .b(1'b1),
    .c(\u2_Display/add101/c4 ),
    .o({\u2_Display/add101/c5 ,\u2_Display/n3260 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u5  (
    .a(\u2_Display/n3252 ),
    .b(1'b1),
    .c(\u2_Display/add101/c5 ),
    .o({\u2_Display/add101/c6 ,\u2_Display/n3260 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u6  (
    .a(\u2_Display/n3251 ),
    .b(1'b1),
    .c(\u2_Display/add101/c6 ),
    .o({\u2_Display/add101/c7 ,\u2_Display/n3260 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u7  (
    .a(\u2_Display/n3250 ),
    .b(1'b1),
    .c(\u2_Display/add101/c7 ),
    .o({\u2_Display/add101/c8 ,\u2_Display/n3260 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u8  (
    .a(\u2_Display/n3249 ),
    .b(1'b0),
    .c(\u2_Display/add101/c8 ),
    .o({\u2_Display/add101/c9 ,\u2_Display/n3260 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add101/u9  (
    .a(\u2_Display/n3248 ),
    .b(1'b0),
    .c(\u2_Display/add101/c9 ),
    .o({\u2_Display/add101/c10 ,\u2_Display/n3260 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add101/ucin  (
    .a(1'b1),
    .o({\u2_Display/add101/c0 ,open_n886}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u0  (
    .a(\u2_Display/n3292 ),
    .b(1'b1),
    .c(\u2_Display/add102/c0 ),
    .o({\u2_Display/add102/c1 ,\u2_Display/n3295 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u1  (
    .a(\u2_Display/n3291 ),
    .b(1'b1),
    .c(\u2_Display/add102/c1 ),
    .o({\u2_Display/add102/c2 ,\u2_Display/n3295 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u10  (
    .a(\u2_Display/n3282 ),
    .b(1'b0),
    .c(\u2_Display/add102/c10 ),
    .o({\u2_Display/add102/c11 ,\u2_Display/n3295 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u11  (
    .a(\u2_Display/n3281 ),
    .b(1'b1),
    .c(\u2_Display/add102/c11 ),
    .o({\u2_Display/add102/c12 ,\u2_Display/n3295 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u12  (
    .a(\u2_Display/n3280 ),
    .b(1'b1),
    .c(\u2_Display/add102/c12 ),
    .o({\u2_Display/add102/c13 ,\u2_Display/n3295 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u13  (
    .a(\u2_Display/n3279 ),
    .b(1'b0),
    .c(\u2_Display/add102/c13 ),
    .o({\u2_Display/add102/c14 ,\u2_Display/n3295 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u14  (
    .a(\u2_Display/n3278 ),
    .b(1'b1),
    .c(\u2_Display/add102/c14 ),
    .o({\u2_Display/add102/c15 ,\u2_Display/n3295 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u15  (
    .a(\u2_Display/n3277 ),
    .b(1'b1),
    .c(\u2_Display/add102/c15 ),
    .o({\u2_Display/add102/c16 ,\u2_Display/n3295 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u16  (
    .a(\u2_Display/n3276 ),
    .b(1'b1),
    .c(\u2_Display/add102/c16 ),
    .o({\u2_Display/add102/c17 ,\u2_Display/n3295 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u17  (
    .a(\u2_Display/n3275 ),
    .b(1'b1),
    .c(\u2_Display/add102/c17 ),
    .o({\u2_Display/add102/c18 ,\u2_Display/n3295 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u18  (
    .a(\u2_Display/n3274 ),
    .b(1'b1),
    .c(\u2_Display/add102/c18 ),
    .o({\u2_Display/add102/c19 ,\u2_Display/n3295 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u19  (
    .a(\u2_Display/n3273 ),
    .b(1'b1),
    .c(\u2_Display/add102/c19 ),
    .o({\u2_Display/add102/c20 ,\u2_Display/n3295 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u2  (
    .a(\u2_Display/n3290 ),
    .b(1'b1),
    .c(\u2_Display/add102/c2 ),
    .o({\u2_Display/add102/c3 ,\u2_Display/n3295 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u20  (
    .a(\u2_Display/n3272 ),
    .b(1'b1),
    .c(\u2_Display/add102/c20 ),
    .o({\u2_Display/add102/c21 ,\u2_Display/n3295 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u21  (
    .a(\u2_Display/n3271 ),
    .b(1'b1),
    .c(\u2_Display/add102/c21 ),
    .o({\u2_Display/add102/c22 ,\u2_Display/n3295 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u22  (
    .a(\u2_Display/n3270 ),
    .b(1'b1),
    .c(\u2_Display/add102/c22 ),
    .o({\u2_Display/add102/c23 ,\u2_Display/n3295 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u23  (
    .a(\u2_Display/n3269 ),
    .b(1'b1),
    .c(\u2_Display/add102/c23 ),
    .o({\u2_Display/add102/c24 ,\u2_Display/n3295 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u24  (
    .a(\u2_Display/n3268 ),
    .b(1'b1),
    .c(\u2_Display/add102/c24 ),
    .o({\u2_Display/add102/c25 ,\u2_Display/n3295 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u25  (
    .a(\u2_Display/n3267 ),
    .b(1'b1),
    .c(\u2_Display/add102/c25 ),
    .o({\u2_Display/add102/c26 ,\u2_Display/n3295 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u26  (
    .a(\u2_Display/n3266 ),
    .b(1'b1),
    .c(\u2_Display/add102/c26 ),
    .o({\u2_Display/add102/c27 ,\u2_Display/n3295 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u27  (
    .a(\u2_Display/n3265 ),
    .b(1'b1),
    .c(\u2_Display/add102/c27 ),
    .o({\u2_Display/add102/c28 ,\u2_Display/n3295 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u28  (
    .a(\u2_Display/n3264 ),
    .b(1'b1),
    .c(\u2_Display/add102/c28 ),
    .o({\u2_Display/add102/c29 ,\u2_Display/n3295 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u29  (
    .a(\u2_Display/n3263 ),
    .b(1'b1),
    .c(\u2_Display/add102/c29 ),
    .o({\u2_Display/add102/c30 ,\u2_Display/n3295 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u3  (
    .a(\u2_Display/n3289 ),
    .b(1'b1),
    .c(\u2_Display/add102/c3 ),
    .o({\u2_Display/add102/c4 ,\u2_Display/n3295 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u30  (
    .a(\u2_Display/n3262 ),
    .b(1'b1),
    .c(\u2_Display/add102/c30 ),
    .o({\u2_Display/add102/c31 ,\u2_Display/n3295 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u31  (
    .a(\u2_Display/n3261 ),
    .b(1'b1),
    .c(\u2_Display/add102/c31 ),
    .o({open_n887,\u2_Display/n3295 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u4  (
    .a(\u2_Display/n3288 ),
    .b(1'b1),
    .c(\u2_Display/add102/c4 ),
    .o({\u2_Display/add102/c5 ,\u2_Display/n3295 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u5  (
    .a(\u2_Display/n3287 ),
    .b(1'b1),
    .c(\u2_Display/add102/c5 ),
    .o({\u2_Display/add102/c6 ,\u2_Display/n3295 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u6  (
    .a(\u2_Display/n3286 ),
    .b(1'b1),
    .c(\u2_Display/add102/c6 ),
    .o({\u2_Display/add102/c7 ,\u2_Display/n3295 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u7  (
    .a(\u2_Display/n3285 ),
    .b(1'b0),
    .c(\u2_Display/add102/c7 ),
    .o({\u2_Display/add102/c8 ,\u2_Display/n3295 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u8  (
    .a(\u2_Display/n3284 ),
    .b(1'b0),
    .c(\u2_Display/add102/c8 ),
    .o({\u2_Display/add102/c9 ,\u2_Display/n3295 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add102/u9  (
    .a(\u2_Display/n3283 ),
    .b(1'b1),
    .c(\u2_Display/add102/c9 ),
    .o({\u2_Display/add102/c10 ,\u2_Display/n3295 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add102/ucin  (
    .a(1'b1),
    .o({\u2_Display/add102/c0 ,open_n890}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u0  (
    .a(\u2_Display/n3327 ),
    .b(1'b1),
    .c(\u2_Display/add103/c0 ),
    .o({\u2_Display/add103/c1 ,\u2_Display/n3330 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u1  (
    .a(\u2_Display/n3326 ),
    .b(1'b1),
    .c(\u2_Display/add103/c1 ),
    .o({\u2_Display/add103/c2 ,\u2_Display/n3330 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u10  (
    .a(\u2_Display/n3317 ),
    .b(1'b1),
    .c(\u2_Display/add103/c10 ),
    .o({\u2_Display/add103/c11 ,\u2_Display/n3330 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u11  (
    .a(\u2_Display/n3316 ),
    .b(1'b1),
    .c(\u2_Display/add103/c11 ),
    .o({\u2_Display/add103/c12 ,\u2_Display/n3330 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u12  (
    .a(\u2_Display/n3315 ),
    .b(1'b0),
    .c(\u2_Display/add103/c12 ),
    .o({\u2_Display/add103/c13 ,\u2_Display/n3330 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u13  (
    .a(\u2_Display/n3314 ),
    .b(1'b1),
    .c(\u2_Display/add103/c13 ),
    .o({\u2_Display/add103/c14 ,\u2_Display/n3330 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u14  (
    .a(\u2_Display/n3313 ),
    .b(1'b1),
    .c(\u2_Display/add103/c14 ),
    .o({\u2_Display/add103/c15 ,\u2_Display/n3330 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u15  (
    .a(\u2_Display/n3312 ),
    .b(1'b1),
    .c(\u2_Display/add103/c15 ),
    .o({\u2_Display/add103/c16 ,\u2_Display/n3330 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u16  (
    .a(\u2_Display/n3311 ),
    .b(1'b1),
    .c(\u2_Display/add103/c16 ),
    .o({\u2_Display/add103/c17 ,\u2_Display/n3330 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u17  (
    .a(\u2_Display/n3310 ),
    .b(1'b1),
    .c(\u2_Display/add103/c17 ),
    .o({\u2_Display/add103/c18 ,\u2_Display/n3330 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u18  (
    .a(\u2_Display/n3309 ),
    .b(1'b1),
    .c(\u2_Display/add103/c18 ),
    .o({\u2_Display/add103/c19 ,\u2_Display/n3330 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u19  (
    .a(\u2_Display/n3308 ),
    .b(1'b1),
    .c(\u2_Display/add103/c19 ),
    .o({\u2_Display/add103/c20 ,\u2_Display/n3330 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u2  (
    .a(\u2_Display/n3325 ),
    .b(1'b1),
    .c(\u2_Display/add103/c2 ),
    .o({\u2_Display/add103/c3 ,\u2_Display/n3330 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u20  (
    .a(\u2_Display/n3307 ),
    .b(1'b1),
    .c(\u2_Display/add103/c20 ),
    .o({\u2_Display/add103/c21 ,\u2_Display/n3330 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u21  (
    .a(\u2_Display/n3306 ),
    .b(1'b1),
    .c(\u2_Display/add103/c21 ),
    .o({\u2_Display/add103/c22 ,\u2_Display/n3330 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u22  (
    .a(\u2_Display/n3305 ),
    .b(1'b1),
    .c(\u2_Display/add103/c22 ),
    .o({\u2_Display/add103/c23 ,\u2_Display/n3330 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u23  (
    .a(\u2_Display/n3304 ),
    .b(1'b1),
    .c(\u2_Display/add103/c23 ),
    .o({\u2_Display/add103/c24 ,\u2_Display/n3330 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u24  (
    .a(\u2_Display/n3303 ),
    .b(1'b1),
    .c(\u2_Display/add103/c24 ),
    .o({\u2_Display/add103/c25 ,\u2_Display/n3330 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u25  (
    .a(\u2_Display/n3302 ),
    .b(1'b1),
    .c(\u2_Display/add103/c25 ),
    .o({\u2_Display/add103/c26 ,\u2_Display/n3330 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u26  (
    .a(\u2_Display/n3301 ),
    .b(1'b1),
    .c(\u2_Display/add103/c26 ),
    .o({\u2_Display/add103/c27 ,\u2_Display/n3330 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u27  (
    .a(\u2_Display/n3300 ),
    .b(1'b1),
    .c(\u2_Display/add103/c27 ),
    .o({\u2_Display/add103/c28 ,\u2_Display/n3330 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u28  (
    .a(\u2_Display/n3299 ),
    .b(1'b1),
    .c(\u2_Display/add103/c28 ),
    .o({\u2_Display/add103/c29 ,\u2_Display/n3330 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u29  (
    .a(\u2_Display/n3298 ),
    .b(1'b1),
    .c(\u2_Display/add103/c29 ),
    .o({\u2_Display/add103/c30 ,\u2_Display/n3330 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u3  (
    .a(\u2_Display/n3324 ),
    .b(1'b1),
    .c(\u2_Display/add103/c3 ),
    .o({\u2_Display/add103/c4 ,\u2_Display/n3330 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u30  (
    .a(\u2_Display/n3297 ),
    .b(1'b1),
    .c(\u2_Display/add103/c30 ),
    .o({\u2_Display/add103/c31 ,\u2_Display/n3330 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u31  (
    .a(\u2_Display/n3296 ),
    .b(1'b1),
    .c(\u2_Display/add103/c31 ),
    .o({open_n891,\u2_Display/n3330 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u4  (
    .a(\u2_Display/n3323 ),
    .b(1'b1),
    .c(\u2_Display/add103/c4 ),
    .o({\u2_Display/add103/c5 ,\u2_Display/n3330 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u5  (
    .a(\u2_Display/n3322 ),
    .b(1'b1),
    .c(\u2_Display/add103/c5 ),
    .o({\u2_Display/add103/c6 ,\u2_Display/n3330 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u6  (
    .a(\u2_Display/n3321 ),
    .b(1'b0),
    .c(\u2_Display/add103/c6 ),
    .o({\u2_Display/add103/c7 ,\u2_Display/n3330 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u7  (
    .a(\u2_Display/n3320 ),
    .b(1'b0),
    .c(\u2_Display/add103/c7 ),
    .o({\u2_Display/add103/c8 ,\u2_Display/n3330 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u8  (
    .a(\u2_Display/n3319 ),
    .b(1'b1),
    .c(\u2_Display/add103/c8 ),
    .o({\u2_Display/add103/c9 ,\u2_Display/n3330 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add103/u9  (
    .a(\u2_Display/n3318 ),
    .b(1'b0),
    .c(\u2_Display/add103/c9 ),
    .o({\u2_Display/add103/c10 ,\u2_Display/n3330 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add103/ucin  (
    .a(1'b1),
    .o({\u2_Display/add103/c0 ,open_n894}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u0  (
    .a(\u2_Display/n3362 ),
    .b(1'b1),
    .c(\u2_Display/add104/c0 ),
    .o({\u2_Display/add104/c1 ,\u2_Display/n3365 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u1  (
    .a(\u2_Display/n3361 ),
    .b(1'b1),
    .c(\u2_Display/add104/c1 ),
    .o({\u2_Display/add104/c2 ,\u2_Display/n3365 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u10  (
    .a(\u2_Display/n3352 ),
    .b(1'b1),
    .c(\u2_Display/add104/c10 ),
    .o({\u2_Display/add104/c11 ,\u2_Display/n3365 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u11  (
    .a(\u2_Display/n3351 ),
    .b(1'b0),
    .c(\u2_Display/add104/c11 ),
    .o({\u2_Display/add104/c12 ,\u2_Display/n3365 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u12  (
    .a(\u2_Display/n3350 ),
    .b(1'b1),
    .c(\u2_Display/add104/c12 ),
    .o({\u2_Display/add104/c13 ,\u2_Display/n3365 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u13  (
    .a(\u2_Display/n3349 ),
    .b(1'b1),
    .c(\u2_Display/add104/c13 ),
    .o({\u2_Display/add104/c14 ,\u2_Display/n3365 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u14  (
    .a(\u2_Display/n3348 ),
    .b(1'b1),
    .c(\u2_Display/add104/c14 ),
    .o({\u2_Display/add104/c15 ,\u2_Display/n3365 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u15  (
    .a(\u2_Display/n3347 ),
    .b(1'b1),
    .c(\u2_Display/add104/c15 ),
    .o({\u2_Display/add104/c16 ,\u2_Display/n3365 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u16  (
    .a(\u2_Display/n3346 ),
    .b(1'b1),
    .c(\u2_Display/add104/c16 ),
    .o({\u2_Display/add104/c17 ,\u2_Display/n3365 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u17  (
    .a(\u2_Display/n3345 ),
    .b(1'b1),
    .c(\u2_Display/add104/c17 ),
    .o({\u2_Display/add104/c18 ,\u2_Display/n3365 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u18  (
    .a(\u2_Display/n3344 ),
    .b(1'b1),
    .c(\u2_Display/add104/c18 ),
    .o({\u2_Display/add104/c19 ,\u2_Display/n3365 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u19  (
    .a(\u2_Display/n3343 ),
    .b(1'b1),
    .c(\u2_Display/add104/c19 ),
    .o({\u2_Display/add104/c20 ,\u2_Display/n3365 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u2  (
    .a(\u2_Display/n3360 ),
    .b(1'b1),
    .c(\u2_Display/add104/c2 ),
    .o({\u2_Display/add104/c3 ,\u2_Display/n3365 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u20  (
    .a(\u2_Display/n3342 ),
    .b(1'b1),
    .c(\u2_Display/add104/c20 ),
    .o({\u2_Display/add104/c21 ,\u2_Display/n3365 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u21  (
    .a(\u2_Display/n3341 ),
    .b(1'b1),
    .c(\u2_Display/add104/c21 ),
    .o({\u2_Display/add104/c22 ,\u2_Display/n3365 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u22  (
    .a(\u2_Display/n3340 ),
    .b(1'b1),
    .c(\u2_Display/add104/c22 ),
    .o({\u2_Display/add104/c23 ,\u2_Display/n3365 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u23  (
    .a(\u2_Display/n3339 ),
    .b(1'b1),
    .c(\u2_Display/add104/c23 ),
    .o({\u2_Display/add104/c24 ,\u2_Display/n3365 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u24  (
    .a(\u2_Display/n3338 ),
    .b(1'b1),
    .c(\u2_Display/add104/c24 ),
    .o({\u2_Display/add104/c25 ,\u2_Display/n3365 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u25  (
    .a(\u2_Display/n3337 ),
    .b(1'b1),
    .c(\u2_Display/add104/c25 ),
    .o({\u2_Display/add104/c26 ,\u2_Display/n3365 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u26  (
    .a(\u2_Display/n3336 ),
    .b(1'b1),
    .c(\u2_Display/add104/c26 ),
    .o({\u2_Display/add104/c27 ,\u2_Display/n3365 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u27  (
    .a(\u2_Display/n3335 ),
    .b(1'b1),
    .c(\u2_Display/add104/c27 ),
    .o({\u2_Display/add104/c28 ,\u2_Display/n3365 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u28  (
    .a(\u2_Display/n3334 ),
    .b(1'b1),
    .c(\u2_Display/add104/c28 ),
    .o({\u2_Display/add104/c29 ,\u2_Display/n3365 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u29  (
    .a(\u2_Display/n3333 ),
    .b(1'b1),
    .c(\u2_Display/add104/c29 ),
    .o({\u2_Display/add104/c30 ,\u2_Display/n3365 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u3  (
    .a(\u2_Display/n3359 ),
    .b(1'b1),
    .c(\u2_Display/add104/c3 ),
    .o({\u2_Display/add104/c4 ,\u2_Display/n3365 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u30  (
    .a(\u2_Display/n3332 ),
    .b(1'b1),
    .c(\u2_Display/add104/c30 ),
    .o({\u2_Display/add104/c31 ,\u2_Display/n3365 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u31  (
    .a(\u2_Display/n3331 ),
    .b(1'b1),
    .c(\u2_Display/add104/c31 ),
    .o({open_n895,\u2_Display/n3365 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u4  (
    .a(\u2_Display/n3358 ),
    .b(1'b1),
    .c(\u2_Display/add104/c4 ),
    .o({\u2_Display/add104/c5 ,\u2_Display/n3365 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u5  (
    .a(\u2_Display/n3357 ),
    .b(1'b0),
    .c(\u2_Display/add104/c5 ),
    .o({\u2_Display/add104/c6 ,\u2_Display/n3365 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u6  (
    .a(\u2_Display/n3356 ),
    .b(1'b0),
    .c(\u2_Display/add104/c6 ),
    .o({\u2_Display/add104/c7 ,\u2_Display/n3365 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u7  (
    .a(\u2_Display/n3355 ),
    .b(1'b1),
    .c(\u2_Display/add104/c7 ),
    .o({\u2_Display/add104/c8 ,\u2_Display/n3365 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u8  (
    .a(\u2_Display/n3354 ),
    .b(1'b0),
    .c(\u2_Display/add104/c8 ),
    .o({\u2_Display/add104/c9 ,\u2_Display/n3365 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add104/u9  (
    .a(\u2_Display/n3353 ),
    .b(1'b1),
    .c(\u2_Display/add104/c9 ),
    .o({\u2_Display/add104/c10 ,\u2_Display/n3365 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add104/ucin  (
    .a(1'b1),
    .o({\u2_Display/add104/c0 ,open_n898}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u0  (
    .a(\u2_Display/n3397 ),
    .b(1'b1),
    .c(\u2_Display/add105/c0 ),
    .o({\u2_Display/add105/c1 ,\u2_Display/n3400 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u1  (
    .a(\u2_Display/n3396 ),
    .b(1'b1),
    .c(\u2_Display/add105/c1 ),
    .o({\u2_Display/add105/c2 ,\u2_Display/n3400 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u10  (
    .a(\u2_Display/n3387 ),
    .b(1'b0),
    .c(\u2_Display/add105/c10 ),
    .o({\u2_Display/add105/c11 ,\u2_Display/n3400 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u11  (
    .a(\u2_Display/n3386 ),
    .b(1'b1),
    .c(\u2_Display/add105/c11 ),
    .o({\u2_Display/add105/c12 ,\u2_Display/n3400 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u12  (
    .a(\u2_Display/n3385 ),
    .b(1'b1),
    .c(\u2_Display/add105/c12 ),
    .o({\u2_Display/add105/c13 ,\u2_Display/n3400 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u13  (
    .a(\u2_Display/n3384 ),
    .b(1'b1),
    .c(\u2_Display/add105/c13 ),
    .o({\u2_Display/add105/c14 ,\u2_Display/n3400 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u14  (
    .a(\u2_Display/n3383 ),
    .b(1'b1),
    .c(\u2_Display/add105/c14 ),
    .o({\u2_Display/add105/c15 ,\u2_Display/n3400 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u15  (
    .a(\u2_Display/n3382 ),
    .b(1'b1),
    .c(\u2_Display/add105/c15 ),
    .o({\u2_Display/add105/c16 ,\u2_Display/n3400 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u16  (
    .a(\u2_Display/n3381 ),
    .b(1'b1),
    .c(\u2_Display/add105/c16 ),
    .o({\u2_Display/add105/c17 ,\u2_Display/n3400 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u17  (
    .a(\u2_Display/n3380 ),
    .b(1'b1),
    .c(\u2_Display/add105/c17 ),
    .o({\u2_Display/add105/c18 ,\u2_Display/n3400 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u18  (
    .a(\u2_Display/n3379 ),
    .b(1'b1),
    .c(\u2_Display/add105/c18 ),
    .o({\u2_Display/add105/c19 ,\u2_Display/n3400 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u19  (
    .a(\u2_Display/n3378 ),
    .b(1'b1),
    .c(\u2_Display/add105/c19 ),
    .o({\u2_Display/add105/c20 ,\u2_Display/n3400 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u2  (
    .a(\u2_Display/n3395 ),
    .b(1'b1),
    .c(\u2_Display/add105/c2 ),
    .o({\u2_Display/add105/c3 ,\u2_Display/n3400 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u20  (
    .a(\u2_Display/n3377 ),
    .b(1'b1),
    .c(\u2_Display/add105/c20 ),
    .o({\u2_Display/add105/c21 ,\u2_Display/n3400 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u21  (
    .a(\u2_Display/n3376 ),
    .b(1'b1),
    .c(\u2_Display/add105/c21 ),
    .o({\u2_Display/add105/c22 ,\u2_Display/n3400 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u22  (
    .a(\u2_Display/n3375 ),
    .b(1'b1),
    .c(\u2_Display/add105/c22 ),
    .o({\u2_Display/add105/c23 ,\u2_Display/n3400 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u23  (
    .a(\u2_Display/n3374 ),
    .b(1'b1),
    .c(\u2_Display/add105/c23 ),
    .o({\u2_Display/add105/c24 ,\u2_Display/n3400 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u24  (
    .a(\u2_Display/n3373 ),
    .b(1'b1),
    .c(\u2_Display/add105/c24 ),
    .o({\u2_Display/add105/c25 ,\u2_Display/n3400 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u25  (
    .a(\u2_Display/n3372 ),
    .b(1'b1),
    .c(\u2_Display/add105/c25 ),
    .o({\u2_Display/add105/c26 ,\u2_Display/n3400 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u26  (
    .a(\u2_Display/n3371 ),
    .b(1'b1),
    .c(\u2_Display/add105/c26 ),
    .o({\u2_Display/add105/c27 ,\u2_Display/n3400 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u27  (
    .a(\u2_Display/n3370 ),
    .b(1'b1),
    .c(\u2_Display/add105/c27 ),
    .o({\u2_Display/add105/c28 ,\u2_Display/n3400 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u28  (
    .a(\u2_Display/n3369 ),
    .b(1'b1),
    .c(\u2_Display/add105/c28 ),
    .o({\u2_Display/add105/c29 ,\u2_Display/n3400 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u29  (
    .a(\u2_Display/n3368 ),
    .b(1'b1),
    .c(\u2_Display/add105/c29 ),
    .o({\u2_Display/add105/c30 ,\u2_Display/n3400 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u3  (
    .a(\u2_Display/n3394 ),
    .b(1'b1),
    .c(\u2_Display/add105/c3 ),
    .o({\u2_Display/add105/c4 ,\u2_Display/n3400 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u30  (
    .a(\u2_Display/n3367 ),
    .b(1'b1),
    .c(\u2_Display/add105/c30 ),
    .o({\u2_Display/add105/c31 ,\u2_Display/n3400 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u31  (
    .a(\u2_Display/n3366 ),
    .b(1'b1),
    .c(\u2_Display/add105/c31 ),
    .o({open_n899,\u2_Display/n3400 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u4  (
    .a(\u2_Display/n3393 ),
    .b(1'b0),
    .c(\u2_Display/add105/c4 ),
    .o({\u2_Display/add105/c5 ,\u2_Display/n3400 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u5  (
    .a(\u2_Display/n3392 ),
    .b(1'b0),
    .c(\u2_Display/add105/c5 ),
    .o({\u2_Display/add105/c6 ,\u2_Display/n3400 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u6  (
    .a(\u2_Display/n3391 ),
    .b(1'b1),
    .c(\u2_Display/add105/c6 ),
    .o({\u2_Display/add105/c7 ,\u2_Display/n3400 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u7  (
    .a(\u2_Display/n3390 ),
    .b(1'b0),
    .c(\u2_Display/add105/c7 ),
    .o({\u2_Display/add105/c8 ,\u2_Display/n3400 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u8  (
    .a(\u2_Display/n3389 ),
    .b(1'b1),
    .c(\u2_Display/add105/c8 ),
    .o({\u2_Display/add105/c9 ,\u2_Display/n3400 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add105/u9  (
    .a(\u2_Display/n3388 ),
    .b(1'b1),
    .c(\u2_Display/add105/c9 ),
    .o({\u2_Display/add105/c10 ,\u2_Display/n3400 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add105/ucin  (
    .a(1'b1),
    .o({\u2_Display/add105/c0 ,open_n902}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add106/u0  (
    .a(\u2_Display/n3432 ),
    .b(1'b1),
    .c(\u2_Display/add106/c0 ),
    .o({\u2_Display/add106/c1 ,\u2_Display/n3435 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add106/u1  (
    .a(\u2_Display/n3431 ),
    .b(1'b1),
    .c(\u2_Display/add106/c1 ),
    .o({\u2_Display/add106/c2 ,\u2_Display/n3435 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add106/u2  (
    .a(\u2_Display/n3430 ),
    .b(1'b1),
    .c(\u2_Display/add106/c2 ),
    .o({\u2_Display/add106/c3 ,\u2_Display/n3435 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add106/u3  (
    .a(\u2_Display/n3429 ),
    .b(1'b0),
    .c(\u2_Display/add106/c3 ),
    .o({\u2_Display/add106/c4 ,\u2_Display/n3435 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add106/u4  (
    .a(\u2_Display/n3428 ),
    .b(1'b0),
    .c(\u2_Display/add106/c4 ),
    .o({\u2_Display/add106/c5 ,\u2_Display/n3435 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add106/u5  (
    .a(\u2_Display/n3427 ),
    .b(1'b1),
    .c(\u2_Display/add106/c5 ),
    .o({\u2_Display/add106/c6 ,\u2_Display/n3435 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add106/u6  (
    .a(\u2_Display/n3426 ),
    .b(1'b0),
    .c(\u2_Display/add106/c6 ),
    .o({\u2_Display/add106/c7 ,\u2_Display/n3435 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add106/u7  (
    .a(\u2_Display/n3425 ),
    .b(1'b1),
    .c(\u2_Display/add106/c7 ),
    .o({\u2_Display/add106/c8 ,\u2_Display/n3435 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add106/u8  (
    .a(\u2_Display/n3424 ),
    .b(1'b1),
    .c(\u2_Display/add106/c8 ),
    .o({\u2_Display/add106/c9 ,\u2_Display/n3435 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add106/u9  (
    .a(\u2_Display/n3423 ),
    .b(1'b0),
    .c(\u2_Display/add106/c9 ),
    .o({open_n903,\u2_Display/n3435 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add106/ucin  (
    .a(1'b1),
    .o({\u2_Display/add106/c0 ,open_n906}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u0  (
    .a(\u2_Display/counta [0]),
    .b(1'b1),
    .c(\u2_Display/add117/c0 ),
    .o({\u2_Display/add117/c1 ,\u2_Display/n3788 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u1  (
    .a(\u2_Display/counta [1]),
    .b(1'b1),
    .c(\u2_Display/add117/c1 ),
    .o({\u2_Display/add117/c2 ,\u2_Display/n3788 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u10  (
    .a(\u2_Display/counta [10]),
    .b(1'b1),
    .c(\u2_Display/add117/c10 ),
    .o({\u2_Display/add117/c11 ,\u2_Display/n3788 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u11  (
    .a(\u2_Display/counta [11]),
    .b(1'b1),
    .c(\u2_Display/add117/c11 ),
    .o({\u2_Display/add117/c12 ,\u2_Display/n3788 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u12  (
    .a(\u2_Display/counta [12]),
    .b(1'b1),
    .c(\u2_Display/add117/c12 ),
    .o({\u2_Display/add117/c13 ,\u2_Display/n3788 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u13  (
    .a(\u2_Display/counta [13]),
    .b(1'b1),
    .c(\u2_Display/add117/c13 ),
    .o({\u2_Display/add117/c14 ,\u2_Display/n3788 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u14  (
    .a(\u2_Display/counta [14]),
    .b(1'b1),
    .c(\u2_Display/add117/c14 ),
    .o({\u2_Display/add117/c15 ,\u2_Display/n3788 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u15  (
    .a(\u2_Display/counta [15]),
    .b(1'b1),
    .c(\u2_Display/add117/c15 ),
    .o({\u2_Display/add117/c16 ,\u2_Display/n3788 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u16  (
    .a(\u2_Display/counta [16]),
    .b(1'b1),
    .c(\u2_Display/add117/c16 ),
    .o({\u2_Display/add117/c17 ,\u2_Display/n3788 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u17  (
    .a(\u2_Display/counta [17]),
    .b(1'b1),
    .c(\u2_Display/add117/c17 ),
    .o({\u2_Display/add117/c18 ,\u2_Display/n3788 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u18  (
    .a(\u2_Display/counta [18]),
    .b(1'b1),
    .c(\u2_Display/add117/c18 ),
    .o({\u2_Display/add117/c19 ,\u2_Display/n3788 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u19  (
    .a(\u2_Display/counta [19]),
    .b(1'b1),
    .c(\u2_Display/add117/c19 ),
    .o({\u2_Display/add117/c20 ,\u2_Display/n3788 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u2  (
    .a(\u2_Display/counta [2]),
    .b(1'b1),
    .c(\u2_Display/add117/c2 ),
    .o({\u2_Display/add117/c3 ,\u2_Display/n3788 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u20  (
    .a(\u2_Display/counta [20]),
    .b(1'b1),
    .c(\u2_Display/add117/c20 ),
    .o({\u2_Display/add117/c21 ,\u2_Display/n3788 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u21  (
    .a(\u2_Display/counta [21]),
    .b(1'b1),
    .c(\u2_Display/add117/c21 ),
    .o({\u2_Display/add117/c22 ,\u2_Display/n3788 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u22  (
    .a(\u2_Display/counta [22]),
    .b(1'b1),
    .c(\u2_Display/add117/c22 ),
    .o({\u2_Display/add117/c23 ,\u2_Display/n3788 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u23  (
    .a(\u2_Display/counta [23]),
    .b(1'b1),
    .c(\u2_Display/add117/c23 ),
    .o({\u2_Display/add117/c24 ,\u2_Display/n3788 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u24  (
    .a(\u2_Display/counta [24]),
    .b(1'b1),
    .c(\u2_Display/add117/c24 ),
    .o({\u2_Display/add117/c25 ,\u2_Display/n3788 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u25  (
    .a(\u2_Display/counta [25]),
    .b(1'b1),
    .c(\u2_Display/add117/c25 ),
    .o({\u2_Display/add117/c26 ,\u2_Display/n3788 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u26  (
    .a(\u2_Display/counta [26]),
    .b(1'b1),
    .c(\u2_Display/add117/c26 ),
    .o({\u2_Display/add117/c27 ,\u2_Display/n3788 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u27  (
    .a(\u2_Display/counta [27]),
    .b(1'b0),
    .c(\u2_Display/add117/c27 ),
    .o({\u2_Display/add117/c28 ,\u2_Display/n3788 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u28  (
    .a(\u2_Display/counta [28]),
    .b(1'b1),
    .c(\u2_Display/add117/c28 ),
    .o({\u2_Display/add117/c29 ,\u2_Display/n3788 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u29  (
    .a(\u2_Display/counta [29]),
    .b(1'b1),
    .c(\u2_Display/add117/c29 ),
    .o({\u2_Display/add117/c30 ,\u2_Display/n3788 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u3  (
    .a(\u2_Display/counta [3]),
    .b(1'b1),
    .c(\u2_Display/add117/c3 ),
    .o({\u2_Display/add117/c4 ,\u2_Display/n3788 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u30  (
    .a(\u2_Display/counta [30]),
    .b(1'b0),
    .c(\u2_Display/add117/c30 ),
    .o({\u2_Display/add117/c31 ,\u2_Display/n3788 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u31  (
    .a(\u2_Display/counta [31]),
    .b(1'b0),
    .c(\u2_Display/add117/c31 ),
    .o({open_n907,\u2_Display/n3788 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u4  (
    .a(\u2_Display/counta [4]),
    .b(1'b1),
    .c(\u2_Display/add117/c4 ),
    .o({\u2_Display/add117/c5 ,\u2_Display/n3788 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u5  (
    .a(\u2_Display/counta [5]),
    .b(1'b1),
    .c(\u2_Display/add117/c5 ),
    .o({\u2_Display/add117/c6 ,\u2_Display/n3788 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u6  (
    .a(\u2_Display/counta [6]),
    .b(1'b1),
    .c(\u2_Display/add117/c6 ),
    .o({\u2_Display/add117/c7 ,\u2_Display/n3788 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u7  (
    .a(\u2_Display/counta [7]),
    .b(1'b1),
    .c(\u2_Display/add117/c7 ),
    .o({\u2_Display/add117/c8 ,\u2_Display/n3788 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u8  (
    .a(\u2_Display/counta [8]),
    .b(1'b1),
    .c(\u2_Display/add117/c8 ),
    .o({\u2_Display/add117/c9 ,\u2_Display/n3788 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add117/u9  (
    .a(\u2_Display/counta [9]),
    .b(1'b1),
    .c(\u2_Display/add117/c9 ),
    .o({\u2_Display/add117/c10 ,\u2_Display/n3788 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add117/ucin  (
    .a(1'b1),
    .o({\u2_Display/add117/c0 ,open_n910}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u0  (
    .a(\u2_Display/n3820 ),
    .b(1'b1),
    .c(\u2_Display/add118/c0 ),
    .o({\u2_Display/add118/c1 ,\u2_Display/n3823 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u1  (
    .a(\u2_Display/n3819 ),
    .b(1'b1),
    .c(\u2_Display/add118/c1 ),
    .o({\u2_Display/add118/c2 ,\u2_Display/n3823 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u10  (
    .a(\u2_Display/n3810 ),
    .b(1'b1),
    .c(\u2_Display/add118/c10 ),
    .o({\u2_Display/add118/c11 ,\u2_Display/n3823 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u11  (
    .a(\u2_Display/n3809 ),
    .b(1'b1),
    .c(\u2_Display/add118/c11 ),
    .o({\u2_Display/add118/c12 ,\u2_Display/n3823 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u12  (
    .a(\u2_Display/n3808 ),
    .b(1'b1),
    .c(\u2_Display/add118/c12 ),
    .o({\u2_Display/add118/c13 ,\u2_Display/n3823 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u13  (
    .a(\u2_Display/n3807 ),
    .b(1'b1),
    .c(\u2_Display/add118/c13 ),
    .o({\u2_Display/add118/c14 ,\u2_Display/n3823 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u14  (
    .a(\u2_Display/n3806 ),
    .b(1'b1),
    .c(\u2_Display/add118/c14 ),
    .o({\u2_Display/add118/c15 ,\u2_Display/n3823 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u15  (
    .a(\u2_Display/n3805 ),
    .b(1'b1),
    .c(\u2_Display/add118/c15 ),
    .o({\u2_Display/add118/c16 ,\u2_Display/n3823 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u16  (
    .a(\u2_Display/n3804 ),
    .b(1'b1),
    .c(\u2_Display/add118/c16 ),
    .o({\u2_Display/add118/c17 ,\u2_Display/n3823 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u17  (
    .a(\u2_Display/n3803 ),
    .b(1'b1),
    .c(\u2_Display/add118/c17 ),
    .o({\u2_Display/add118/c18 ,\u2_Display/n3823 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u18  (
    .a(\u2_Display/n3802 ),
    .b(1'b1),
    .c(\u2_Display/add118/c18 ),
    .o({\u2_Display/add118/c19 ,\u2_Display/n3823 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u19  (
    .a(\u2_Display/n3801 ),
    .b(1'b1),
    .c(\u2_Display/add118/c19 ),
    .o({\u2_Display/add118/c20 ,\u2_Display/n3823 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u2  (
    .a(\u2_Display/n3818 ),
    .b(1'b1),
    .c(\u2_Display/add118/c2 ),
    .o({\u2_Display/add118/c3 ,\u2_Display/n3823 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u20  (
    .a(\u2_Display/n3800 ),
    .b(1'b1),
    .c(\u2_Display/add118/c20 ),
    .o({\u2_Display/add118/c21 ,\u2_Display/n3823 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u21  (
    .a(\u2_Display/n3799 ),
    .b(1'b1),
    .c(\u2_Display/add118/c21 ),
    .o({\u2_Display/add118/c22 ,\u2_Display/n3823 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u22  (
    .a(\u2_Display/n3798 ),
    .b(1'b1),
    .c(\u2_Display/add118/c22 ),
    .o({\u2_Display/add118/c23 ,\u2_Display/n3823 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u23  (
    .a(\u2_Display/n3797 ),
    .b(1'b1),
    .c(\u2_Display/add118/c23 ),
    .o({\u2_Display/add118/c24 ,\u2_Display/n3823 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u24  (
    .a(\u2_Display/n3796 ),
    .b(1'b1),
    .c(\u2_Display/add118/c24 ),
    .o({\u2_Display/add118/c25 ,\u2_Display/n3823 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u25  (
    .a(\u2_Display/n3795 ),
    .b(1'b1),
    .c(\u2_Display/add118/c25 ),
    .o({\u2_Display/add118/c26 ,\u2_Display/n3823 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u26  (
    .a(\u2_Display/n3794 ),
    .b(1'b0),
    .c(\u2_Display/add118/c26 ),
    .o({\u2_Display/add118/c27 ,\u2_Display/n3823 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u27  (
    .a(\u2_Display/n3793 ),
    .b(1'b1),
    .c(\u2_Display/add118/c27 ),
    .o({\u2_Display/add118/c28 ,\u2_Display/n3823 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u28  (
    .a(\u2_Display/n3792 ),
    .b(1'b1),
    .c(\u2_Display/add118/c28 ),
    .o({\u2_Display/add118/c29 ,\u2_Display/n3823 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u29  (
    .a(\u2_Display/n3791 ),
    .b(1'b0),
    .c(\u2_Display/add118/c29 ),
    .o({\u2_Display/add118/c30 ,\u2_Display/n3823 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u3  (
    .a(\u2_Display/n3817 ),
    .b(1'b1),
    .c(\u2_Display/add118/c3 ),
    .o({\u2_Display/add118/c4 ,\u2_Display/n3823 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u30  (
    .a(\u2_Display/n3790 ),
    .b(1'b0),
    .c(\u2_Display/add118/c30 ),
    .o({\u2_Display/add118/c31 ,\u2_Display/n3823 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u31  (
    .a(\u2_Display/n3789 ),
    .b(1'b1),
    .c(\u2_Display/add118/c31 ),
    .o({open_n911,\u2_Display/n3823 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u4  (
    .a(\u2_Display/n3816 ),
    .b(1'b1),
    .c(\u2_Display/add118/c4 ),
    .o({\u2_Display/add118/c5 ,\u2_Display/n3823 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u5  (
    .a(\u2_Display/n3815 ),
    .b(1'b1),
    .c(\u2_Display/add118/c5 ),
    .o({\u2_Display/add118/c6 ,\u2_Display/n3823 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u6  (
    .a(\u2_Display/n3814 ),
    .b(1'b1),
    .c(\u2_Display/add118/c6 ),
    .o({\u2_Display/add118/c7 ,\u2_Display/n3823 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u7  (
    .a(\u2_Display/n3813 ),
    .b(1'b1),
    .c(\u2_Display/add118/c7 ),
    .o({\u2_Display/add118/c8 ,\u2_Display/n3823 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u8  (
    .a(\u2_Display/n3812 ),
    .b(1'b1),
    .c(\u2_Display/add118/c8 ),
    .o({\u2_Display/add118/c9 ,\u2_Display/n3823 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add118/u9  (
    .a(\u2_Display/n3811 ),
    .b(1'b1),
    .c(\u2_Display/add118/c9 ),
    .o({\u2_Display/add118/c10 ,\u2_Display/n3823 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add118/ucin  (
    .a(1'b1),
    .o({\u2_Display/add118/c0 ,open_n914}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u0  (
    .a(\u2_Display/n3855 ),
    .b(1'b1),
    .c(\u2_Display/add119/c0 ),
    .o({\u2_Display/add119/c1 ,\u2_Display/n3858 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u1  (
    .a(\u2_Display/n3854 ),
    .b(1'b1),
    .c(\u2_Display/add119/c1 ),
    .o({\u2_Display/add119/c2 ,\u2_Display/n3858 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u10  (
    .a(\u2_Display/n3845 ),
    .b(1'b1),
    .c(\u2_Display/add119/c10 ),
    .o({\u2_Display/add119/c11 ,\u2_Display/n3858 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u11  (
    .a(\u2_Display/n3844 ),
    .b(1'b1),
    .c(\u2_Display/add119/c11 ),
    .o({\u2_Display/add119/c12 ,\u2_Display/n3858 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u12  (
    .a(\u2_Display/n3843 ),
    .b(1'b1),
    .c(\u2_Display/add119/c12 ),
    .o({\u2_Display/add119/c13 ,\u2_Display/n3858 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u13  (
    .a(\u2_Display/n3842 ),
    .b(1'b1),
    .c(\u2_Display/add119/c13 ),
    .o({\u2_Display/add119/c14 ,\u2_Display/n3858 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u14  (
    .a(\u2_Display/n3841 ),
    .b(1'b1),
    .c(\u2_Display/add119/c14 ),
    .o({\u2_Display/add119/c15 ,\u2_Display/n3858 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u15  (
    .a(\u2_Display/n3840 ),
    .b(1'b1),
    .c(\u2_Display/add119/c15 ),
    .o({\u2_Display/add119/c16 ,\u2_Display/n3858 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u16  (
    .a(\u2_Display/n3839 ),
    .b(1'b1),
    .c(\u2_Display/add119/c16 ),
    .o({\u2_Display/add119/c17 ,\u2_Display/n3858 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u17  (
    .a(\u2_Display/n3838 ),
    .b(1'b1),
    .c(\u2_Display/add119/c17 ),
    .o({\u2_Display/add119/c18 ,\u2_Display/n3858 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u18  (
    .a(\u2_Display/n3837 ),
    .b(1'b1),
    .c(\u2_Display/add119/c18 ),
    .o({\u2_Display/add119/c19 ,\u2_Display/n3858 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u19  (
    .a(\u2_Display/n3836 ),
    .b(1'b1),
    .c(\u2_Display/add119/c19 ),
    .o({\u2_Display/add119/c20 ,\u2_Display/n3858 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u2  (
    .a(\u2_Display/n3853 ),
    .b(1'b1),
    .c(\u2_Display/add119/c2 ),
    .o({\u2_Display/add119/c3 ,\u2_Display/n3858 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u20  (
    .a(\u2_Display/n3835 ),
    .b(1'b1),
    .c(\u2_Display/add119/c20 ),
    .o({\u2_Display/add119/c21 ,\u2_Display/n3858 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u21  (
    .a(\u2_Display/n3834 ),
    .b(1'b1),
    .c(\u2_Display/add119/c21 ),
    .o({\u2_Display/add119/c22 ,\u2_Display/n3858 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u22  (
    .a(\u2_Display/n3833 ),
    .b(1'b1),
    .c(\u2_Display/add119/c22 ),
    .o({\u2_Display/add119/c23 ,\u2_Display/n3858 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u23  (
    .a(\u2_Display/n3832 ),
    .b(1'b1),
    .c(\u2_Display/add119/c23 ),
    .o({\u2_Display/add119/c24 ,\u2_Display/n3858 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u24  (
    .a(\u2_Display/n3831 ),
    .b(1'b1),
    .c(\u2_Display/add119/c24 ),
    .o({\u2_Display/add119/c25 ,\u2_Display/n3858 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u25  (
    .a(\u2_Display/n3830 ),
    .b(1'b0),
    .c(\u2_Display/add119/c25 ),
    .o({\u2_Display/add119/c26 ,\u2_Display/n3858 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u26  (
    .a(\u2_Display/n3829 ),
    .b(1'b1),
    .c(\u2_Display/add119/c26 ),
    .o({\u2_Display/add119/c27 ,\u2_Display/n3858 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u27  (
    .a(\u2_Display/n3828 ),
    .b(1'b1),
    .c(\u2_Display/add119/c27 ),
    .o({\u2_Display/add119/c28 ,\u2_Display/n3858 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u28  (
    .a(\u2_Display/n3827 ),
    .b(1'b0),
    .c(\u2_Display/add119/c28 ),
    .o({\u2_Display/add119/c29 ,\u2_Display/n3858 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u29  (
    .a(\u2_Display/n3826 ),
    .b(1'b0),
    .c(\u2_Display/add119/c29 ),
    .o({\u2_Display/add119/c30 ,\u2_Display/n3858 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u3  (
    .a(\u2_Display/n3852 ),
    .b(1'b1),
    .c(\u2_Display/add119/c3 ),
    .o({\u2_Display/add119/c4 ,\u2_Display/n3858 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u30  (
    .a(\u2_Display/n3825 ),
    .b(1'b1),
    .c(\u2_Display/add119/c30 ),
    .o({\u2_Display/add119/c31 ,\u2_Display/n3858 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u31  (
    .a(\u2_Display/n3824 ),
    .b(1'b1),
    .c(\u2_Display/add119/c31 ),
    .o({open_n915,\u2_Display/n3858 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u4  (
    .a(\u2_Display/n3851 ),
    .b(1'b1),
    .c(\u2_Display/add119/c4 ),
    .o({\u2_Display/add119/c5 ,\u2_Display/n3858 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u5  (
    .a(\u2_Display/n3850 ),
    .b(1'b1),
    .c(\u2_Display/add119/c5 ),
    .o({\u2_Display/add119/c6 ,\u2_Display/n3858 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u6  (
    .a(\u2_Display/n3849 ),
    .b(1'b1),
    .c(\u2_Display/add119/c6 ),
    .o({\u2_Display/add119/c7 ,\u2_Display/n3858 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u7  (
    .a(\u2_Display/n3848 ),
    .b(1'b1),
    .c(\u2_Display/add119/c7 ),
    .o({\u2_Display/add119/c8 ,\u2_Display/n3858 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u8  (
    .a(\u2_Display/n3847 ),
    .b(1'b1),
    .c(\u2_Display/add119/c8 ),
    .o({\u2_Display/add119/c9 ,\u2_Display/n3858 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add119/u9  (
    .a(\u2_Display/n3846 ),
    .b(1'b1),
    .c(\u2_Display/add119/c9 ),
    .o({\u2_Display/add119/c10 ,\u2_Display/n3858 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add119/ucin  (
    .a(1'b1),
    .o({\u2_Display/add119/c0 ,open_n918}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u0  (
    .a(\u2_Display/n3890 ),
    .b(1'b1),
    .c(\u2_Display/add120/c0 ),
    .o({\u2_Display/add120/c1 ,\u2_Display/n3893 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u1  (
    .a(\u2_Display/n3889 ),
    .b(1'b1),
    .c(\u2_Display/add120/c1 ),
    .o({\u2_Display/add120/c2 ,\u2_Display/n3893 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u10  (
    .a(\u2_Display/n3880 ),
    .b(1'b1),
    .c(\u2_Display/add120/c10 ),
    .o({\u2_Display/add120/c11 ,\u2_Display/n3893 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u11  (
    .a(\u2_Display/n3879 ),
    .b(1'b1),
    .c(\u2_Display/add120/c11 ),
    .o({\u2_Display/add120/c12 ,\u2_Display/n3893 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u12  (
    .a(\u2_Display/n3878 ),
    .b(1'b1),
    .c(\u2_Display/add120/c12 ),
    .o({\u2_Display/add120/c13 ,\u2_Display/n3893 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u13  (
    .a(\u2_Display/n3877 ),
    .b(1'b1),
    .c(\u2_Display/add120/c13 ),
    .o({\u2_Display/add120/c14 ,\u2_Display/n3893 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u14  (
    .a(\u2_Display/n3876 ),
    .b(1'b1),
    .c(\u2_Display/add120/c14 ),
    .o({\u2_Display/add120/c15 ,\u2_Display/n3893 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u15  (
    .a(\u2_Display/n3875 ),
    .b(1'b1),
    .c(\u2_Display/add120/c15 ),
    .o({\u2_Display/add120/c16 ,\u2_Display/n3893 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u16  (
    .a(\u2_Display/n3874 ),
    .b(1'b1),
    .c(\u2_Display/add120/c16 ),
    .o({\u2_Display/add120/c17 ,\u2_Display/n3893 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u17  (
    .a(\u2_Display/n3873 ),
    .b(1'b1),
    .c(\u2_Display/add120/c17 ),
    .o({\u2_Display/add120/c18 ,\u2_Display/n3893 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u18  (
    .a(\u2_Display/n3872 ),
    .b(1'b1),
    .c(\u2_Display/add120/c18 ),
    .o({\u2_Display/add120/c19 ,\u2_Display/n3893 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u19  (
    .a(\u2_Display/n3871 ),
    .b(1'b1),
    .c(\u2_Display/add120/c19 ),
    .o({\u2_Display/add120/c20 ,\u2_Display/n3893 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u2  (
    .a(\u2_Display/n3888 ),
    .b(1'b1),
    .c(\u2_Display/add120/c2 ),
    .o({\u2_Display/add120/c3 ,\u2_Display/n3893 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u20  (
    .a(\u2_Display/n3870 ),
    .b(1'b1),
    .c(\u2_Display/add120/c20 ),
    .o({\u2_Display/add120/c21 ,\u2_Display/n3893 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u21  (
    .a(\u2_Display/n3869 ),
    .b(1'b1),
    .c(\u2_Display/add120/c21 ),
    .o({\u2_Display/add120/c22 ,\u2_Display/n3893 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u22  (
    .a(\u2_Display/n3868 ),
    .b(1'b1),
    .c(\u2_Display/add120/c22 ),
    .o({\u2_Display/add120/c23 ,\u2_Display/n3893 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u23  (
    .a(\u2_Display/n3867 ),
    .b(1'b1),
    .c(\u2_Display/add120/c23 ),
    .o({\u2_Display/add120/c24 ,\u2_Display/n3893 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u24  (
    .a(\u2_Display/n3866 ),
    .b(1'b0),
    .c(\u2_Display/add120/c24 ),
    .o({\u2_Display/add120/c25 ,\u2_Display/n3893 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u25  (
    .a(\u2_Display/n3865 ),
    .b(1'b1),
    .c(\u2_Display/add120/c25 ),
    .o({\u2_Display/add120/c26 ,\u2_Display/n3893 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u26  (
    .a(\u2_Display/n3864 ),
    .b(1'b1),
    .c(\u2_Display/add120/c26 ),
    .o({\u2_Display/add120/c27 ,\u2_Display/n3893 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u27  (
    .a(\u2_Display/n3863 ),
    .b(1'b0),
    .c(\u2_Display/add120/c27 ),
    .o({\u2_Display/add120/c28 ,\u2_Display/n3893 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u28  (
    .a(\u2_Display/n3862 ),
    .b(1'b0),
    .c(\u2_Display/add120/c28 ),
    .o({\u2_Display/add120/c29 ,\u2_Display/n3893 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u29  (
    .a(\u2_Display/n3861 ),
    .b(1'b1),
    .c(\u2_Display/add120/c29 ),
    .o({\u2_Display/add120/c30 ,\u2_Display/n3893 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u3  (
    .a(\u2_Display/n3887 ),
    .b(1'b1),
    .c(\u2_Display/add120/c3 ),
    .o({\u2_Display/add120/c4 ,\u2_Display/n3893 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u30  (
    .a(\u2_Display/n3860 ),
    .b(1'b1),
    .c(\u2_Display/add120/c30 ),
    .o({\u2_Display/add120/c31 ,\u2_Display/n3893 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u31  (
    .a(\u2_Display/n3859 ),
    .b(1'b1),
    .c(\u2_Display/add120/c31 ),
    .o({open_n919,\u2_Display/n3893 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u4  (
    .a(\u2_Display/n3886 ),
    .b(1'b1),
    .c(\u2_Display/add120/c4 ),
    .o({\u2_Display/add120/c5 ,\u2_Display/n3893 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u5  (
    .a(\u2_Display/n3885 ),
    .b(1'b1),
    .c(\u2_Display/add120/c5 ),
    .o({\u2_Display/add120/c6 ,\u2_Display/n3893 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u6  (
    .a(\u2_Display/n3884 ),
    .b(1'b1),
    .c(\u2_Display/add120/c6 ),
    .o({\u2_Display/add120/c7 ,\u2_Display/n3893 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u7  (
    .a(\u2_Display/n3883 ),
    .b(1'b1),
    .c(\u2_Display/add120/c7 ),
    .o({\u2_Display/add120/c8 ,\u2_Display/n3893 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u8  (
    .a(\u2_Display/n3882 ),
    .b(1'b1),
    .c(\u2_Display/add120/c8 ),
    .o({\u2_Display/add120/c9 ,\u2_Display/n3893 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add120/u9  (
    .a(\u2_Display/n3881 ),
    .b(1'b1),
    .c(\u2_Display/add120/c9 ),
    .o({\u2_Display/add120/c10 ,\u2_Display/n3893 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add120/ucin  (
    .a(1'b1),
    .o({\u2_Display/add120/c0 ,open_n922}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u0  (
    .a(\u2_Display/n3925 ),
    .b(1'b1),
    .c(\u2_Display/add121/c0 ),
    .o({\u2_Display/add121/c1 ,\u2_Display/n3928 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u1  (
    .a(\u2_Display/n3924 ),
    .b(1'b1),
    .c(\u2_Display/add121/c1 ),
    .o({\u2_Display/add121/c2 ,\u2_Display/n3928 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u10  (
    .a(\u2_Display/n3915 ),
    .b(1'b1),
    .c(\u2_Display/add121/c10 ),
    .o({\u2_Display/add121/c11 ,\u2_Display/n3928 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u11  (
    .a(\u2_Display/n3914 ),
    .b(1'b1),
    .c(\u2_Display/add121/c11 ),
    .o({\u2_Display/add121/c12 ,\u2_Display/n3928 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u12  (
    .a(\u2_Display/n3913 ),
    .b(1'b1),
    .c(\u2_Display/add121/c12 ),
    .o({\u2_Display/add121/c13 ,\u2_Display/n3928 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u13  (
    .a(\u2_Display/n3912 ),
    .b(1'b1),
    .c(\u2_Display/add121/c13 ),
    .o({\u2_Display/add121/c14 ,\u2_Display/n3928 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u14  (
    .a(\u2_Display/n3911 ),
    .b(1'b1),
    .c(\u2_Display/add121/c14 ),
    .o({\u2_Display/add121/c15 ,\u2_Display/n3928 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u15  (
    .a(\u2_Display/n3910 ),
    .b(1'b1),
    .c(\u2_Display/add121/c15 ),
    .o({\u2_Display/add121/c16 ,\u2_Display/n3928 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u16  (
    .a(\u2_Display/n3909 ),
    .b(1'b1),
    .c(\u2_Display/add121/c16 ),
    .o({\u2_Display/add121/c17 ,\u2_Display/n3928 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u17  (
    .a(\u2_Display/n3908 ),
    .b(1'b1),
    .c(\u2_Display/add121/c17 ),
    .o({\u2_Display/add121/c18 ,\u2_Display/n3928 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u18  (
    .a(\u2_Display/n3907 ),
    .b(1'b1),
    .c(\u2_Display/add121/c18 ),
    .o({\u2_Display/add121/c19 ,\u2_Display/n3928 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u19  (
    .a(\u2_Display/n3906 ),
    .b(1'b1),
    .c(\u2_Display/add121/c19 ),
    .o({\u2_Display/add121/c20 ,\u2_Display/n3928 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u2  (
    .a(\u2_Display/n3923 ),
    .b(1'b1),
    .c(\u2_Display/add121/c2 ),
    .o({\u2_Display/add121/c3 ,\u2_Display/n3928 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u20  (
    .a(\u2_Display/n3905 ),
    .b(1'b1),
    .c(\u2_Display/add121/c20 ),
    .o({\u2_Display/add121/c21 ,\u2_Display/n3928 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u21  (
    .a(\u2_Display/n3904 ),
    .b(1'b1),
    .c(\u2_Display/add121/c21 ),
    .o({\u2_Display/add121/c22 ,\u2_Display/n3928 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u22  (
    .a(\u2_Display/n3903 ),
    .b(1'b1),
    .c(\u2_Display/add121/c22 ),
    .o({\u2_Display/add121/c23 ,\u2_Display/n3928 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u23  (
    .a(\u2_Display/n3902 ),
    .b(1'b0),
    .c(\u2_Display/add121/c23 ),
    .o({\u2_Display/add121/c24 ,\u2_Display/n3928 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u24  (
    .a(\u2_Display/n3901 ),
    .b(1'b1),
    .c(\u2_Display/add121/c24 ),
    .o({\u2_Display/add121/c25 ,\u2_Display/n3928 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u25  (
    .a(\u2_Display/n3900 ),
    .b(1'b1),
    .c(\u2_Display/add121/c25 ),
    .o({\u2_Display/add121/c26 ,\u2_Display/n3928 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u26  (
    .a(\u2_Display/n3899 ),
    .b(1'b0),
    .c(\u2_Display/add121/c26 ),
    .o({\u2_Display/add121/c27 ,\u2_Display/n3928 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u27  (
    .a(\u2_Display/n3898 ),
    .b(1'b0),
    .c(\u2_Display/add121/c27 ),
    .o({\u2_Display/add121/c28 ,\u2_Display/n3928 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u28  (
    .a(\u2_Display/n3897 ),
    .b(1'b1),
    .c(\u2_Display/add121/c28 ),
    .o({\u2_Display/add121/c29 ,\u2_Display/n3928 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u29  (
    .a(\u2_Display/n3896 ),
    .b(1'b1),
    .c(\u2_Display/add121/c29 ),
    .o({\u2_Display/add121/c30 ,\u2_Display/n3928 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u3  (
    .a(\u2_Display/n3922 ),
    .b(1'b1),
    .c(\u2_Display/add121/c3 ),
    .o({\u2_Display/add121/c4 ,\u2_Display/n3928 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u30  (
    .a(\u2_Display/n3895 ),
    .b(1'b1),
    .c(\u2_Display/add121/c30 ),
    .o({\u2_Display/add121/c31 ,\u2_Display/n3928 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u31  (
    .a(\u2_Display/n3894 ),
    .b(1'b1),
    .c(\u2_Display/add121/c31 ),
    .o({open_n923,\u2_Display/n3928 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u4  (
    .a(\u2_Display/n3921 ),
    .b(1'b1),
    .c(\u2_Display/add121/c4 ),
    .o({\u2_Display/add121/c5 ,\u2_Display/n3928 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u5  (
    .a(\u2_Display/n3920 ),
    .b(1'b1),
    .c(\u2_Display/add121/c5 ),
    .o({\u2_Display/add121/c6 ,\u2_Display/n3928 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u6  (
    .a(\u2_Display/n3919 ),
    .b(1'b1),
    .c(\u2_Display/add121/c6 ),
    .o({\u2_Display/add121/c7 ,\u2_Display/n3928 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u7  (
    .a(\u2_Display/n3918 ),
    .b(1'b1),
    .c(\u2_Display/add121/c7 ),
    .o({\u2_Display/add121/c8 ,\u2_Display/n3928 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u8  (
    .a(\u2_Display/n3917 ),
    .b(1'b1),
    .c(\u2_Display/add121/c8 ),
    .o({\u2_Display/add121/c9 ,\u2_Display/n3928 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add121/u9  (
    .a(\u2_Display/n3916 ),
    .b(1'b1),
    .c(\u2_Display/add121/c9 ),
    .o({\u2_Display/add121/c10 ,\u2_Display/n3928 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add121/ucin  (
    .a(1'b1),
    .o({\u2_Display/add121/c0 ,open_n926}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u0  (
    .a(\u2_Display/n3960 ),
    .b(1'b1),
    .c(\u2_Display/add122/c0 ),
    .o({\u2_Display/add122/c1 ,\u2_Display/n3963 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u1  (
    .a(\u2_Display/n3959 ),
    .b(1'b1),
    .c(\u2_Display/add122/c1 ),
    .o({\u2_Display/add122/c2 ,\u2_Display/n3963 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u10  (
    .a(\u2_Display/n3950 ),
    .b(1'b1),
    .c(\u2_Display/add122/c10 ),
    .o({\u2_Display/add122/c11 ,\u2_Display/n3963 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u11  (
    .a(\u2_Display/n3949 ),
    .b(1'b1),
    .c(\u2_Display/add122/c11 ),
    .o({\u2_Display/add122/c12 ,\u2_Display/n3963 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u12  (
    .a(\u2_Display/n3948 ),
    .b(1'b1),
    .c(\u2_Display/add122/c12 ),
    .o({\u2_Display/add122/c13 ,\u2_Display/n3963 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u13  (
    .a(\u2_Display/n3947 ),
    .b(1'b1),
    .c(\u2_Display/add122/c13 ),
    .o({\u2_Display/add122/c14 ,\u2_Display/n3963 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u14  (
    .a(\u2_Display/n3946 ),
    .b(1'b1),
    .c(\u2_Display/add122/c14 ),
    .o({\u2_Display/add122/c15 ,\u2_Display/n3963 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u15  (
    .a(\u2_Display/n3945 ),
    .b(1'b1),
    .c(\u2_Display/add122/c15 ),
    .o({\u2_Display/add122/c16 ,\u2_Display/n3963 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u16  (
    .a(\u2_Display/n3944 ),
    .b(1'b1),
    .c(\u2_Display/add122/c16 ),
    .o({\u2_Display/add122/c17 ,\u2_Display/n3963 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u17  (
    .a(\u2_Display/n3943 ),
    .b(1'b1),
    .c(\u2_Display/add122/c17 ),
    .o({\u2_Display/add122/c18 ,\u2_Display/n3963 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u18  (
    .a(\u2_Display/n3942 ),
    .b(1'b1),
    .c(\u2_Display/add122/c18 ),
    .o({\u2_Display/add122/c19 ,\u2_Display/n3963 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u19  (
    .a(\u2_Display/n3941 ),
    .b(1'b1),
    .c(\u2_Display/add122/c19 ),
    .o({\u2_Display/add122/c20 ,\u2_Display/n3963 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u2  (
    .a(\u2_Display/n3958 ),
    .b(1'b1),
    .c(\u2_Display/add122/c2 ),
    .o({\u2_Display/add122/c3 ,\u2_Display/n3963 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u20  (
    .a(\u2_Display/n3940 ),
    .b(1'b1),
    .c(\u2_Display/add122/c20 ),
    .o({\u2_Display/add122/c21 ,\u2_Display/n3963 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u21  (
    .a(\u2_Display/n3939 ),
    .b(1'b1),
    .c(\u2_Display/add122/c21 ),
    .o({\u2_Display/add122/c22 ,\u2_Display/n3963 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u22  (
    .a(\u2_Display/n3938 ),
    .b(1'b0),
    .c(\u2_Display/add122/c22 ),
    .o({\u2_Display/add122/c23 ,\u2_Display/n3963 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u23  (
    .a(\u2_Display/n3937 ),
    .b(1'b1),
    .c(\u2_Display/add122/c23 ),
    .o({\u2_Display/add122/c24 ,\u2_Display/n3963 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u24  (
    .a(\u2_Display/n3936 ),
    .b(1'b1),
    .c(\u2_Display/add122/c24 ),
    .o({\u2_Display/add122/c25 ,\u2_Display/n3963 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u25  (
    .a(\u2_Display/n3935 ),
    .b(1'b0),
    .c(\u2_Display/add122/c25 ),
    .o({\u2_Display/add122/c26 ,\u2_Display/n3963 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u26  (
    .a(\u2_Display/n3934 ),
    .b(1'b0),
    .c(\u2_Display/add122/c26 ),
    .o({\u2_Display/add122/c27 ,\u2_Display/n3963 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u27  (
    .a(\u2_Display/n3933 ),
    .b(1'b1),
    .c(\u2_Display/add122/c27 ),
    .o({\u2_Display/add122/c28 ,\u2_Display/n3963 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u28  (
    .a(\u2_Display/n3932 ),
    .b(1'b1),
    .c(\u2_Display/add122/c28 ),
    .o({\u2_Display/add122/c29 ,\u2_Display/n3963 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u29  (
    .a(\u2_Display/n3931 ),
    .b(1'b1),
    .c(\u2_Display/add122/c29 ),
    .o({\u2_Display/add122/c30 ,\u2_Display/n3963 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u3  (
    .a(\u2_Display/n3957 ),
    .b(1'b1),
    .c(\u2_Display/add122/c3 ),
    .o({\u2_Display/add122/c4 ,\u2_Display/n3963 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u30  (
    .a(\u2_Display/n3930 ),
    .b(1'b1),
    .c(\u2_Display/add122/c30 ),
    .o({\u2_Display/add122/c31 ,\u2_Display/n3963 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u31  (
    .a(\u2_Display/n3929 ),
    .b(1'b1),
    .c(\u2_Display/add122/c31 ),
    .o({open_n927,\u2_Display/n3963 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u4  (
    .a(\u2_Display/n3956 ),
    .b(1'b1),
    .c(\u2_Display/add122/c4 ),
    .o({\u2_Display/add122/c5 ,\u2_Display/n3963 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u5  (
    .a(\u2_Display/n3955 ),
    .b(1'b1),
    .c(\u2_Display/add122/c5 ),
    .o({\u2_Display/add122/c6 ,\u2_Display/n3963 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u6  (
    .a(\u2_Display/n3954 ),
    .b(1'b1),
    .c(\u2_Display/add122/c6 ),
    .o({\u2_Display/add122/c7 ,\u2_Display/n3963 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u7  (
    .a(\u2_Display/n3953 ),
    .b(1'b1),
    .c(\u2_Display/add122/c7 ),
    .o({\u2_Display/add122/c8 ,\u2_Display/n3963 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u8  (
    .a(\u2_Display/n3952 ),
    .b(1'b1),
    .c(\u2_Display/add122/c8 ),
    .o({\u2_Display/add122/c9 ,\u2_Display/n3963 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add122/u9  (
    .a(\u2_Display/n3951 ),
    .b(1'b1),
    .c(\u2_Display/add122/c9 ),
    .o({\u2_Display/add122/c10 ,\u2_Display/n3963 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add122/ucin  (
    .a(1'b1),
    .o({\u2_Display/add122/c0 ,open_n930}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u0  (
    .a(\u2_Display/n3995 ),
    .b(1'b1),
    .c(\u2_Display/add123/c0 ),
    .o({\u2_Display/add123/c1 ,\u2_Display/n3998 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u1  (
    .a(\u2_Display/n3994 ),
    .b(1'b1),
    .c(\u2_Display/add123/c1 ),
    .o({\u2_Display/add123/c2 ,\u2_Display/n3998 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u10  (
    .a(\u2_Display/n3985 ),
    .b(1'b1),
    .c(\u2_Display/add123/c10 ),
    .o({\u2_Display/add123/c11 ,\u2_Display/n3998 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u11  (
    .a(\u2_Display/n3984 ),
    .b(1'b1),
    .c(\u2_Display/add123/c11 ),
    .o({\u2_Display/add123/c12 ,\u2_Display/n3998 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u12  (
    .a(\u2_Display/n3983 ),
    .b(1'b1),
    .c(\u2_Display/add123/c12 ),
    .o({\u2_Display/add123/c13 ,\u2_Display/n3998 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u13  (
    .a(\u2_Display/n3982 ),
    .b(1'b1),
    .c(\u2_Display/add123/c13 ),
    .o({\u2_Display/add123/c14 ,\u2_Display/n3998 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u14  (
    .a(\u2_Display/n3981 ),
    .b(1'b1),
    .c(\u2_Display/add123/c14 ),
    .o({\u2_Display/add123/c15 ,\u2_Display/n3998 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u15  (
    .a(\u2_Display/n3980 ),
    .b(1'b1),
    .c(\u2_Display/add123/c15 ),
    .o({\u2_Display/add123/c16 ,\u2_Display/n3998 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u16  (
    .a(\u2_Display/n3979 ),
    .b(1'b1),
    .c(\u2_Display/add123/c16 ),
    .o({\u2_Display/add123/c17 ,\u2_Display/n3998 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u17  (
    .a(\u2_Display/n3978 ),
    .b(1'b1),
    .c(\u2_Display/add123/c17 ),
    .o({\u2_Display/add123/c18 ,\u2_Display/n3998 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u18  (
    .a(\u2_Display/n3977 ),
    .b(1'b1),
    .c(\u2_Display/add123/c18 ),
    .o({\u2_Display/add123/c19 ,\u2_Display/n3998 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u19  (
    .a(\u2_Display/n3976 ),
    .b(1'b1),
    .c(\u2_Display/add123/c19 ),
    .o({\u2_Display/add123/c20 ,\u2_Display/n3998 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u2  (
    .a(\u2_Display/n3993 ),
    .b(1'b1),
    .c(\u2_Display/add123/c2 ),
    .o({\u2_Display/add123/c3 ,\u2_Display/n3998 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u20  (
    .a(\u2_Display/n3975 ),
    .b(1'b1),
    .c(\u2_Display/add123/c20 ),
    .o({\u2_Display/add123/c21 ,\u2_Display/n3998 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u21  (
    .a(\u2_Display/n3974 ),
    .b(1'b0),
    .c(\u2_Display/add123/c21 ),
    .o({\u2_Display/add123/c22 ,\u2_Display/n3998 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u22  (
    .a(\u2_Display/n3973 ),
    .b(1'b1),
    .c(\u2_Display/add123/c22 ),
    .o({\u2_Display/add123/c23 ,\u2_Display/n3998 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u23  (
    .a(\u2_Display/n3972 ),
    .b(1'b1),
    .c(\u2_Display/add123/c23 ),
    .o({\u2_Display/add123/c24 ,\u2_Display/n3998 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u24  (
    .a(\u2_Display/n3971 ),
    .b(1'b0),
    .c(\u2_Display/add123/c24 ),
    .o({\u2_Display/add123/c25 ,\u2_Display/n3998 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u25  (
    .a(\u2_Display/n3970 ),
    .b(1'b0),
    .c(\u2_Display/add123/c25 ),
    .o({\u2_Display/add123/c26 ,\u2_Display/n3998 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u26  (
    .a(\u2_Display/n3969 ),
    .b(1'b1),
    .c(\u2_Display/add123/c26 ),
    .o({\u2_Display/add123/c27 ,\u2_Display/n3998 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u27  (
    .a(\u2_Display/n3968 ),
    .b(1'b1),
    .c(\u2_Display/add123/c27 ),
    .o({\u2_Display/add123/c28 ,\u2_Display/n3998 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u28  (
    .a(\u2_Display/n3967 ),
    .b(1'b1),
    .c(\u2_Display/add123/c28 ),
    .o({\u2_Display/add123/c29 ,\u2_Display/n3998 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u29  (
    .a(\u2_Display/n3966 ),
    .b(1'b1),
    .c(\u2_Display/add123/c29 ),
    .o({\u2_Display/add123/c30 ,\u2_Display/n3998 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u3  (
    .a(\u2_Display/n3992 ),
    .b(1'b1),
    .c(\u2_Display/add123/c3 ),
    .o({\u2_Display/add123/c4 ,\u2_Display/n3998 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u30  (
    .a(\u2_Display/n3965 ),
    .b(1'b1),
    .c(\u2_Display/add123/c30 ),
    .o({\u2_Display/add123/c31 ,\u2_Display/n3998 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u31  (
    .a(\u2_Display/n3964 ),
    .b(1'b1),
    .c(\u2_Display/add123/c31 ),
    .o({open_n931,\u2_Display/n3998 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u4  (
    .a(\u2_Display/n3991 ),
    .b(1'b1),
    .c(\u2_Display/add123/c4 ),
    .o({\u2_Display/add123/c5 ,\u2_Display/n3998 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u5  (
    .a(\u2_Display/n3990 ),
    .b(1'b1),
    .c(\u2_Display/add123/c5 ),
    .o({\u2_Display/add123/c6 ,\u2_Display/n3998 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u6  (
    .a(\u2_Display/n3989 ),
    .b(1'b1),
    .c(\u2_Display/add123/c6 ),
    .o({\u2_Display/add123/c7 ,\u2_Display/n3998 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u7  (
    .a(\u2_Display/n3988 ),
    .b(1'b1),
    .c(\u2_Display/add123/c7 ),
    .o({\u2_Display/add123/c8 ,\u2_Display/n3998 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u8  (
    .a(\u2_Display/n3987 ),
    .b(1'b1),
    .c(\u2_Display/add123/c8 ),
    .o({\u2_Display/add123/c9 ,\u2_Display/n3998 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add123/u9  (
    .a(\u2_Display/n3986 ),
    .b(1'b1),
    .c(\u2_Display/add123/c9 ),
    .o({\u2_Display/add123/c10 ,\u2_Display/n3998 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add123/ucin  (
    .a(1'b1),
    .o({\u2_Display/add123/c0 ,open_n934}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u0  (
    .a(\u2_Display/n4030 ),
    .b(1'b1),
    .c(\u2_Display/add124/c0 ),
    .o({\u2_Display/add124/c1 ,\u2_Display/n4033 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u1  (
    .a(\u2_Display/n4029 ),
    .b(1'b1),
    .c(\u2_Display/add124/c1 ),
    .o({\u2_Display/add124/c2 ,\u2_Display/n4033 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u10  (
    .a(\u2_Display/n4020 ),
    .b(1'b1),
    .c(\u2_Display/add124/c10 ),
    .o({\u2_Display/add124/c11 ,\u2_Display/n4033 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u11  (
    .a(\u2_Display/n4019 ),
    .b(1'b1),
    .c(\u2_Display/add124/c11 ),
    .o({\u2_Display/add124/c12 ,\u2_Display/n4033 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u12  (
    .a(\u2_Display/n4018 ),
    .b(1'b1),
    .c(\u2_Display/add124/c12 ),
    .o({\u2_Display/add124/c13 ,\u2_Display/n4033 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u13  (
    .a(\u2_Display/n4017 ),
    .b(1'b1),
    .c(\u2_Display/add124/c13 ),
    .o({\u2_Display/add124/c14 ,\u2_Display/n4033 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u14  (
    .a(\u2_Display/n4016 ),
    .b(1'b1),
    .c(\u2_Display/add124/c14 ),
    .o({\u2_Display/add124/c15 ,\u2_Display/n4033 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u15  (
    .a(\u2_Display/n4015 ),
    .b(1'b1),
    .c(\u2_Display/add124/c15 ),
    .o({\u2_Display/add124/c16 ,\u2_Display/n4033 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u16  (
    .a(\u2_Display/n4014 ),
    .b(1'b1),
    .c(\u2_Display/add124/c16 ),
    .o({\u2_Display/add124/c17 ,\u2_Display/n4033 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u17  (
    .a(\u2_Display/n4013 ),
    .b(1'b1),
    .c(\u2_Display/add124/c17 ),
    .o({\u2_Display/add124/c18 ,\u2_Display/n4033 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u18  (
    .a(\u2_Display/n4012 ),
    .b(1'b1),
    .c(\u2_Display/add124/c18 ),
    .o({\u2_Display/add124/c19 ,\u2_Display/n4033 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u19  (
    .a(\u2_Display/n4011 ),
    .b(1'b1),
    .c(\u2_Display/add124/c19 ),
    .o({\u2_Display/add124/c20 ,\u2_Display/n4033 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u2  (
    .a(\u2_Display/n4028 ),
    .b(1'b1),
    .c(\u2_Display/add124/c2 ),
    .o({\u2_Display/add124/c3 ,\u2_Display/n4033 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u20  (
    .a(\u2_Display/n4010 ),
    .b(1'b0),
    .c(\u2_Display/add124/c20 ),
    .o({\u2_Display/add124/c21 ,\u2_Display/n4033 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u21  (
    .a(\u2_Display/n4009 ),
    .b(1'b1),
    .c(\u2_Display/add124/c21 ),
    .o({\u2_Display/add124/c22 ,\u2_Display/n4033 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u22  (
    .a(\u2_Display/n4008 ),
    .b(1'b1),
    .c(\u2_Display/add124/c22 ),
    .o({\u2_Display/add124/c23 ,\u2_Display/n4033 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u23  (
    .a(\u2_Display/n4007 ),
    .b(1'b0),
    .c(\u2_Display/add124/c23 ),
    .o({\u2_Display/add124/c24 ,\u2_Display/n4033 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u24  (
    .a(\u2_Display/n4006 ),
    .b(1'b0),
    .c(\u2_Display/add124/c24 ),
    .o({\u2_Display/add124/c25 ,\u2_Display/n4033 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u25  (
    .a(\u2_Display/n4005 ),
    .b(1'b1),
    .c(\u2_Display/add124/c25 ),
    .o({\u2_Display/add124/c26 ,\u2_Display/n4033 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u26  (
    .a(\u2_Display/n4004 ),
    .b(1'b1),
    .c(\u2_Display/add124/c26 ),
    .o({\u2_Display/add124/c27 ,\u2_Display/n4033 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u27  (
    .a(\u2_Display/n4003 ),
    .b(1'b1),
    .c(\u2_Display/add124/c27 ),
    .o({\u2_Display/add124/c28 ,\u2_Display/n4033 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u28  (
    .a(\u2_Display/n4002 ),
    .b(1'b1),
    .c(\u2_Display/add124/c28 ),
    .o({\u2_Display/add124/c29 ,\u2_Display/n4033 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u29  (
    .a(\u2_Display/n4001 ),
    .b(1'b1),
    .c(\u2_Display/add124/c29 ),
    .o({\u2_Display/add124/c30 ,\u2_Display/n4033 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u3  (
    .a(\u2_Display/n4027 ),
    .b(1'b1),
    .c(\u2_Display/add124/c3 ),
    .o({\u2_Display/add124/c4 ,\u2_Display/n4033 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u30  (
    .a(\u2_Display/n4000 ),
    .b(1'b1),
    .c(\u2_Display/add124/c30 ),
    .o({\u2_Display/add124/c31 ,\u2_Display/n4033 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u31  (
    .a(\u2_Display/n3999 ),
    .b(1'b1),
    .c(\u2_Display/add124/c31 ),
    .o({open_n935,\u2_Display/n4033 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u4  (
    .a(\u2_Display/n4026 ),
    .b(1'b1),
    .c(\u2_Display/add124/c4 ),
    .o({\u2_Display/add124/c5 ,\u2_Display/n4033 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u5  (
    .a(\u2_Display/n4025 ),
    .b(1'b1),
    .c(\u2_Display/add124/c5 ),
    .o({\u2_Display/add124/c6 ,\u2_Display/n4033 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u6  (
    .a(\u2_Display/n4024 ),
    .b(1'b1),
    .c(\u2_Display/add124/c6 ),
    .o({\u2_Display/add124/c7 ,\u2_Display/n4033 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u7  (
    .a(\u2_Display/n4023 ),
    .b(1'b1),
    .c(\u2_Display/add124/c7 ),
    .o({\u2_Display/add124/c8 ,\u2_Display/n4033 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u8  (
    .a(\u2_Display/n4022 ),
    .b(1'b1),
    .c(\u2_Display/add124/c8 ),
    .o({\u2_Display/add124/c9 ,\u2_Display/n4033 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add124/u9  (
    .a(\u2_Display/n4021 ),
    .b(1'b1),
    .c(\u2_Display/add124/c9 ),
    .o({\u2_Display/add124/c10 ,\u2_Display/n4033 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add124/ucin  (
    .a(1'b1),
    .o({\u2_Display/add124/c0 ,open_n938}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u0  (
    .a(\u2_Display/n4065 ),
    .b(1'b1),
    .c(\u2_Display/add125/c0 ),
    .o({\u2_Display/add125/c1 ,\u2_Display/n4068 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u1  (
    .a(\u2_Display/n4064 ),
    .b(1'b1),
    .c(\u2_Display/add125/c1 ),
    .o({\u2_Display/add125/c2 ,\u2_Display/n4068 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u10  (
    .a(\u2_Display/n4055 ),
    .b(1'b1),
    .c(\u2_Display/add125/c10 ),
    .o({\u2_Display/add125/c11 ,\u2_Display/n4068 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u11  (
    .a(\u2_Display/n4054 ),
    .b(1'b1),
    .c(\u2_Display/add125/c11 ),
    .o({\u2_Display/add125/c12 ,\u2_Display/n4068 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u12  (
    .a(\u2_Display/n4053 ),
    .b(1'b1),
    .c(\u2_Display/add125/c12 ),
    .o({\u2_Display/add125/c13 ,\u2_Display/n4068 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u13  (
    .a(\u2_Display/n4052 ),
    .b(1'b1),
    .c(\u2_Display/add125/c13 ),
    .o({\u2_Display/add125/c14 ,\u2_Display/n4068 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u14  (
    .a(\u2_Display/n4051 ),
    .b(1'b1),
    .c(\u2_Display/add125/c14 ),
    .o({\u2_Display/add125/c15 ,\u2_Display/n4068 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u15  (
    .a(\u2_Display/n4050 ),
    .b(1'b1),
    .c(\u2_Display/add125/c15 ),
    .o({\u2_Display/add125/c16 ,\u2_Display/n4068 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u16  (
    .a(\u2_Display/n4049 ),
    .b(1'b1),
    .c(\u2_Display/add125/c16 ),
    .o({\u2_Display/add125/c17 ,\u2_Display/n4068 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u17  (
    .a(\u2_Display/n4048 ),
    .b(1'b1),
    .c(\u2_Display/add125/c17 ),
    .o({\u2_Display/add125/c18 ,\u2_Display/n4068 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u18  (
    .a(\u2_Display/n4047 ),
    .b(1'b1),
    .c(\u2_Display/add125/c18 ),
    .o({\u2_Display/add125/c19 ,\u2_Display/n4068 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u19  (
    .a(\u2_Display/n4046 ),
    .b(1'b0),
    .c(\u2_Display/add125/c19 ),
    .o({\u2_Display/add125/c20 ,\u2_Display/n4068 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u2  (
    .a(\u2_Display/n4063 ),
    .b(1'b1),
    .c(\u2_Display/add125/c2 ),
    .o({\u2_Display/add125/c3 ,\u2_Display/n4068 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u20  (
    .a(\u2_Display/n4045 ),
    .b(1'b1),
    .c(\u2_Display/add125/c20 ),
    .o({\u2_Display/add125/c21 ,\u2_Display/n4068 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u21  (
    .a(\u2_Display/n4044 ),
    .b(1'b1),
    .c(\u2_Display/add125/c21 ),
    .o({\u2_Display/add125/c22 ,\u2_Display/n4068 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u22  (
    .a(\u2_Display/n4043 ),
    .b(1'b0),
    .c(\u2_Display/add125/c22 ),
    .o({\u2_Display/add125/c23 ,\u2_Display/n4068 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u23  (
    .a(\u2_Display/n4042 ),
    .b(1'b0),
    .c(\u2_Display/add125/c23 ),
    .o({\u2_Display/add125/c24 ,\u2_Display/n4068 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u24  (
    .a(\u2_Display/n4041 ),
    .b(1'b1),
    .c(\u2_Display/add125/c24 ),
    .o({\u2_Display/add125/c25 ,\u2_Display/n4068 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u25  (
    .a(\u2_Display/n4040 ),
    .b(1'b1),
    .c(\u2_Display/add125/c25 ),
    .o({\u2_Display/add125/c26 ,\u2_Display/n4068 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u26  (
    .a(\u2_Display/n4039 ),
    .b(1'b1),
    .c(\u2_Display/add125/c26 ),
    .o({\u2_Display/add125/c27 ,\u2_Display/n4068 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u27  (
    .a(\u2_Display/n4038 ),
    .b(1'b1),
    .c(\u2_Display/add125/c27 ),
    .o({\u2_Display/add125/c28 ,\u2_Display/n4068 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u28  (
    .a(\u2_Display/n4037 ),
    .b(1'b1),
    .c(\u2_Display/add125/c28 ),
    .o({\u2_Display/add125/c29 ,\u2_Display/n4068 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u29  (
    .a(\u2_Display/n4036 ),
    .b(1'b1),
    .c(\u2_Display/add125/c29 ),
    .o({\u2_Display/add125/c30 ,\u2_Display/n4068 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u3  (
    .a(\u2_Display/n4062 ),
    .b(1'b1),
    .c(\u2_Display/add125/c3 ),
    .o({\u2_Display/add125/c4 ,\u2_Display/n4068 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u30  (
    .a(\u2_Display/n4035 ),
    .b(1'b1),
    .c(\u2_Display/add125/c30 ),
    .o({\u2_Display/add125/c31 ,\u2_Display/n4068 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u31  (
    .a(\u2_Display/n4034 ),
    .b(1'b1),
    .c(\u2_Display/add125/c31 ),
    .o({open_n939,\u2_Display/n4068 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u4  (
    .a(\u2_Display/n4061 ),
    .b(1'b1),
    .c(\u2_Display/add125/c4 ),
    .o({\u2_Display/add125/c5 ,\u2_Display/n4068 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u5  (
    .a(\u2_Display/n4060 ),
    .b(1'b1),
    .c(\u2_Display/add125/c5 ),
    .o({\u2_Display/add125/c6 ,\u2_Display/n4068 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u6  (
    .a(\u2_Display/n4059 ),
    .b(1'b1),
    .c(\u2_Display/add125/c6 ),
    .o({\u2_Display/add125/c7 ,\u2_Display/n4068 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u7  (
    .a(\u2_Display/n4058 ),
    .b(1'b1),
    .c(\u2_Display/add125/c7 ),
    .o({\u2_Display/add125/c8 ,\u2_Display/n4068 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u8  (
    .a(\u2_Display/n4057 ),
    .b(1'b1),
    .c(\u2_Display/add125/c8 ),
    .o({\u2_Display/add125/c9 ,\u2_Display/n4068 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add125/u9  (
    .a(\u2_Display/n4056 ),
    .b(1'b1),
    .c(\u2_Display/add125/c9 ),
    .o({\u2_Display/add125/c10 ,\u2_Display/n4068 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add125/ucin  (
    .a(1'b1),
    .o({\u2_Display/add125/c0 ,open_n942}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u0  (
    .a(\u2_Display/n4100 ),
    .b(1'b1),
    .c(\u2_Display/add126/c0 ),
    .o({\u2_Display/add126/c1 ,\u2_Display/n4103 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u1  (
    .a(\u2_Display/n4099 ),
    .b(1'b1),
    .c(\u2_Display/add126/c1 ),
    .o({\u2_Display/add126/c2 ,\u2_Display/n4103 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u10  (
    .a(\u2_Display/n4090 ),
    .b(1'b1),
    .c(\u2_Display/add126/c10 ),
    .o({\u2_Display/add126/c11 ,\u2_Display/n4103 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u11  (
    .a(\u2_Display/n4089 ),
    .b(1'b1),
    .c(\u2_Display/add126/c11 ),
    .o({\u2_Display/add126/c12 ,\u2_Display/n4103 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u12  (
    .a(\u2_Display/n4088 ),
    .b(1'b1),
    .c(\u2_Display/add126/c12 ),
    .o({\u2_Display/add126/c13 ,\u2_Display/n4103 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u13  (
    .a(\u2_Display/n4087 ),
    .b(1'b1),
    .c(\u2_Display/add126/c13 ),
    .o({\u2_Display/add126/c14 ,\u2_Display/n4103 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u14  (
    .a(\u2_Display/n4086 ),
    .b(1'b1),
    .c(\u2_Display/add126/c14 ),
    .o({\u2_Display/add126/c15 ,\u2_Display/n4103 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u15  (
    .a(\u2_Display/n4085 ),
    .b(1'b1),
    .c(\u2_Display/add126/c15 ),
    .o({\u2_Display/add126/c16 ,\u2_Display/n4103 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u16  (
    .a(\u2_Display/n4084 ),
    .b(1'b1),
    .c(\u2_Display/add126/c16 ),
    .o({\u2_Display/add126/c17 ,\u2_Display/n4103 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u17  (
    .a(\u2_Display/n4083 ),
    .b(1'b1),
    .c(\u2_Display/add126/c17 ),
    .o({\u2_Display/add126/c18 ,\u2_Display/n4103 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u18  (
    .a(\u2_Display/n4082 ),
    .b(1'b0),
    .c(\u2_Display/add126/c18 ),
    .o({\u2_Display/add126/c19 ,\u2_Display/n4103 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u19  (
    .a(\u2_Display/n4081 ),
    .b(1'b1),
    .c(\u2_Display/add126/c19 ),
    .o({\u2_Display/add126/c20 ,\u2_Display/n4103 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u2  (
    .a(\u2_Display/n4098 ),
    .b(1'b1),
    .c(\u2_Display/add126/c2 ),
    .o({\u2_Display/add126/c3 ,\u2_Display/n4103 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u20  (
    .a(\u2_Display/n4080 ),
    .b(1'b1),
    .c(\u2_Display/add126/c20 ),
    .o({\u2_Display/add126/c21 ,\u2_Display/n4103 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u21  (
    .a(\u2_Display/n4079 ),
    .b(1'b0),
    .c(\u2_Display/add126/c21 ),
    .o({\u2_Display/add126/c22 ,\u2_Display/n4103 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u22  (
    .a(\u2_Display/n4078 ),
    .b(1'b0),
    .c(\u2_Display/add126/c22 ),
    .o({\u2_Display/add126/c23 ,\u2_Display/n4103 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u23  (
    .a(\u2_Display/n4077 ),
    .b(1'b1),
    .c(\u2_Display/add126/c23 ),
    .o({\u2_Display/add126/c24 ,\u2_Display/n4103 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u24  (
    .a(\u2_Display/n4076 ),
    .b(1'b1),
    .c(\u2_Display/add126/c24 ),
    .o({\u2_Display/add126/c25 ,\u2_Display/n4103 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u25  (
    .a(\u2_Display/n4075 ),
    .b(1'b1),
    .c(\u2_Display/add126/c25 ),
    .o({\u2_Display/add126/c26 ,\u2_Display/n4103 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u26  (
    .a(\u2_Display/n4074 ),
    .b(1'b1),
    .c(\u2_Display/add126/c26 ),
    .o({\u2_Display/add126/c27 ,\u2_Display/n4103 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u27  (
    .a(\u2_Display/n4073 ),
    .b(1'b1),
    .c(\u2_Display/add126/c27 ),
    .o({\u2_Display/add126/c28 ,\u2_Display/n4103 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u28  (
    .a(\u2_Display/n4072 ),
    .b(1'b1),
    .c(\u2_Display/add126/c28 ),
    .o({\u2_Display/add126/c29 ,\u2_Display/n4103 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u29  (
    .a(\u2_Display/n4071 ),
    .b(1'b1),
    .c(\u2_Display/add126/c29 ),
    .o({\u2_Display/add126/c30 ,\u2_Display/n4103 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u3  (
    .a(\u2_Display/n4097 ),
    .b(1'b1),
    .c(\u2_Display/add126/c3 ),
    .o({\u2_Display/add126/c4 ,\u2_Display/n4103 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u30  (
    .a(\u2_Display/n4070 ),
    .b(1'b1),
    .c(\u2_Display/add126/c30 ),
    .o({\u2_Display/add126/c31 ,\u2_Display/n4103 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u31  (
    .a(\u2_Display/n4069 ),
    .b(1'b1),
    .c(\u2_Display/add126/c31 ),
    .o({open_n943,\u2_Display/n4103 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u4  (
    .a(\u2_Display/n4096 ),
    .b(1'b1),
    .c(\u2_Display/add126/c4 ),
    .o({\u2_Display/add126/c5 ,\u2_Display/n4103 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u5  (
    .a(\u2_Display/n4095 ),
    .b(1'b1),
    .c(\u2_Display/add126/c5 ),
    .o({\u2_Display/add126/c6 ,\u2_Display/n4103 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u6  (
    .a(\u2_Display/n4094 ),
    .b(1'b1),
    .c(\u2_Display/add126/c6 ),
    .o({\u2_Display/add126/c7 ,\u2_Display/n4103 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u7  (
    .a(\u2_Display/n4093 ),
    .b(1'b1),
    .c(\u2_Display/add126/c7 ),
    .o({\u2_Display/add126/c8 ,\u2_Display/n4103 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u8  (
    .a(\u2_Display/n4092 ),
    .b(1'b1),
    .c(\u2_Display/add126/c8 ),
    .o({\u2_Display/add126/c9 ,\u2_Display/n4103 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add126/u9  (
    .a(\u2_Display/n4091 ),
    .b(1'b1),
    .c(\u2_Display/add126/c9 ),
    .o({\u2_Display/add126/c10 ,\u2_Display/n4103 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add126/ucin  (
    .a(1'b1),
    .o({\u2_Display/add126/c0 ,open_n946}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u0  (
    .a(\u2_Display/n4135 ),
    .b(1'b1),
    .c(\u2_Display/add127/c0 ),
    .o({\u2_Display/add127/c1 ,\u2_Display/n4138 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u1  (
    .a(\u2_Display/n4134 ),
    .b(1'b1),
    .c(\u2_Display/add127/c1 ),
    .o({\u2_Display/add127/c2 ,\u2_Display/n4138 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u10  (
    .a(\u2_Display/n4125 ),
    .b(1'b1),
    .c(\u2_Display/add127/c10 ),
    .o({\u2_Display/add127/c11 ,\u2_Display/n4138 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u11  (
    .a(\u2_Display/n4124 ),
    .b(1'b1),
    .c(\u2_Display/add127/c11 ),
    .o({\u2_Display/add127/c12 ,\u2_Display/n4138 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u12  (
    .a(\u2_Display/n4123 ),
    .b(1'b1),
    .c(\u2_Display/add127/c12 ),
    .o({\u2_Display/add127/c13 ,\u2_Display/n4138 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u13  (
    .a(\u2_Display/n4122 ),
    .b(1'b1),
    .c(\u2_Display/add127/c13 ),
    .o({\u2_Display/add127/c14 ,\u2_Display/n4138 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u14  (
    .a(\u2_Display/n4121 ),
    .b(1'b1),
    .c(\u2_Display/add127/c14 ),
    .o({\u2_Display/add127/c15 ,\u2_Display/n4138 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u15  (
    .a(\u2_Display/n4120 ),
    .b(1'b1),
    .c(\u2_Display/add127/c15 ),
    .o({\u2_Display/add127/c16 ,\u2_Display/n4138 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u16  (
    .a(\u2_Display/n4119 ),
    .b(1'b1),
    .c(\u2_Display/add127/c16 ),
    .o({\u2_Display/add127/c17 ,\u2_Display/n4138 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u17  (
    .a(\u2_Display/n4118 ),
    .b(1'b0),
    .c(\u2_Display/add127/c17 ),
    .o({\u2_Display/add127/c18 ,\u2_Display/n4138 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u18  (
    .a(\u2_Display/n4117 ),
    .b(1'b1),
    .c(\u2_Display/add127/c18 ),
    .o({\u2_Display/add127/c19 ,\u2_Display/n4138 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u19  (
    .a(\u2_Display/n4116 ),
    .b(1'b1),
    .c(\u2_Display/add127/c19 ),
    .o({\u2_Display/add127/c20 ,\u2_Display/n4138 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u2  (
    .a(\u2_Display/n4133 ),
    .b(1'b1),
    .c(\u2_Display/add127/c2 ),
    .o({\u2_Display/add127/c3 ,\u2_Display/n4138 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u20  (
    .a(\u2_Display/n4115 ),
    .b(1'b0),
    .c(\u2_Display/add127/c20 ),
    .o({\u2_Display/add127/c21 ,\u2_Display/n4138 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u21  (
    .a(\u2_Display/n4114 ),
    .b(1'b0),
    .c(\u2_Display/add127/c21 ),
    .o({\u2_Display/add127/c22 ,\u2_Display/n4138 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u22  (
    .a(\u2_Display/n4113 ),
    .b(1'b1),
    .c(\u2_Display/add127/c22 ),
    .o({\u2_Display/add127/c23 ,\u2_Display/n4138 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u23  (
    .a(\u2_Display/n4112 ),
    .b(1'b1),
    .c(\u2_Display/add127/c23 ),
    .o({\u2_Display/add127/c24 ,\u2_Display/n4138 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u24  (
    .a(\u2_Display/n4111 ),
    .b(1'b1),
    .c(\u2_Display/add127/c24 ),
    .o({\u2_Display/add127/c25 ,\u2_Display/n4138 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u25  (
    .a(\u2_Display/n4110 ),
    .b(1'b1),
    .c(\u2_Display/add127/c25 ),
    .o({\u2_Display/add127/c26 ,\u2_Display/n4138 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u26  (
    .a(\u2_Display/n4109 ),
    .b(1'b1),
    .c(\u2_Display/add127/c26 ),
    .o({\u2_Display/add127/c27 ,\u2_Display/n4138 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u27  (
    .a(\u2_Display/n4108 ),
    .b(1'b1),
    .c(\u2_Display/add127/c27 ),
    .o({\u2_Display/add127/c28 ,\u2_Display/n4138 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u28  (
    .a(\u2_Display/n4107 ),
    .b(1'b1),
    .c(\u2_Display/add127/c28 ),
    .o({\u2_Display/add127/c29 ,\u2_Display/n4138 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u29  (
    .a(\u2_Display/n4106 ),
    .b(1'b1),
    .c(\u2_Display/add127/c29 ),
    .o({\u2_Display/add127/c30 ,\u2_Display/n4138 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u3  (
    .a(\u2_Display/n4132 ),
    .b(1'b1),
    .c(\u2_Display/add127/c3 ),
    .o({\u2_Display/add127/c4 ,\u2_Display/n4138 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u30  (
    .a(\u2_Display/n4105 ),
    .b(1'b1),
    .c(\u2_Display/add127/c30 ),
    .o({\u2_Display/add127/c31 ,\u2_Display/n4138 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u31  (
    .a(\u2_Display/n4104 ),
    .b(1'b1),
    .c(\u2_Display/add127/c31 ),
    .o({open_n947,\u2_Display/n4138 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u4  (
    .a(\u2_Display/n4131 ),
    .b(1'b1),
    .c(\u2_Display/add127/c4 ),
    .o({\u2_Display/add127/c5 ,\u2_Display/n4138 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u5  (
    .a(\u2_Display/n4130 ),
    .b(1'b1),
    .c(\u2_Display/add127/c5 ),
    .o({\u2_Display/add127/c6 ,\u2_Display/n4138 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u6  (
    .a(\u2_Display/n4129 ),
    .b(1'b1),
    .c(\u2_Display/add127/c6 ),
    .o({\u2_Display/add127/c7 ,\u2_Display/n4138 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u7  (
    .a(\u2_Display/n4128 ),
    .b(1'b1),
    .c(\u2_Display/add127/c7 ),
    .o({\u2_Display/add127/c8 ,\u2_Display/n4138 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u8  (
    .a(\u2_Display/n4127 ),
    .b(1'b1),
    .c(\u2_Display/add127/c8 ),
    .o({\u2_Display/add127/c9 ,\u2_Display/n4138 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add127/u9  (
    .a(\u2_Display/n4126 ),
    .b(1'b1),
    .c(\u2_Display/add127/c9 ),
    .o({\u2_Display/add127/c10 ,\u2_Display/n4138 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add127/ucin  (
    .a(1'b1),
    .o({\u2_Display/add127/c0 ,open_n950}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u0  (
    .a(\u2_Display/n4170 ),
    .b(1'b1),
    .c(\u2_Display/add128/c0 ),
    .o({\u2_Display/add128/c1 ,\u2_Display/n4173 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u1  (
    .a(\u2_Display/n4169 ),
    .b(1'b1),
    .c(\u2_Display/add128/c1 ),
    .o({\u2_Display/add128/c2 ,\u2_Display/n4173 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u10  (
    .a(\u2_Display/n4160 ),
    .b(1'b1),
    .c(\u2_Display/add128/c10 ),
    .o({\u2_Display/add128/c11 ,\u2_Display/n4173 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u11  (
    .a(\u2_Display/n4159 ),
    .b(1'b1),
    .c(\u2_Display/add128/c11 ),
    .o({\u2_Display/add128/c12 ,\u2_Display/n4173 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u12  (
    .a(\u2_Display/n4158 ),
    .b(1'b1),
    .c(\u2_Display/add128/c12 ),
    .o({\u2_Display/add128/c13 ,\u2_Display/n4173 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u13  (
    .a(\u2_Display/n4157 ),
    .b(1'b1),
    .c(\u2_Display/add128/c13 ),
    .o({\u2_Display/add128/c14 ,\u2_Display/n4173 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u14  (
    .a(\u2_Display/n4156 ),
    .b(1'b1),
    .c(\u2_Display/add128/c14 ),
    .o({\u2_Display/add128/c15 ,\u2_Display/n4173 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u15  (
    .a(\u2_Display/n4155 ),
    .b(1'b1),
    .c(\u2_Display/add128/c15 ),
    .o({\u2_Display/add128/c16 ,\u2_Display/n4173 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u16  (
    .a(\u2_Display/n4154 ),
    .b(1'b0),
    .c(\u2_Display/add128/c16 ),
    .o({\u2_Display/add128/c17 ,\u2_Display/n4173 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u17  (
    .a(\u2_Display/n4153 ),
    .b(1'b1),
    .c(\u2_Display/add128/c17 ),
    .o({\u2_Display/add128/c18 ,\u2_Display/n4173 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u18  (
    .a(\u2_Display/n4152 ),
    .b(1'b1),
    .c(\u2_Display/add128/c18 ),
    .o({\u2_Display/add128/c19 ,\u2_Display/n4173 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u19  (
    .a(\u2_Display/n4151 ),
    .b(1'b0),
    .c(\u2_Display/add128/c19 ),
    .o({\u2_Display/add128/c20 ,\u2_Display/n4173 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u2  (
    .a(\u2_Display/n4168 ),
    .b(1'b1),
    .c(\u2_Display/add128/c2 ),
    .o({\u2_Display/add128/c3 ,\u2_Display/n4173 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u20  (
    .a(\u2_Display/n4150 ),
    .b(1'b0),
    .c(\u2_Display/add128/c20 ),
    .o({\u2_Display/add128/c21 ,\u2_Display/n4173 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u21  (
    .a(\u2_Display/n4149 ),
    .b(1'b1),
    .c(\u2_Display/add128/c21 ),
    .o({\u2_Display/add128/c22 ,\u2_Display/n4173 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u22  (
    .a(\u2_Display/n4148 ),
    .b(1'b1),
    .c(\u2_Display/add128/c22 ),
    .o({\u2_Display/add128/c23 ,\u2_Display/n4173 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u23  (
    .a(\u2_Display/n4147 ),
    .b(1'b1),
    .c(\u2_Display/add128/c23 ),
    .o({\u2_Display/add128/c24 ,\u2_Display/n4173 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u24  (
    .a(\u2_Display/n4146 ),
    .b(1'b1),
    .c(\u2_Display/add128/c24 ),
    .o({\u2_Display/add128/c25 ,\u2_Display/n4173 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u25  (
    .a(\u2_Display/n4145 ),
    .b(1'b1),
    .c(\u2_Display/add128/c25 ),
    .o({\u2_Display/add128/c26 ,\u2_Display/n4173 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u26  (
    .a(\u2_Display/n4144 ),
    .b(1'b1),
    .c(\u2_Display/add128/c26 ),
    .o({\u2_Display/add128/c27 ,\u2_Display/n4173 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u27  (
    .a(\u2_Display/n4143 ),
    .b(1'b1),
    .c(\u2_Display/add128/c27 ),
    .o({\u2_Display/add128/c28 ,\u2_Display/n4173 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u28  (
    .a(\u2_Display/n4142 ),
    .b(1'b1),
    .c(\u2_Display/add128/c28 ),
    .o({\u2_Display/add128/c29 ,\u2_Display/n4173 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u29  (
    .a(\u2_Display/n4141 ),
    .b(1'b1),
    .c(\u2_Display/add128/c29 ),
    .o({\u2_Display/add128/c30 ,\u2_Display/n4173 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u3  (
    .a(\u2_Display/n4167 ),
    .b(1'b1),
    .c(\u2_Display/add128/c3 ),
    .o({\u2_Display/add128/c4 ,\u2_Display/n4173 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u30  (
    .a(\u2_Display/n4140 ),
    .b(1'b1),
    .c(\u2_Display/add128/c30 ),
    .o({\u2_Display/add128/c31 ,\u2_Display/n4173 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u31  (
    .a(\u2_Display/n4139 ),
    .b(1'b1),
    .c(\u2_Display/add128/c31 ),
    .o({open_n951,\u2_Display/n4173 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u4  (
    .a(\u2_Display/n4166 ),
    .b(1'b1),
    .c(\u2_Display/add128/c4 ),
    .o({\u2_Display/add128/c5 ,\u2_Display/n4173 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u5  (
    .a(\u2_Display/n4165 ),
    .b(1'b1),
    .c(\u2_Display/add128/c5 ),
    .o({\u2_Display/add128/c6 ,\u2_Display/n4173 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u6  (
    .a(\u2_Display/n4164 ),
    .b(1'b1),
    .c(\u2_Display/add128/c6 ),
    .o({\u2_Display/add128/c7 ,\u2_Display/n4173 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u7  (
    .a(\u2_Display/n4163 ),
    .b(1'b1),
    .c(\u2_Display/add128/c7 ),
    .o({\u2_Display/add128/c8 ,\u2_Display/n4173 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u8  (
    .a(\u2_Display/n4162 ),
    .b(1'b1),
    .c(\u2_Display/add128/c8 ),
    .o({\u2_Display/add128/c9 ,\u2_Display/n4173 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add128/u9  (
    .a(\u2_Display/n4161 ),
    .b(1'b1),
    .c(\u2_Display/add128/c9 ),
    .o({\u2_Display/add128/c10 ,\u2_Display/n4173 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add128/ucin  (
    .a(1'b1),
    .o({\u2_Display/add128/c0 ,open_n954}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u0  (
    .a(\u2_Display/n4205 ),
    .b(1'b1),
    .c(\u2_Display/add129/c0 ),
    .o({\u2_Display/add129/c1 ,\u2_Display/n4208 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u1  (
    .a(\u2_Display/n4204 ),
    .b(1'b1),
    .c(\u2_Display/add129/c1 ),
    .o({\u2_Display/add129/c2 ,\u2_Display/n4208 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u10  (
    .a(\u2_Display/n4195 ),
    .b(1'b1),
    .c(\u2_Display/add129/c10 ),
    .o({\u2_Display/add129/c11 ,\u2_Display/n4208 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u11  (
    .a(\u2_Display/n4194 ),
    .b(1'b1),
    .c(\u2_Display/add129/c11 ),
    .o({\u2_Display/add129/c12 ,\u2_Display/n4208 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u12  (
    .a(\u2_Display/n4193 ),
    .b(1'b1),
    .c(\u2_Display/add129/c12 ),
    .o({\u2_Display/add129/c13 ,\u2_Display/n4208 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u13  (
    .a(\u2_Display/n4192 ),
    .b(1'b1),
    .c(\u2_Display/add129/c13 ),
    .o({\u2_Display/add129/c14 ,\u2_Display/n4208 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u14  (
    .a(\u2_Display/n4191 ),
    .b(1'b1),
    .c(\u2_Display/add129/c14 ),
    .o({\u2_Display/add129/c15 ,\u2_Display/n4208 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u15  (
    .a(\u2_Display/n4190 ),
    .b(1'b0),
    .c(\u2_Display/add129/c15 ),
    .o({\u2_Display/add129/c16 ,\u2_Display/n4208 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u16  (
    .a(\u2_Display/n4189 ),
    .b(1'b1),
    .c(\u2_Display/add129/c16 ),
    .o({\u2_Display/add129/c17 ,\u2_Display/n4208 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u17  (
    .a(\u2_Display/n4188 ),
    .b(1'b1),
    .c(\u2_Display/add129/c17 ),
    .o({\u2_Display/add129/c18 ,\u2_Display/n4208 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u18  (
    .a(\u2_Display/n4187 ),
    .b(1'b0),
    .c(\u2_Display/add129/c18 ),
    .o({\u2_Display/add129/c19 ,\u2_Display/n4208 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u19  (
    .a(\u2_Display/n4186 ),
    .b(1'b0),
    .c(\u2_Display/add129/c19 ),
    .o({\u2_Display/add129/c20 ,\u2_Display/n4208 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u2  (
    .a(\u2_Display/n4203 ),
    .b(1'b1),
    .c(\u2_Display/add129/c2 ),
    .o({\u2_Display/add129/c3 ,\u2_Display/n4208 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u20  (
    .a(\u2_Display/n4185 ),
    .b(1'b1),
    .c(\u2_Display/add129/c20 ),
    .o({\u2_Display/add129/c21 ,\u2_Display/n4208 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u21  (
    .a(\u2_Display/n4184 ),
    .b(1'b1),
    .c(\u2_Display/add129/c21 ),
    .o({\u2_Display/add129/c22 ,\u2_Display/n4208 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u22  (
    .a(\u2_Display/n4183 ),
    .b(1'b1),
    .c(\u2_Display/add129/c22 ),
    .o({\u2_Display/add129/c23 ,\u2_Display/n4208 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u23  (
    .a(\u2_Display/n4182 ),
    .b(1'b1),
    .c(\u2_Display/add129/c23 ),
    .o({\u2_Display/add129/c24 ,\u2_Display/n4208 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u24  (
    .a(\u2_Display/n4181 ),
    .b(1'b1),
    .c(\u2_Display/add129/c24 ),
    .o({\u2_Display/add129/c25 ,\u2_Display/n4208 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u25  (
    .a(\u2_Display/n4180 ),
    .b(1'b1),
    .c(\u2_Display/add129/c25 ),
    .o({\u2_Display/add129/c26 ,\u2_Display/n4208 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u26  (
    .a(\u2_Display/n4179 ),
    .b(1'b1),
    .c(\u2_Display/add129/c26 ),
    .o({\u2_Display/add129/c27 ,\u2_Display/n4208 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u27  (
    .a(\u2_Display/n4178 ),
    .b(1'b1),
    .c(\u2_Display/add129/c27 ),
    .o({\u2_Display/add129/c28 ,\u2_Display/n4208 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u28  (
    .a(\u2_Display/n4177 ),
    .b(1'b1),
    .c(\u2_Display/add129/c28 ),
    .o({\u2_Display/add129/c29 ,\u2_Display/n4208 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u29  (
    .a(\u2_Display/n4176 ),
    .b(1'b1),
    .c(\u2_Display/add129/c29 ),
    .o({\u2_Display/add129/c30 ,\u2_Display/n4208 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u3  (
    .a(\u2_Display/n4202 ),
    .b(1'b1),
    .c(\u2_Display/add129/c3 ),
    .o({\u2_Display/add129/c4 ,\u2_Display/n4208 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u30  (
    .a(\u2_Display/n4175 ),
    .b(1'b1),
    .c(\u2_Display/add129/c30 ),
    .o({\u2_Display/add129/c31 ,\u2_Display/n4208 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u31  (
    .a(\u2_Display/n4174 ),
    .b(1'b1),
    .c(\u2_Display/add129/c31 ),
    .o({open_n955,\u2_Display/n4208 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u4  (
    .a(\u2_Display/n4201 ),
    .b(1'b1),
    .c(\u2_Display/add129/c4 ),
    .o({\u2_Display/add129/c5 ,\u2_Display/n4208 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u5  (
    .a(\u2_Display/n4200 ),
    .b(1'b1),
    .c(\u2_Display/add129/c5 ),
    .o({\u2_Display/add129/c6 ,\u2_Display/n4208 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u6  (
    .a(\u2_Display/n4199 ),
    .b(1'b1),
    .c(\u2_Display/add129/c6 ),
    .o({\u2_Display/add129/c7 ,\u2_Display/n4208 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u7  (
    .a(\u2_Display/n4198 ),
    .b(1'b1),
    .c(\u2_Display/add129/c7 ),
    .o({\u2_Display/add129/c8 ,\u2_Display/n4208 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u8  (
    .a(\u2_Display/n4197 ),
    .b(1'b1),
    .c(\u2_Display/add129/c8 ),
    .o({\u2_Display/add129/c9 ,\u2_Display/n4208 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add129/u9  (
    .a(\u2_Display/n4196 ),
    .b(1'b1),
    .c(\u2_Display/add129/c9 ),
    .o({\u2_Display/add129/c10 ,\u2_Display/n4208 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add129/ucin  (
    .a(1'b1),
    .o({\u2_Display/add129/c0 ,open_n958}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u0  (
    .a(\u2_Display/n4240 ),
    .b(1'b1),
    .c(\u2_Display/add130/c0 ),
    .o({\u2_Display/add130/c1 ,\u2_Display/n4243 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u1  (
    .a(\u2_Display/n4239 ),
    .b(1'b1),
    .c(\u2_Display/add130/c1 ),
    .o({\u2_Display/add130/c2 ,\u2_Display/n4243 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u10  (
    .a(\u2_Display/n4230 ),
    .b(1'b1),
    .c(\u2_Display/add130/c10 ),
    .o({\u2_Display/add130/c11 ,\u2_Display/n4243 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u11  (
    .a(\u2_Display/n4229 ),
    .b(1'b1),
    .c(\u2_Display/add130/c11 ),
    .o({\u2_Display/add130/c12 ,\u2_Display/n4243 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u12  (
    .a(\u2_Display/n4228 ),
    .b(1'b1),
    .c(\u2_Display/add130/c12 ),
    .o({\u2_Display/add130/c13 ,\u2_Display/n4243 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u13  (
    .a(\u2_Display/n4227 ),
    .b(1'b1),
    .c(\u2_Display/add130/c13 ),
    .o({\u2_Display/add130/c14 ,\u2_Display/n4243 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u14  (
    .a(\u2_Display/n4226 ),
    .b(1'b0),
    .c(\u2_Display/add130/c14 ),
    .o({\u2_Display/add130/c15 ,\u2_Display/n4243 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u15  (
    .a(\u2_Display/n4225 ),
    .b(1'b1),
    .c(\u2_Display/add130/c15 ),
    .o({\u2_Display/add130/c16 ,\u2_Display/n4243 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u16  (
    .a(\u2_Display/n4224 ),
    .b(1'b1),
    .c(\u2_Display/add130/c16 ),
    .o({\u2_Display/add130/c17 ,\u2_Display/n4243 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u17  (
    .a(\u2_Display/n4223 ),
    .b(1'b0),
    .c(\u2_Display/add130/c17 ),
    .o({\u2_Display/add130/c18 ,\u2_Display/n4243 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u18  (
    .a(\u2_Display/n4222 ),
    .b(1'b0),
    .c(\u2_Display/add130/c18 ),
    .o({\u2_Display/add130/c19 ,\u2_Display/n4243 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u19  (
    .a(\u2_Display/n4221 ),
    .b(1'b1),
    .c(\u2_Display/add130/c19 ),
    .o({\u2_Display/add130/c20 ,\u2_Display/n4243 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u2  (
    .a(\u2_Display/n4238 ),
    .b(1'b1),
    .c(\u2_Display/add130/c2 ),
    .o({\u2_Display/add130/c3 ,\u2_Display/n4243 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u20  (
    .a(\u2_Display/n4220 ),
    .b(1'b1),
    .c(\u2_Display/add130/c20 ),
    .o({\u2_Display/add130/c21 ,\u2_Display/n4243 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u21  (
    .a(\u2_Display/n4219 ),
    .b(1'b1),
    .c(\u2_Display/add130/c21 ),
    .o({\u2_Display/add130/c22 ,\u2_Display/n4243 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u22  (
    .a(\u2_Display/n4218 ),
    .b(1'b1),
    .c(\u2_Display/add130/c22 ),
    .o({\u2_Display/add130/c23 ,\u2_Display/n4243 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u23  (
    .a(\u2_Display/n4217 ),
    .b(1'b1),
    .c(\u2_Display/add130/c23 ),
    .o({\u2_Display/add130/c24 ,\u2_Display/n4243 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u24  (
    .a(\u2_Display/n4216 ),
    .b(1'b1),
    .c(\u2_Display/add130/c24 ),
    .o({\u2_Display/add130/c25 ,\u2_Display/n4243 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u25  (
    .a(\u2_Display/n4215 ),
    .b(1'b1),
    .c(\u2_Display/add130/c25 ),
    .o({\u2_Display/add130/c26 ,\u2_Display/n4243 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u26  (
    .a(\u2_Display/n4214 ),
    .b(1'b1),
    .c(\u2_Display/add130/c26 ),
    .o({\u2_Display/add130/c27 ,\u2_Display/n4243 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u27  (
    .a(\u2_Display/n4213 ),
    .b(1'b1),
    .c(\u2_Display/add130/c27 ),
    .o({\u2_Display/add130/c28 ,\u2_Display/n4243 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u28  (
    .a(\u2_Display/n4212 ),
    .b(1'b1),
    .c(\u2_Display/add130/c28 ),
    .o({\u2_Display/add130/c29 ,\u2_Display/n4243 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u29  (
    .a(\u2_Display/n4211 ),
    .b(1'b1),
    .c(\u2_Display/add130/c29 ),
    .o({\u2_Display/add130/c30 ,\u2_Display/n4243 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u3  (
    .a(\u2_Display/n4237 ),
    .b(1'b1),
    .c(\u2_Display/add130/c3 ),
    .o({\u2_Display/add130/c4 ,\u2_Display/n4243 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u30  (
    .a(\u2_Display/n4210 ),
    .b(1'b1),
    .c(\u2_Display/add130/c30 ),
    .o({\u2_Display/add130/c31 ,\u2_Display/n4243 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u31  (
    .a(\u2_Display/n4209 ),
    .b(1'b1),
    .c(\u2_Display/add130/c31 ),
    .o({open_n959,\u2_Display/n4243 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u4  (
    .a(\u2_Display/n4236 ),
    .b(1'b1),
    .c(\u2_Display/add130/c4 ),
    .o({\u2_Display/add130/c5 ,\u2_Display/n4243 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u5  (
    .a(\u2_Display/n4235 ),
    .b(1'b1),
    .c(\u2_Display/add130/c5 ),
    .o({\u2_Display/add130/c6 ,\u2_Display/n4243 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u6  (
    .a(\u2_Display/n4234 ),
    .b(1'b1),
    .c(\u2_Display/add130/c6 ),
    .o({\u2_Display/add130/c7 ,\u2_Display/n4243 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u7  (
    .a(\u2_Display/n4233 ),
    .b(1'b1),
    .c(\u2_Display/add130/c7 ),
    .o({\u2_Display/add130/c8 ,\u2_Display/n4243 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u8  (
    .a(\u2_Display/n4232 ),
    .b(1'b1),
    .c(\u2_Display/add130/c8 ),
    .o({\u2_Display/add130/c9 ,\u2_Display/n4243 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add130/u9  (
    .a(\u2_Display/n4231 ),
    .b(1'b1),
    .c(\u2_Display/add130/c9 ),
    .o({\u2_Display/add130/c10 ,\u2_Display/n4243 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add130/ucin  (
    .a(1'b1),
    .o({\u2_Display/add130/c0 ,open_n962}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u0  (
    .a(\u2_Display/n4275 ),
    .b(1'b1),
    .c(\u2_Display/add131/c0 ),
    .o({\u2_Display/add131/c1 ,\u2_Display/n4278 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u1  (
    .a(\u2_Display/n4274 ),
    .b(1'b1),
    .c(\u2_Display/add131/c1 ),
    .o({\u2_Display/add131/c2 ,\u2_Display/n4278 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u10  (
    .a(\u2_Display/n4265 ),
    .b(1'b1),
    .c(\u2_Display/add131/c10 ),
    .o({\u2_Display/add131/c11 ,\u2_Display/n4278 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u11  (
    .a(\u2_Display/n4264 ),
    .b(1'b1),
    .c(\u2_Display/add131/c11 ),
    .o({\u2_Display/add131/c12 ,\u2_Display/n4278 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u12  (
    .a(\u2_Display/n4263 ),
    .b(1'b1),
    .c(\u2_Display/add131/c12 ),
    .o({\u2_Display/add131/c13 ,\u2_Display/n4278 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u13  (
    .a(\u2_Display/n4262 ),
    .b(1'b0),
    .c(\u2_Display/add131/c13 ),
    .o({\u2_Display/add131/c14 ,\u2_Display/n4278 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u14  (
    .a(\u2_Display/n4261 ),
    .b(1'b1),
    .c(\u2_Display/add131/c14 ),
    .o({\u2_Display/add131/c15 ,\u2_Display/n4278 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u15  (
    .a(\u2_Display/n4260 ),
    .b(1'b1),
    .c(\u2_Display/add131/c15 ),
    .o({\u2_Display/add131/c16 ,\u2_Display/n4278 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u16  (
    .a(\u2_Display/n4259 ),
    .b(1'b0),
    .c(\u2_Display/add131/c16 ),
    .o({\u2_Display/add131/c17 ,\u2_Display/n4278 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u17  (
    .a(\u2_Display/n4258 ),
    .b(1'b0),
    .c(\u2_Display/add131/c17 ),
    .o({\u2_Display/add131/c18 ,\u2_Display/n4278 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u18  (
    .a(\u2_Display/n4257 ),
    .b(1'b1),
    .c(\u2_Display/add131/c18 ),
    .o({\u2_Display/add131/c19 ,\u2_Display/n4278 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u19  (
    .a(\u2_Display/n4256 ),
    .b(1'b1),
    .c(\u2_Display/add131/c19 ),
    .o({\u2_Display/add131/c20 ,\u2_Display/n4278 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u2  (
    .a(\u2_Display/n4273 ),
    .b(1'b1),
    .c(\u2_Display/add131/c2 ),
    .o({\u2_Display/add131/c3 ,\u2_Display/n4278 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u20  (
    .a(\u2_Display/n4255 ),
    .b(1'b1),
    .c(\u2_Display/add131/c20 ),
    .o({\u2_Display/add131/c21 ,\u2_Display/n4278 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u21  (
    .a(\u2_Display/n4254 ),
    .b(1'b1),
    .c(\u2_Display/add131/c21 ),
    .o({\u2_Display/add131/c22 ,\u2_Display/n4278 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u22  (
    .a(\u2_Display/n4253 ),
    .b(1'b1),
    .c(\u2_Display/add131/c22 ),
    .o({\u2_Display/add131/c23 ,\u2_Display/n4278 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u23  (
    .a(\u2_Display/n4252 ),
    .b(1'b1),
    .c(\u2_Display/add131/c23 ),
    .o({\u2_Display/add131/c24 ,\u2_Display/n4278 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u24  (
    .a(\u2_Display/n4251 ),
    .b(1'b1),
    .c(\u2_Display/add131/c24 ),
    .o({\u2_Display/add131/c25 ,\u2_Display/n4278 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u25  (
    .a(\u2_Display/n4250 ),
    .b(1'b1),
    .c(\u2_Display/add131/c25 ),
    .o({\u2_Display/add131/c26 ,\u2_Display/n4278 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u26  (
    .a(\u2_Display/n4249 ),
    .b(1'b1),
    .c(\u2_Display/add131/c26 ),
    .o({\u2_Display/add131/c27 ,\u2_Display/n4278 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u27  (
    .a(\u2_Display/n4248 ),
    .b(1'b1),
    .c(\u2_Display/add131/c27 ),
    .o({\u2_Display/add131/c28 ,\u2_Display/n4278 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u28  (
    .a(\u2_Display/n4247 ),
    .b(1'b1),
    .c(\u2_Display/add131/c28 ),
    .o({\u2_Display/add131/c29 ,\u2_Display/n4278 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u29  (
    .a(\u2_Display/n4246 ),
    .b(1'b1),
    .c(\u2_Display/add131/c29 ),
    .o({\u2_Display/add131/c30 ,\u2_Display/n4278 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u3  (
    .a(\u2_Display/n4272 ),
    .b(1'b1),
    .c(\u2_Display/add131/c3 ),
    .o({\u2_Display/add131/c4 ,\u2_Display/n4278 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u30  (
    .a(\u2_Display/n4245 ),
    .b(1'b1),
    .c(\u2_Display/add131/c30 ),
    .o({\u2_Display/add131/c31 ,\u2_Display/n4278 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u31  (
    .a(\u2_Display/n4244 ),
    .b(1'b1),
    .c(\u2_Display/add131/c31 ),
    .o({open_n963,\u2_Display/n4278 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u4  (
    .a(\u2_Display/n4271 ),
    .b(1'b1),
    .c(\u2_Display/add131/c4 ),
    .o({\u2_Display/add131/c5 ,\u2_Display/n4278 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u5  (
    .a(\u2_Display/n4270 ),
    .b(1'b1),
    .c(\u2_Display/add131/c5 ),
    .o({\u2_Display/add131/c6 ,\u2_Display/n4278 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u6  (
    .a(\u2_Display/n4269 ),
    .b(1'b1),
    .c(\u2_Display/add131/c6 ),
    .o({\u2_Display/add131/c7 ,\u2_Display/n4278 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u7  (
    .a(\u2_Display/n4268 ),
    .b(1'b1),
    .c(\u2_Display/add131/c7 ),
    .o({\u2_Display/add131/c8 ,\u2_Display/n4278 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u8  (
    .a(\u2_Display/n4267 ),
    .b(1'b1),
    .c(\u2_Display/add131/c8 ),
    .o({\u2_Display/add131/c9 ,\u2_Display/n4278 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add131/u9  (
    .a(\u2_Display/n4266 ),
    .b(1'b1),
    .c(\u2_Display/add131/c9 ),
    .o({\u2_Display/add131/c10 ,\u2_Display/n4278 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add131/ucin  (
    .a(1'b1),
    .o({\u2_Display/add131/c0 ,open_n966}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u0  (
    .a(\u2_Display/n4310 ),
    .b(1'b1),
    .c(\u2_Display/add132/c0 ),
    .o({\u2_Display/add132/c1 ,\u2_Display/n4313 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u1  (
    .a(\u2_Display/n4309 ),
    .b(1'b1),
    .c(\u2_Display/add132/c1 ),
    .o({\u2_Display/add132/c2 ,\u2_Display/n4313 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u10  (
    .a(\u2_Display/n4300 ),
    .b(1'b1),
    .c(\u2_Display/add132/c10 ),
    .o({\u2_Display/add132/c11 ,\u2_Display/n4313 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u11  (
    .a(\u2_Display/n4299 ),
    .b(1'b1),
    .c(\u2_Display/add132/c11 ),
    .o({\u2_Display/add132/c12 ,\u2_Display/n4313 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u12  (
    .a(\u2_Display/n4298 ),
    .b(1'b0),
    .c(\u2_Display/add132/c12 ),
    .o({\u2_Display/add132/c13 ,\u2_Display/n4313 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u13  (
    .a(\u2_Display/n4297 ),
    .b(1'b1),
    .c(\u2_Display/add132/c13 ),
    .o({\u2_Display/add132/c14 ,\u2_Display/n4313 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u14  (
    .a(\u2_Display/n4296 ),
    .b(1'b1),
    .c(\u2_Display/add132/c14 ),
    .o({\u2_Display/add132/c15 ,\u2_Display/n4313 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u15  (
    .a(\u2_Display/n4295 ),
    .b(1'b0),
    .c(\u2_Display/add132/c15 ),
    .o({\u2_Display/add132/c16 ,\u2_Display/n4313 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u16  (
    .a(\u2_Display/n4294 ),
    .b(1'b0),
    .c(\u2_Display/add132/c16 ),
    .o({\u2_Display/add132/c17 ,\u2_Display/n4313 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u17  (
    .a(\u2_Display/n4293 ),
    .b(1'b1),
    .c(\u2_Display/add132/c17 ),
    .o({\u2_Display/add132/c18 ,\u2_Display/n4313 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u18  (
    .a(\u2_Display/n4292 ),
    .b(1'b1),
    .c(\u2_Display/add132/c18 ),
    .o({\u2_Display/add132/c19 ,\u2_Display/n4313 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u19  (
    .a(\u2_Display/n4291 ),
    .b(1'b1),
    .c(\u2_Display/add132/c19 ),
    .o({\u2_Display/add132/c20 ,\u2_Display/n4313 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u2  (
    .a(\u2_Display/n4308 ),
    .b(1'b1),
    .c(\u2_Display/add132/c2 ),
    .o({\u2_Display/add132/c3 ,\u2_Display/n4313 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u20  (
    .a(\u2_Display/n4290 ),
    .b(1'b1),
    .c(\u2_Display/add132/c20 ),
    .o({\u2_Display/add132/c21 ,\u2_Display/n4313 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u21  (
    .a(\u2_Display/n4289 ),
    .b(1'b1),
    .c(\u2_Display/add132/c21 ),
    .o({\u2_Display/add132/c22 ,\u2_Display/n4313 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u22  (
    .a(\u2_Display/n4288 ),
    .b(1'b1),
    .c(\u2_Display/add132/c22 ),
    .o({\u2_Display/add132/c23 ,\u2_Display/n4313 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u23  (
    .a(\u2_Display/n4287 ),
    .b(1'b1),
    .c(\u2_Display/add132/c23 ),
    .o({\u2_Display/add132/c24 ,\u2_Display/n4313 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u24  (
    .a(\u2_Display/n4286 ),
    .b(1'b1),
    .c(\u2_Display/add132/c24 ),
    .o({\u2_Display/add132/c25 ,\u2_Display/n4313 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u25  (
    .a(\u2_Display/n4285 ),
    .b(1'b1),
    .c(\u2_Display/add132/c25 ),
    .o({\u2_Display/add132/c26 ,\u2_Display/n4313 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u26  (
    .a(\u2_Display/n4284 ),
    .b(1'b1),
    .c(\u2_Display/add132/c26 ),
    .o({\u2_Display/add132/c27 ,\u2_Display/n4313 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u27  (
    .a(\u2_Display/n4283 ),
    .b(1'b1),
    .c(\u2_Display/add132/c27 ),
    .o({\u2_Display/add132/c28 ,\u2_Display/n4313 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u28  (
    .a(\u2_Display/n4282 ),
    .b(1'b1),
    .c(\u2_Display/add132/c28 ),
    .o({\u2_Display/add132/c29 ,\u2_Display/n4313 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u29  (
    .a(\u2_Display/n4281 ),
    .b(1'b1),
    .c(\u2_Display/add132/c29 ),
    .o({\u2_Display/add132/c30 ,\u2_Display/n4313 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u3  (
    .a(\u2_Display/n4307 ),
    .b(1'b1),
    .c(\u2_Display/add132/c3 ),
    .o({\u2_Display/add132/c4 ,\u2_Display/n4313 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u30  (
    .a(\u2_Display/n4280 ),
    .b(1'b1),
    .c(\u2_Display/add132/c30 ),
    .o({\u2_Display/add132/c31 ,\u2_Display/n4313 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u31  (
    .a(\u2_Display/n4279 ),
    .b(1'b1),
    .c(\u2_Display/add132/c31 ),
    .o({open_n967,\u2_Display/n4313 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u4  (
    .a(\u2_Display/n4306 ),
    .b(1'b1),
    .c(\u2_Display/add132/c4 ),
    .o({\u2_Display/add132/c5 ,\u2_Display/n4313 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u5  (
    .a(\u2_Display/n4305 ),
    .b(1'b1),
    .c(\u2_Display/add132/c5 ),
    .o({\u2_Display/add132/c6 ,\u2_Display/n4313 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u6  (
    .a(\u2_Display/n4304 ),
    .b(1'b1),
    .c(\u2_Display/add132/c6 ),
    .o({\u2_Display/add132/c7 ,\u2_Display/n4313 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u7  (
    .a(\u2_Display/n4303 ),
    .b(1'b1),
    .c(\u2_Display/add132/c7 ),
    .o({\u2_Display/add132/c8 ,\u2_Display/n4313 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u8  (
    .a(\u2_Display/n4302 ),
    .b(1'b1),
    .c(\u2_Display/add132/c8 ),
    .o({\u2_Display/add132/c9 ,\u2_Display/n4313 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add132/u9  (
    .a(\u2_Display/n4301 ),
    .b(1'b1),
    .c(\u2_Display/add132/c9 ),
    .o({\u2_Display/add132/c10 ,\u2_Display/n4313 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add132/ucin  (
    .a(1'b1),
    .o({\u2_Display/add132/c0 ,open_n970}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u0  (
    .a(\u2_Display/n4345 ),
    .b(1'b1),
    .c(\u2_Display/add133/c0 ),
    .o({\u2_Display/add133/c1 ,\u2_Display/n4348 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u1  (
    .a(\u2_Display/n4344 ),
    .b(1'b1),
    .c(\u2_Display/add133/c1 ),
    .o({\u2_Display/add133/c2 ,\u2_Display/n4348 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u10  (
    .a(\u2_Display/n4335 ),
    .b(1'b1),
    .c(\u2_Display/add133/c10 ),
    .o({\u2_Display/add133/c11 ,\u2_Display/n4348 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u11  (
    .a(\u2_Display/n4334 ),
    .b(1'b0),
    .c(\u2_Display/add133/c11 ),
    .o({\u2_Display/add133/c12 ,\u2_Display/n4348 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u12  (
    .a(\u2_Display/n4333 ),
    .b(1'b1),
    .c(\u2_Display/add133/c12 ),
    .o({\u2_Display/add133/c13 ,\u2_Display/n4348 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u13  (
    .a(\u2_Display/n4332 ),
    .b(1'b1),
    .c(\u2_Display/add133/c13 ),
    .o({\u2_Display/add133/c14 ,\u2_Display/n4348 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u14  (
    .a(\u2_Display/n4331 ),
    .b(1'b0),
    .c(\u2_Display/add133/c14 ),
    .o({\u2_Display/add133/c15 ,\u2_Display/n4348 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u15  (
    .a(\u2_Display/n4330 ),
    .b(1'b0),
    .c(\u2_Display/add133/c15 ),
    .o({\u2_Display/add133/c16 ,\u2_Display/n4348 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u16  (
    .a(\u2_Display/n4329 ),
    .b(1'b1),
    .c(\u2_Display/add133/c16 ),
    .o({\u2_Display/add133/c17 ,\u2_Display/n4348 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u17  (
    .a(\u2_Display/n4328 ),
    .b(1'b1),
    .c(\u2_Display/add133/c17 ),
    .o({\u2_Display/add133/c18 ,\u2_Display/n4348 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u18  (
    .a(\u2_Display/n4327 ),
    .b(1'b1),
    .c(\u2_Display/add133/c18 ),
    .o({\u2_Display/add133/c19 ,\u2_Display/n4348 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u19  (
    .a(\u2_Display/n4326 ),
    .b(1'b1),
    .c(\u2_Display/add133/c19 ),
    .o({\u2_Display/add133/c20 ,\u2_Display/n4348 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u2  (
    .a(\u2_Display/n4343 ),
    .b(1'b1),
    .c(\u2_Display/add133/c2 ),
    .o({\u2_Display/add133/c3 ,\u2_Display/n4348 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u20  (
    .a(\u2_Display/n4325 ),
    .b(1'b1),
    .c(\u2_Display/add133/c20 ),
    .o({\u2_Display/add133/c21 ,\u2_Display/n4348 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u21  (
    .a(\u2_Display/n4324 ),
    .b(1'b1),
    .c(\u2_Display/add133/c21 ),
    .o({\u2_Display/add133/c22 ,\u2_Display/n4348 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u22  (
    .a(\u2_Display/n4323 ),
    .b(1'b1),
    .c(\u2_Display/add133/c22 ),
    .o({\u2_Display/add133/c23 ,\u2_Display/n4348 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u23  (
    .a(\u2_Display/n4322 ),
    .b(1'b1),
    .c(\u2_Display/add133/c23 ),
    .o({\u2_Display/add133/c24 ,\u2_Display/n4348 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u24  (
    .a(\u2_Display/n4321 ),
    .b(1'b1),
    .c(\u2_Display/add133/c24 ),
    .o({\u2_Display/add133/c25 ,\u2_Display/n4348 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u25  (
    .a(\u2_Display/n4320 ),
    .b(1'b1),
    .c(\u2_Display/add133/c25 ),
    .o({\u2_Display/add133/c26 ,\u2_Display/n4348 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u26  (
    .a(\u2_Display/n4319 ),
    .b(1'b1),
    .c(\u2_Display/add133/c26 ),
    .o({\u2_Display/add133/c27 ,\u2_Display/n4348 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u27  (
    .a(\u2_Display/n4318 ),
    .b(1'b1),
    .c(\u2_Display/add133/c27 ),
    .o({\u2_Display/add133/c28 ,\u2_Display/n4348 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u28  (
    .a(\u2_Display/n4317 ),
    .b(1'b1),
    .c(\u2_Display/add133/c28 ),
    .o({\u2_Display/add133/c29 ,\u2_Display/n4348 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u29  (
    .a(\u2_Display/n4316 ),
    .b(1'b1),
    .c(\u2_Display/add133/c29 ),
    .o({\u2_Display/add133/c30 ,\u2_Display/n4348 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u3  (
    .a(\u2_Display/n4342 ),
    .b(1'b1),
    .c(\u2_Display/add133/c3 ),
    .o({\u2_Display/add133/c4 ,\u2_Display/n4348 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u30  (
    .a(\u2_Display/n4315 ),
    .b(1'b1),
    .c(\u2_Display/add133/c30 ),
    .o({\u2_Display/add133/c31 ,\u2_Display/n4348 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u31  (
    .a(\u2_Display/n4314 ),
    .b(1'b1),
    .c(\u2_Display/add133/c31 ),
    .o({open_n971,\u2_Display/n4348 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u4  (
    .a(\u2_Display/n4341 ),
    .b(1'b1),
    .c(\u2_Display/add133/c4 ),
    .o({\u2_Display/add133/c5 ,\u2_Display/n4348 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u5  (
    .a(\u2_Display/n4340 ),
    .b(1'b1),
    .c(\u2_Display/add133/c5 ),
    .o({\u2_Display/add133/c6 ,\u2_Display/n4348 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u6  (
    .a(\u2_Display/n4339 ),
    .b(1'b1),
    .c(\u2_Display/add133/c6 ),
    .o({\u2_Display/add133/c7 ,\u2_Display/n4348 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u7  (
    .a(\u2_Display/n4338 ),
    .b(1'b1),
    .c(\u2_Display/add133/c7 ),
    .o({\u2_Display/add133/c8 ,\u2_Display/n4348 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u8  (
    .a(\u2_Display/n4337 ),
    .b(1'b1),
    .c(\u2_Display/add133/c8 ),
    .o({\u2_Display/add133/c9 ,\u2_Display/n4348 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add133/u9  (
    .a(\u2_Display/n4336 ),
    .b(1'b1),
    .c(\u2_Display/add133/c9 ),
    .o({\u2_Display/add133/c10 ,\u2_Display/n4348 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add133/ucin  (
    .a(1'b1),
    .o({\u2_Display/add133/c0 ,open_n974}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u0  (
    .a(\u2_Display/n4380 ),
    .b(1'b1),
    .c(\u2_Display/add134/c0 ),
    .o({\u2_Display/add134/c1 ,\u2_Display/n4383 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u1  (
    .a(\u2_Display/n4379 ),
    .b(1'b1),
    .c(\u2_Display/add134/c1 ),
    .o({\u2_Display/add134/c2 ,\u2_Display/n4383 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u10  (
    .a(\u2_Display/n4370 ),
    .b(1'b0),
    .c(\u2_Display/add134/c10 ),
    .o({\u2_Display/add134/c11 ,\u2_Display/n4383 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u11  (
    .a(\u2_Display/n4369 ),
    .b(1'b1),
    .c(\u2_Display/add134/c11 ),
    .o({\u2_Display/add134/c12 ,\u2_Display/n4383 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u12  (
    .a(\u2_Display/n4368 ),
    .b(1'b1),
    .c(\u2_Display/add134/c12 ),
    .o({\u2_Display/add134/c13 ,\u2_Display/n4383 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u13  (
    .a(\u2_Display/n4367 ),
    .b(1'b0),
    .c(\u2_Display/add134/c13 ),
    .o({\u2_Display/add134/c14 ,\u2_Display/n4383 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u14  (
    .a(\u2_Display/n4366 ),
    .b(1'b0),
    .c(\u2_Display/add134/c14 ),
    .o({\u2_Display/add134/c15 ,\u2_Display/n4383 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u15  (
    .a(\u2_Display/n4365 ),
    .b(1'b1),
    .c(\u2_Display/add134/c15 ),
    .o({\u2_Display/add134/c16 ,\u2_Display/n4383 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u16  (
    .a(\u2_Display/n4364 ),
    .b(1'b1),
    .c(\u2_Display/add134/c16 ),
    .o({\u2_Display/add134/c17 ,\u2_Display/n4383 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u17  (
    .a(\u2_Display/n4363 ),
    .b(1'b1),
    .c(\u2_Display/add134/c17 ),
    .o({\u2_Display/add134/c18 ,\u2_Display/n4383 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u18  (
    .a(\u2_Display/n4362 ),
    .b(1'b1),
    .c(\u2_Display/add134/c18 ),
    .o({\u2_Display/add134/c19 ,\u2_Display/n4383 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u19  (
    .a(\u2_Display/n4361 ),
    .b(1'b1),
    .c(\u2_Display/add134/c19 ),
    .o({\u2_Display/add134/c20 ,\u2_Display/n4383 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u2  (
    .a(\u2_Display/n4378 ),
    .b(1'b1),
    .c(\u2_Display/add134/c2 ),
    .o({\u2_Display/add134/c3 ,\u2_Display/n4383 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u20  (
    .a(\u2_Display/n4360 ),
    .b(1'b1),
    .c(\u2_Display/add134/c20 ),
    .o({\u2_Display/add134/c21 ,\u2_Display/n4383 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u21  (
    .a(\u2_Display/n4359 ),
    .b(1'b1),
    .c(\u2_Display/add134/c21 ),
    .o({\u2_Display/add134/c22 ,\u2_Display/n4383 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u22  (
    .a(\u2_Display/n4358 ),
    .b(1'b1),
    .c(\u2_Display/add134/c22 ),
    .o({\u2_Display/add134/c23 ,\u2_Display/n4383 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u23  (
    .a(\u2_Display/n4357 ),
    .b(1'b1),
    .c(\u2_Display/add134/c23 ),
    .o({\u2_Display/add134/c24 ,\u2_Display/n4383 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u24  (
    .a(\u2_Display/n4356 ),
    .b(1'b1),
    .c(\u2_Display/add134/c24 ),
    .o({\u2_Display/add134/c25 ,\u2_Display/n4383 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u25  (
    .a(\u2_Display/n4355 ),
    .b(1'b1),
    .c(\u2_Display/add134/c25 ),
    .o({\u2_Display/add134/c26 ,\u2_Display/n4383 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u26  (
    .a(\u2_Display/n4354 ),
    .b(1'b1),
    .c(\u2_Display/add134/c26 ),
    .o({\u2_Display/add134/c27 ,\u2_Display/n4383 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u27  (
    .a(\u2_Display/n4353 ),
    .b(1'b1),
    .c(\u2_Display/add134/c27 ),
    .o({\u2_Display/add134/c28 ,\u2_Display/n4383 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u28  (
    .a(\u2_Display/n4352 ),
    .b(1'b1),
    .c(\u2_Display/add134/c28 ),
    .o({\u2_Display/add134/c29 ,\u2_Display/n4383 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u29  (
    .a(\u2_Display/n4351 ),
    .b(1'b1),
    .c(\u2_Display/add134/c29 ),
    .o({\u2_Display/add134/c30 ,\u2_Display/n4383 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u3  (
    .a(\u2_Display/n4377 ),
    .b(1'b1),
    .c(\u2_Display/add134/c3 ),
    .o({\u2_Display/add134/c4 ,\u2_Display/n4383 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u30  (
    .a(\u2_Display/n4350 ),
    .b(1'b1),
    .c(\u2_Display/add134/c30 ),
    .o({\u2_Display/add134/c31 ,\u2_Display/n4383 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u31  (
    .a(\u2_Display/n4349 ),
    .b(1'b1),
    .c(\u2_Display/add134/c31 ),
    .o({open_n975,\u2_Display/n4383 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u4  (
    .a(\u2_Display/n4376 ),
    .b(1'b1),
    .c(\u2_Display/add134/c4 ),
    .o({\u2_Display/add134/c5 ,\u2_Display/n4383 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u5  (
    .a(\u2_Display/n4375 ),
    .b(1'b1),
    .c(\u2_Display/add134/c5 ),
    .o({\u2_Display/add134/c6 ,\u2_Display/n4383 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u6  (
    .a(\u2_Display/n4374 ),
    .b(1'b1),
    .c(\u2_Display/add134/c6 ),
    .o({\u2_Display/add134/c7 ,\u2_Display/n4383 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u7  (
    .a(\u2_Display/n4373 ),
    .b(1'b1),
    .c(\u2_Display/add134/c7 ),
    .o({\u2_Display/add134/c8 ,\u2_Display/n4383 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u8  (
    .a(\u2_Display/n4372 ),
    .b(1'b1),
    .c(\u2_Display/add134/c8 ),
    .o({\u2_Display/add134/c9 ,\u2_Display/n4383 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add134/u9  (
    .a(\u2_Display/n4371 ),
    .b(1'b1),
    .c(\u2_Display/add134/c9 ),
    .o({\u2_Display/add134/c10 ,\u2_Display/n4383 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add134/ucin  (
    .a(1'b1),
    .o({\u2_Display/add134/c0 ,open_n978}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u0  (
    .a(\u2_Display/n4415 ),
    .b(1'b1),
    .c(\u2_Display/add135/c0 ),
    .o({\u2_Display/add135/c1 ,\u2_Display/n4418 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u1  (
    .a(\u2_Display/n4414 ),
    .b(1'b1),
    .c(\u2_Display/add135/c1 ),
    .o({\u2_Display/add135/c2 ,\u2_Display/n4418 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u10  (
    .a(\u2_Display/n4405 ),
    .b(1'b1),
    .c(\u2_Display/add135/c10 ),
    .o({\u2_Display/add135/c11 ,\u2_Display/n4418 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u11  (
    .a(\u2_Display/n4404 ),
    .b(1'b1),
    .c(\u2_Display/add135/c11 ),
    .o({\u2_Display/add135/c12 ,\u2_Display/n4418 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u12  (
    .a(\u2_Display/n4403 ),
    .b(1'b0),
    .c(\u2_Display/add135/c12 ),
    .o({\u2_Display/add135/c13 ,\u2_Display/n4418 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u13  (
    .a(\u2_Display/n4402 ),
    .b(1'b0),
    .c(\u2_Display/add135/c13 ),
    .o({\u2_Display/add135/c14 ,\u2_Display/n4418 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u14  (
    .a(\u2_Display/n4401 ),
    .b(1'b1),
    .c(\u2_Display/add135/c14 ),
    .o({\u2_Display/add135/c15 ,\u2_Display/n4418 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u15  (
    .a(\u2_Display/n4400 ),
    .b(1'b1),
    .c(\u2_Display/add135/c15 ),
    .o({\u2_Display/add135/c16 ,\u2_Display/n4418 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u16  (
    .a(\u2_Display/n4399 ),
    .b(1'b1),
    .c(\u2_Display/add135/c16 ),
    .o({\u2_Display/add135/c17 ,\u2_Display/n4418 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u17  (
    .a(\u2_Display/n4398 ),
    .b(1'b1),
    .c(\u2_Display/add135/c17 ),
    .o({\u2_Display/add135/c18 ,\u2_Display/n4418 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u18  (
    .a(\u2_Display/n4397 ),
    .b(1'b1),
    .c(\u2_Display/add135/c18 ),
    .o({\u2_Display/add135/c19 ,\u2_Display/n4418 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u19  (
    .a(\u2_Display/n4396 ),
    .b(1'b1),
    .c(\u2_Display/add135/c19 ),
    .o({\u2_Display/add135/c20 ,\u2_Display/n4418 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u2  (
    .a(\u2_Display/n4413 ),
    .b(1'b1),
    .c(\u2_Display/add135/c2 ),
    .o({\u2_Display/add135/c3 ,\u2_Display/n4418 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u20  (
    .a(\u2_Display/n4395 ),
    .b(1'b1),
    .c(\u2_Display/add135/c20 ),
    .o({\u2_Display/add135/c21 ,\u2_Display/n4418 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u21  (
    .a(\u2_Display/n4394 ),
    .b(1'b1),
    .c(\u2_Display/add135/c21 ),
    .o({\u2_Display/add135/c22 ,\u2_Display/n4418 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u22  (
    .a(\u2_Display/n4393 ),
    .b(1'b1),
    .c(\u2_Display/add135/c22 ),
    .o({\u2_Display/add135/c23 ,\u2_Display/n4418 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u23  (
    .a(\u2_Display/n4392 ),
    .b(1'b1),
    .c(\u2_Display/add135/c23 ),
    .o({\u2_Display/add135/c24 ,\u2_Display/n4418 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u24  (
    .a(\u2_Display/n4391 ),
    .b(1'b1),
    .c(\u2_Display/add135/c24 ),
    .o({\u2_Display/add135/c25 ,\u2_Display/n4418 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u25  (
    .a(\u2_Display/n4390 ),
    .b(1'b1),
    .c(\u2_Display/add135/c25 ),
    .o({\u2_Display/add135/c26 ,\u2_Display/n4418 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u26  (
    .a(\u2_Display/n4389 ),
    .b(1'b1),
    .c(\u2_Display/add135/c26 ),
    .o({\u2_Display/add135/c27 ,\u2_Display/n4418 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u27  (
    .a(\u2_Display/n4388 ),
    .b(1'b1),
    .c(\u2_Display/add135/c27 ),
    .o({\u2_Display/add135/c28 ,\u2_Display/n4418 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u28  (
    .a(\u2_Display/n4387 ),
    .b(1'b1),
    .c(\u2_Display/add135/c28 ),
    .o({\u2_Display/add135/c29 ,\u2_Display/n4418 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u29  (
    .a(\u2_Display/n4386 ),
    .b(1'b1),
    .c(\u2_Display/add135/c29 ),
    .o({\u2_Display/add135/c30 ,\u2_Display/n4418 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u3  (
    .a(\u2_Display/n4412 ),
    .b(1'b1),
    .c(\u2_Display/add135/c3 ),
    .o({\u2_Display/add135/c4 ,\u2_Display/n4418 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u30  (
    .a(\u2_Display/n4385 ),
    .b(1'b1),
    .c(\u2_Display/add135/c30 ),
    .o({\u2_Display/add135/c31 ,\u2_Display/n4418 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u31  (
    .a(\u2_Display/n4384 ),
    .b(1'b1),
    .c(\u2_Display/add135/c31 ),
    .o({open_n979,\u2_Display/n4418 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u4  (
    .a(\u2_Display/n4411 ),
    .b(1'b1),
    .c(\u2_Display/add135/c4 ),
    .o({\u2_Display/add135/c5 ,\u2_Display/n4418 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u5  (
    .a(\u2_Display/n4410 ),
    .b(1'b1),
    .c(\u2_Display/add135/c5 ),
    .o({\u2_Display/add135/c6 ,\u2_Display/n4418 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u6  (
    .a(\u2_Display/n4409 ),
    .b(1'b1),
    .c(\u2_Display/add135/c6 ),
    .o({\u2_Display/add135/c7 ,\u2_Display/n4418 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u7  (
    .a(\u2_Display/n4408 ),
    .b(1'b1),
    .c(\u2_Display/add135/c7 ),
    .o({\u2_Display/add135/c8 ,\u2_Display/n4418 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u8  (
    .a(\u2_Display/n4407 ),
    .b(1'b1),
    .c(\u2_Display/add135/c8 ),
    .o({\u2_Display/add135/c9 ,\u2_Display/n4418 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add135/u9  (
    .a(\u2_Display/n4406 ),
    .b(1'b0),
    .c(\u2_Display/add135/c9 ),
    .o({\u2_Display/add135/c10 ,\u2_Display/n4418 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add135/ucin  (
    .a(1'b1),
    .o({\u2_Display/add135/c0 ,open_n982}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u0  (
    .a(\u2_Display/n4450 ),
    .b(1'b1),
    .c(\u2_Display/add136/c0 ),
    .o({\u2_Display/add136/c1 ,\u2_Display/n4453 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u1  (
    .a(\u2_Display/n4449 ),
    .b(1'b1),
    .c(\u2_Display/add136/c1 ),
    .o({\u2_Display/add136/c2 ,\u2_Display/n4453 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u10  (
    .a(\u2_Display/n4440 ),
    .b(1'b1),
    .c(\u2_Display/add136/c10 ),
    .o({\u2_Display/add136/c11 ,\u2_Display/n4453 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u11  (
    .a(\u2_Display/n4439 ),
    .b(1'b0),
    .c(\u2_Display/add136/c11 ),
    .o({\u2_Display/add136/c12 ,\u2_Display/n4453 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u12  (
    .a(\u2_Display/n4438 ),
    .b(1'b0),
    .c(\u2_Display/add136/c12 ),
    .o({\u2_Display/add136/c13 ,\u2_Display/n4453 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u13  (
    .a(\u2_Display/n4437 ),
    .b(1'b1),
    .c(\u2_Display/add136/c13 ),
    .o({\u2_Display/add136/c14 ,\u2_Display/n4453 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u14  (
    .a(\u2_Display/n4436 ),
    .b(1'b1),
    .c(\u2_Display/add136/c14 ),
    .o({\u2_Display/add136/c15 ,\u2_Display/n4453 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u15  (
    .a(\u2_Display/n4435 ),
    .b(1'b1),
    .c(\u2_Display/add136/c15 ),
    .o({\u2_Display/add136/c16 ,\u2_Display/n4453 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u16  (
    .a(\u2_Display/n4434 ),
    .b(1'b1),
    .c(\u2_Display/add136/c16 ),
    .o({\u2_Display/add136/c17 ,\u2_Display/n4453 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u17  (
    .a(\u2_Display/n4433 ),
    .b(1'b1),
    .c(\u2_Display/add136/c17 ),
    .o({\u2_Display/add136/c18 ,\u2_Display/n4453 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u18  (
    .a(\u2_Display/n4432 ),
    .b(1'b1),
    .c(\u2_Display/add136/c18 ),
    .o({\u2_Display/add136/c19 ,\u2_Display/n4453 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u19  (
    .a(\u2_Display/n4431 ),
    .b(1'b1),
    .c(\u2_Display/add136/c19 ),
    .o({\u2_Display/add136/c20 ,\u2_Display/n4453 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u2  (
    .a(\u2_Display/n4448 ),
    .b(1'b1),
    .c(\u2_Display/add136/c2 ),
    .o({\u2_Display/add136/c3 ,\u2_Display/n4453 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u20  (
    .a(\u2_Display/n4430 ),
    .b(1'b1),
    .c(\u2_Display/add136/c20 ),
    .o({\u2_Display/add136/c21 ,\u2_Display/n4453 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u21  (
    .a(\u2_Display/n4429 ),
    .b(1'b1),
    .c(\u2_Display/add136/c21 ),
    .o({\u2_Display/add136/c22 ,\u2_Display/n4453 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u22  (
    .a(\u2_Display/n4428 ),
    .b(1'b1),
    .c(\u2_Display/add136/c22 ),
    .o({\u2_Display/add136/c23 ,\u2_Display/n4453 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u23  (
    .a(\u2_Display/n4427 ),
    .b(1'b1),
    .c(\u2_Display/add136/c23 ),
    .o({\u2_Display/add136/c24 ,\u2_Display/n4453 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u24  (
    .a(\u2_Display/n4426 ),
    .b(1'b1),
    .c(\u2_Display/add136/c24 ),
    .o({\u2_Display/add136/c25 ,\u2_Display/n4453 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u25  (
    .a(\u2_Display/n4425 ),
    .b(1'b1),
    .c(\u2_Display/add136/c25 ),
    .o({\u2_Display/add136/c26 ,\u2_Display/n4453 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u26  (
    .a(\u2_Display/n4424 ),
    .b(1'b1),
    .c(\u2_Display/add136/c26 ),
    .o({\u2_Display/add136/c27 ,\u2_Display/n4453 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u27  (
    .a(\u2_Display/n4423 ),
    .b(1'b1),
    .c(\u2_Display/add136/c27 ),
    .o({\u2_Display/add136/c28 ,\u2_Display/n4453 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u28  (
    .a(\u2_Display/n4422 ),
    .b(1'b1),
    .c(\u2_Display/add136/c28 ),
    .o({\u2_Display/add136/c29 ,\u2_Display/n4453 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u29  (
    .a(\u2_Display/n4421 ),
    .b(1'b1),
    .c(\u2_Display/add136/c29 ),
    .o({\u2_Display/add136/c30 ,\u2_Display/n4453 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u3  (
    .a(\u2_Display/n4447 ),
    .b(1'b1),
    .c(\u2_Display/add136/c3 ),
    .o({\u2_Display/add136/c4 ,\u2_Display/n4453 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u30  (
    .a(\u2_Display/n4420 ),
    .b(1'b1),
    .c(\u2_Display/add136/c30 ),
    .o({\u2_Display/add136/c31 ,\u2_Display/n4453 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u31  (
    .a(\u2_Display/n4419 ),
    .b(1'b1),
    .c(\u2_Display/add136/c31 ),
    .o({open_n983,\u2_Display/n4453 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u4  (
    .a(\u2_Display/n4446 ),
    .b(1'b1),
    .c(\u2_Display/add136/c4 ),
    .o({\u2_Display/add136/c5 ,\u2_Display/n4453 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u5  (
    .a(\u2_Display/n4445 ),
    .b(1'b1),
    .c(\u2_Display/add136/c5 ),
    .o({\u2_Display/add136/c6 ,\u2_Display/n4453 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u6  (
    .a(\u2_Display/n4444 ),
    .b(1'b1),
    .c(\u2_Display/add136/c6 ),
    .o({\u2_Display/add136/c7 ,\u2_Display/n4453 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u7  (
    .a(\u2_Display/n4443 ),
    .b(1'b1),
    .c(\u2_Display/add136/c7 ),
    .o({\u2_Display/add136/c8 ,\u2_Display/n4453 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u8  (
    .a(\u2_Display/n4442 ),
    .b(1'b0),
    .c(\u2_Display/add136/c8 ),
    .o({\u2_Display/add136/c9 ,\u2_Display/n4453 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add136/u9  (
    .a(\u2_Display/n4441 ),
    .b(1'b1),
    .c(\u2_Display/add136/c9 ),
    .o({\u2_Display/add136/c10 ,\u2_Display/n4453 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add136/ucin  (
    .a(1'b1),
    .o({\u2_Display/add136/c0 ,open_n986}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u0  (
    .a(\u2_Display/n4485 ),
    .b(1'b1),
    .c(\u2_Display/add137/c0 ),
    .o({\u2_Display/add137/c1 ,\u2_Display/n4488 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u1  (
    .a(\u2_Display/n4484 ),
    .b(1'b1),
    .c(\u2_Display/add137/c1 ),
    .o({\u2_Display/add137/c2 ,\u2_Display/n4488 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u10  (
    .a(\u2_Display/n4475 ),
    .b(1'b0),
    .c(\u2_Display/add137/c10 ),
    .o({\u2_Display/add137/c11 ,\u2_Display/n4488 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u11  (
    .a(\u2_Display/n4474 ),
    .b(1'b0),
    .c(\u2_Display/add137/c11 ),
    .o({\u2_Display/add137/c12 ,\u2_Display/n4488 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u12  (
    .a(\u2_Display/n4473 ),
    .b(1'b1),
    .c(\u2_Display/add137/c12 ),
    .o({\u2_Display/add137/c13 ,\u2_Display/n4488 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u13  (
    .a(\u2_Display/n4472 ),
    .b(1'b1),
    .c(\u2_Display/add137/c13 ),
    .o({\u2_Display/add137/c14 ,\u2_Display/n4488 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u14  (
    .a(\u2_Display/n4471 ),
    .b(1'b1),
    .c(\u2_Display/add137/c14 ),
    .o({\u2_Display/add137/c15 ,\u2_Display/n4488 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u15  (
    .a(\u2_Display/n4470 ),
    .b(1'b1),
    .c(\u2_Display/add137/c15 ),
    .o({\u2_Display/add137/c16 ,\u2_Display/n4488 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u16  (
    .a(\u2_Display/n4469 ),
    .b(1'b1),
    .c(\u2_Display/add137/c16 ),
    .o({\u2_Display/add137/c17 ,\u2_Display/n4488 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u17  (
    .a(\u2_Display/n4468 ),
    .b(1'b1),
    .c(\u2_Display/add137/c17 ),
    .o({\u2_Display/add137/c18 ,\u2_Display/n4488 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u18  (
    .a(\u2_Display/n4467 ),
    .b(1'b1),
    .c(\u2_Display/add137/c18 ),
    .o({\u2_Display/add137/c19 ,\u2_Display/n4488 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u19  (
    .a(\u2_Display/n4466 ),
    .b(1'b1),
    .c(\u2_Display/add137/c19 ),
    .o({\u2_Display/add137/c20 ,\u2_Display/n4488 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u2  (
    .a(\u2_Display/n4483 ),
    .b(1'b1),
    .c(\u2_Display/add137/c2 ),
    .o({\u2_Display/add137/c3 ,\u2_Display/n4488 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u20  (
    .a(\u2_Display/n4465 ),
    .b(1'b1),
    .c(\u2_Display/add137/c20 ),
    .o({\u2_Display/add137/c21 ,\u2_Display/n4488 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u21  (
    .a(\u2_Display/n4464 ),
    .b(1'b1),
    .c(\u2_Display/add137/c21 ),
    .o({\u2_Display/add137/c22 ,\u2_Display/n4488 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u22  (
    .a(\u2_Display/n4463 ),
    .b(1'b1),
    .c(\u2_Display/add137/c22 ),
    .o({\u2_Display/add137/c23 ,\u2_Display/n4488 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u23  (
    .a(\u2_Display/n4462 ),
    .b(1'b1),
    .c(\u2_Display/add137/c23 ),
    .o({\u2_Display/add137/c24 ,\u2_Display/n4488 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u24  (
    .a(\u2_Display/n4461 ),
    .b(1'b1),
    .c(\u2_Display/add137/c24 ),
    .o({\u2_Display/add137/c25 ,\u2_Display/n4488 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u25  (
    .a(\u2_Display/n4460 ),
    .b(1'b1),
    .c(\u2_Display/add137/c25 ),
    .o({\u2_Display/add137/c26 ,\u2_Display/n4488 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u26  (
    .a(\u2_Display/n4459 ),
    .b(1'b1),
    .c(\u2_Display/add137/c26 ),
    .o({\u2_Display/add137/c27 ,\u2_Display/n4488 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u27  (
    .a(\u2_Display/n4458 ),
    .b(1'b1),
    .c(\u2_Display/add137/c27 ),
    .o({\u2_Display/add137/c28 ,\u2_Display/n4488 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u28  (
    .a(\u2_Display/n4457 ),
    .b(1'b1),
    .c(\u2_Display/add137/c28 ),
    .o({\u2_Display/add137/c29 ,\u2_Display/n4488 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u29  (
    .a(\u2_Display/n4456 ),
    .b(1'b1),
    .c(\u2_Display/add137/c29 ),
    .o({\u2_Display/add137/c30 ,\u2_Display/n4488 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u3  (
    .a(\u2_Display/n4482 ),
    .b(1'b1),
    .c(\u2_Display/add137/c3 ),
    .o({\u2_Display/add137/c4 ,\u2_Display/n4488 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u30  (
    .a(\u2_Display/n4455 ),
    .b(1'b1),
    .c(\u2_Display/add137/c30 ),
    .o({\u2_Display/add137/c31 ,\u2_Display/n4488 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u31  (
    .a(\u2_Display/n4454 ),
    .b(1'b1),
    .c(\u2_Display/add137/c31 ),
    .o({open_n987,\u2_Display/n4488 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u4  (
    .a(\u2_Display/n4481 ),
    .b(1'b1),
    .c(\u2_Display/add137/c4 ),
    .o({\u2_Display/add137/c5 ,\u2_Display/n4488 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u5  (
    .a(\u2_Display/n4480 ),
    .b(1'b1),
    .c(\u2_Display/add137/c5 ),
    .o({\u2_Display/add137/c6 ,\u2_Display/n4488 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u6  (
    .a(\u2_Display/n4479 ),
    .b(1'b1),
    .c(\u2_Display/add137/c6 ),
    .o({\u2_Display/add137/c7 ,\u2_Display/n4488 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u7  (
    .a(\u2_Display/n4478 ),
    .b(1'b0),
    .c(\u2_Display/add137/c7 ),
    .o({\u2_Display/add137/c8 ,\u2_Display/n4488 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u8  (
    .a(\u2_Display/n4477 ),
    .b(1'b1),
    .c(\u2_Display/add137/c8 ),
    .o({\u2_Display/add137/c9 ,\u2_Display/n4488 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add137/u9  (
    .a(\u2_Display/n4476 ),
    .b(1'b1),
    .c(\u2_Display/add137/c9 ),
    .o({\u2_Display/add137/c10 ,\u2_Display/n4488 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add137/ucin  (
    .a(1'b1),
    .o({\u2_Display/add137/c0 ,open_n990}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u0  (
    .a(\u2_Display/n4520 ),
    .b(1'b1),
    .c(\u2_Display/add138/c0 ),
    .o({\u2_Display/add138/c1 ,\u2_Display/n4523 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u1  (
    .a(\u2_Display/n4519 ),
    .b(1'b1),
    .c(\u2_Display/add138/c1 ),
    .o({\u2_Display/add138/c2 ,\u2_Display/n4523 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u10  (
    .a(\u2_Display/n4510 ),
    .b(1'b0),
    .c(\u2_Display/add138/c10 ),
    .o({\u2_Display/add138/c11 ,\u2_Display/n4523 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u11  (
    .a(\u2_Display/n4509 ),
    .b(1'b1),
    .c(\u2_Display/add138/c11 ),
    .o({\u2_Display/add138/c12 ,\u2_Display/n4523 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u12  (
    .a(\u2_Display/n4508 ),
    .b(1'b1),
    .c(\u2_Display/add138/c12 ),
    .o({\u2_Display/add138/c13 ,\u2_Display/n4523 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u13  (
    .a(\u2_Display/n4507 ),
    .b(1'b1),
    .c(\u2_Display/add138/c13 ),
    .o({\u2_Display/add138/c14 ,\u2_Display/n4523 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u14  (
    .a(\u2_Display/n4506 ),
    .b(1'b1),
    .c(\u2_Display/add138/c14 ),
    .o({\u2_Display/add138/c15 ,\u2_Display/n4523 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u15  (
    .a(\u2_Display/n4505 ),
    .b(1'b1),
    .c(\u2_Display/add138/c15 ),
    .o({\u2_Display/add138/c16 ,\u2_Display/n4523 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u16  (
    .a(\u2_Display/n4504 ),
    .b(1'b1),
    .c(\u2_Display/add138/c16 ),
    .o({\u2_Display/add138/c17 ,\u2_Display/n4523 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u17  (
    .a(\u2_Display/n4503 ),
    .b(1'b1),
    .c(\u2_Display/add138/c17 ),
    .o({\u2_Display/add138/c18 ,\u2_Display/n4523 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u18  (
    .a(\u2_Display/n4502 ),
    .b(1'b1),
    .c(\u2_Display/add138/c18 ),
    .o({\u2_Display/add138/c19 ,\u2_Display/n4523 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u19  (
    .a(\u2_Display/n4501 ),
    .b(1'b1),
    .c(\u2_Display/add138/c19 ),
    .o({\u2_Display/add138/c20 ,\u2_Display/n4523 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u2  (
    .a(\u2_Display/n4518 ),
    .b(1'b1),
    .c(\u2_Display/add138/c2 ),
    .o({\u2_Display/add138/c3 ,\u2_Display/n4523 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u20  (
    .a(\u2_Display/n4500 ),
    .b(1'b1),
    .c(\u2_Display/add138/c20 ),
    .o({\u2_Display/add138/c21 ,\u2_Display/n4523 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u21  (
    .a(\u2_Display/n4499 ),
    .b(1'b1),
    .c(\u2_Display/add138/c21 ),
    .o({\u2_Display/add138/c22 ,\u2_Display/n4523 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u22  (
    .a(\u2_Display/n4498 ),
    .b(1'b1),
    .c(\u2_Display/add138/c22 ),
    .o({\u2_Display/add138/c23 ,\u2_Display/n4523 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u23  (
    .a(\u2_Display/n4497 ),
    .b(1'b1),
    .c(\u2_Display/add138/c23 ),
    .o({\u2_Display/add138/c24 ,\u2_Display/n4523 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u24  (
    .a(\u2_Display/n4496 ),
    .b(1'b1),
    .c(\u2_Display/add138/c24 ),
    .o({\u2_Display/add138/c25 ,\u2_Display/n4523 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u25  (
    .a(\u2_Display/n4495 ),
    .b(1'b1),
    .c(\u2_Display/add138/c25 ),
    .o({\u2_Display/add138/c26 ,\u2_Display/n4523 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u26  (
    .a(\u2_Display/n4494 ),
    .b(1'b1),
    .c(\u2_Display/add138/c26 ),
    .o({\u2_Display/add138/c27 ,\u2_Display/n4523 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u27  (
    .a(\u2_Display/n4493 ),
    .b(1'b1),
    .c(\u2_Display/add138/c27 ),
    .o({\u2_Display/add138/c28 ,\u2_Display/n4523 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u28  (
    .a(\u2_Display/n4492 ),
    .b(1'b1),
    .c(\u2_Display/add138/c28 ),
    .o({\u2_Display/add138/c29 ,\u2_Display/n4523 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u29  (
    .a(\u2_Display/n4491 ),
    .b(1'b1),
    .c(\u2_Display/add138/c29 ),
    .o({\u2_Display/add138/c30 ,\u2_Display/n4523 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u3  (
    .a(\u2_Display/n4517 ),
    .b(1'b1),
    .c(\u2_Display/add138/c3 ),
    .o({\u2_Display/add138/c4 ,\u2_Display/n4523 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u30  (
    .a(\u2_Display/n4490 ),
    .b(1'b1),
    .c(\u2_Display/add138/c30 ),
    .o({\u2_Display/add138/c31 ,\u2_Display/n4523 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u31  (
    .a(\u2_Display/n4489 ),
    .b(1'b1),
    .c(\u2_Display/add138/c31 ),
    .o({open_n991,\u2_Display/n4523 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u4  (
    .a(\u2_Display/n4516 ),
    .b(1'b1),
    .c(\u2_Display/add138/c4 ),
    .o({\u2_Display/add138/c5 ,\u2_Display/n4523 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u5  (
    .a(\u2_Display/n4515 ),
    .b(1'b1),
    .c(\u2_Display/add138/c5 ),
    .o({\u2_Display/add138/c6 ,\u2_Display/n4523 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u6  (
    .a(\u2_Display/n4514 ),
    .b(1'b0),
    .c(\u2_Display/add138/c6 ),
    .o({\u2_Display/add138/c7 ,\u2_Display/n4523 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u7  (
    .a(\u2_Display/n4513 ),
    .b(1'b1),
    .c(\u2_Display/add138/c7 ),
    .o({\u2_Display/add138/c8 ,\u2_Display/n4523 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u8  (
    .a(\u2_Display/n4512 ),
    .b(1'b1),
    .c(\u2_Display/add138/c8 ),
    .o({\u2_Display/add138/c9 ,\u2_Display/n4523 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add138/u9  (
    .a(\u2_Display/n4511 ),
    .b(1'b0),
    .c(\u2_Display/add138/c9 ),
    .o({\u2_Display/add138/c10 ,\u2_Display/n4523 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add138/ucin  (
    .a(1'b1),
    .o({\u2_Display/add138/c0 ,open_n994}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add139/u0  (
    .a(\u2_Display/n4555 ),
    .b(1'b1),
    .c(\u2_Display/add139/c0 ),
    .o({\u2_Display/add139/c1 ,\u2_Display/n4558 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add139/u1  (
    .a(\u2_Display/n4554 ),
    .b(1'b1),
    .c(\u2_Display/add139/c1 ),
    .o({\u2_Display/add139/c2 ,\u2_Display/n4558 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add139/u2  (
    .a(\u2_Display/n4553 ),
    .b(1'b1),
    .c(\u2_Display/add139/c2 ),
    .o({\u2_Display/add139/c3 ,\u2_Display/n4558 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add139/u3  (
    .a(\u2_Display/n4552 ),
    .b(1'b1),
    .c(\u2_Display/add139/c3 ),
    .o({\u2_Display/add139/c4 ,\u2_Display/n4558 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add139/u4  (
    .a(\u2_Display/n4551 ),
    .b(1'b1),
    .c(\u2_Display/add139/c4 ),
    .o({\u2_Display/add139/c5 ,\u2_Display/n4558 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add139/u5  (
    .a(\u2_Display/n4550 ),
    .b(1'b0),
    .c(\u2_Display/add139/c5 ),
    .o({\u2_Display/add139/c6 ,\u2_Display/n4558 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add139/u6  (
    .a(\u2_Display/n4549 ),
    .b(1'b1),
    .c(\u2_Display/add139/c6 ),
    .o({\u2_Display/add139/c7 ,\u2_Display/n4558 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add139/u7  (
    .a(\u2_Display/n4548 ),
    .b(1'b1),
    .c(\u2_Display/add139/c7 ),
    .o({\u2_Display/add139/c8 ,\u2_Display/n4558 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add139/u8  (
    .a(\u2_Display/n4547 ),
    .b(1'b0),
    .c(\u2_Display/add139/c8 ),
    .o({\u2_Display/add139/c9 ,\u2_Display/n4558 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add139/u9  (
    .a(\u2_Display/n4546 ),
    .b(1'b0),
    .c(\u2_Display/add139/c9 ),
    .o({open_n995,\u2_Display/n4558 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add139/ucin  (
    .a(1'b1),
    .o({\u2_Display/add139/c0 ,open_n998}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u0  (
    .a(\u2_Display/counta [0]),
    .b(1'b1),
    .c(\u2_Display/add14/c0 ),
    .o({\u2_Display/add14/c1 ,\u2_Display/n4911 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u1  (
    .a(\u2_Display/counta [1]),
    .b(1'b1),
    .c(\u2_Display/add14/c1 ),
    .o({\u2_Display/add14/c2 ,\u2_Display/n4911 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u10  (
    .a(\u2_Display/counta [10]),
    .b(1'b1),
    .c(\u2_Display/add14/c10 ),
    .o({\u2_Display/add14/c11 ,\u2_Display/n4911 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u11  (
    .a(\u2_Display/counta [11]),
    .b(1'b1),
    .c(\u2_Display/add14/c11 ),
    .o({\u2_Display/add14/c12 ,\u2_Display/n4911 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u12  (
    .a(\u2_Display/counta [12]),
    .b(1'b1),
    .c(\u2_Display/add14/c12 ),
    .o({\u2_Display/add14/c13 ,\u2_Display/n4911 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u13  (
    .a(\u2_Display/counta [13]),
    .b(1'b1),
    .c(\u2_Display/add14/c13 ),
    .o({\u2_Display/add14/c14 ,\u2_Display/n4911 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u14  (
    .a(\u2_Display/counta [14]),
    .b(1'b1),
    .c(\u2_Display/add14/c14 ),
    .o({\u2_Display/add14/c15 ,\u2_Display/n4911 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u15  (
    .a(\u2_Display/counta [15]),
    .b(1'b1),
    .c(\u2_Display/add14/c15 ),
    .o({\u2_Display/add14/c16 ,\u2_Display/n4911 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u16  (
    .a(\u2_Display/counta [16]),
    .b(1'b1),
    .c(\u2_Display/add14/c16 ),
    .o({\u2_Display/add14/c17 ,\u2_Display/n4911 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u17  (
    .a(\u2_Display/counta [17]),
    .b(1'b1),
    .c(\u2_Display/add14/c17 ),
    .o({\u2_Display/add14/c18 ,\u2_Display/n4911 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u18  (
    .a(\u2_Display/counta [18]),
    .b(1'b1),
    .c(\u2_Display/add14/c18 ),
    .o({\u2_Display/add14/c19 ,\u2_Display/n4911 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u19  (
    .a(\u2_Display/counta [19]),
    .b(1'b1),
    .c(\u2_Display/add14/c19 ),
    .o({\u2_Display/add14/c20 ,\u2_Display/n4911 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u2  (
    .a(\u2_Display/counta [2]),
    .b(1'b1),
    .c(\u2_Display/add14/c2 ),
    .o({\u2_Display/add14/c3 ,\u2_Display/n4911 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u20  (
    .a(\u2_Display/counta [20]),
    .b(1'b1),
    .c(\u2_Display/add14/c20 ),
    .o({\u2_Display/add14/c21 ,\u2_Display/n4911 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u21  (
    .a(\u2_Display/counta [21]),
    .b(1'b1),
    .c(\u2_Display/add14/c21 ),
    .o({\u2_Display/add14/c22 ,\u2_Display/n4911 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u22  (
    .a(\u2_Display/counta [22]),
    .b(1'b1),
    .c(\u2_Display/add14/c22 ),
    .o({\u2_Display/add14/c23 ,\u2_Display/n4911 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u23  (
    .a(\u2_Display/counta [23]),
    .b(1'b1),
    .c(\u2_Display/add14/c23 ),
    .o({\u2_Display/add14/c24 ,\u2_Display/n4911 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u24  (
    .a(\u2_Display/counta [24]),
    .b(1'b1),
    .c(\u2_Display/add14/c24 ),
    .o({\u2_Display/add14/c25 ,\u2_Display/n4911 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u25  (
    .a(\u2_Display/counta [25]),
    .b(1'b1),
    .c(\u2_Display/add14/c25 ),
    .o({\u2_Display/add14/c26 ,\u2_Display/n4911 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u26  (
    .a(\u2_Display/counta [26]),
    .b(1'b1),
    .c(\u2_Display/add14/c26 ),
    .o({\u2_Display/add14/c27 ,\u2_Display/n4911 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u27  (
    .a(\u2_Display/counta [27]),
    .b(1'b1),
    .c(\u2_Display/add14/c27 ),
    .o({\u2_Display/add14/c28 ,\u2_Display/n4911 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u28  (
    .a(\u2_Display/counta [28]),
    .b(1'b1),
    .c(\u2_Display/add14/c28 ),
    .o({\u2_Display/add14/c29 ,\u2_Display/n4911 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u29  (
    .a(\u2_Display/counta [29]),
    .b(1'b0),
    .c(\u2_Display/add14/c29 ),
    .o({\u2_Display/add14/c30 ,\u2_Display/n4911 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u3  (
    .a(\u2_Display/counta [3]),
    .b(1'b1),
    .c(\u2_Display/add14/c3 ),
    .o({\u2_Display/add14/c4 ,\u2_Display/n4911 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u30  (
    .a(\u2_Display/counta [30]),
    .b(1'b1),
    .c(\u2_Display/add14/c30 ),
    .o({\u2_Display/add14/c31 ,\u2_Display/n4911 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u31  (
    .a(\u2_Display/counta [31]),
    .b(1'b0),
    .c(\u2_Display/add14/c31 ),
    .o({open_n999,\u2_Display/n4911 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u4  (
    .a(\u2_Display/counta [4]),
    .b(1'b1),
    .c(\u2_Display/add14/c4 ),
    .o({\u2_Display/add14/c5 ,\u2_Display/n4911 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u5  (
    .a(\u2_Display/counta [5]),
    .b(1'b1),
    .c(\u2_Display/add14/c5 ),
    .o({\u2_Display/add14/c6 ,\u2_Display/n4911 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u6  (
    .a(\u2_Display/counta [6]),
    .b(1'b1),
    .c(\u2_Display/add14/c6 ),
    .o({\u2_Display/add14/c7 ,\u2_Display/n4911 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u7  (
    .a(\u2_Display/counta [7]),
    .b(1'b1),
    .c(\u2_Display/add14/c7 ),
    .o({\u2_Display/add14/c8 ,\u2_Display/n4911 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u8  (
    .a(\u2_Display/counta [8]),
    .b(1'b1),
    .c(\u2_Display/add14/c8 ),
    .o({\u2_Display/add14/c9 ,\u2_Display/n4911 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add14/u9  (
    .a(\u2_Display/counta [9]),
    .b(1'b1),
    .c(\u2_Display/add14/c9 ),
    .o({\u2_Display/add14/c10 ,\u2_Display/n4911 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add14/ucin  (
    .a(1'b1),
    .o({\u2_Display/add14/c0 ,open_n1002}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u0  (
    .a(\u2_Display/n6101 ),
    .b(1'b1),
    .c(\u2_Display/add151/c0 ),
    .o({\u2_Display/add151/c1 ,\u2_Display/n4946 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u1  (
    .a(\u2_Display/n6100 ),
    .b(1'b1),
    .c(\u2_Display/add151/c1 ),
    .o({\u2_Display/add151/c2 ,\u2_Display/n4946 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u10  (
    .a(\u2_Display/n6091 ),
    .b(1'b1),
    .c(\u2_Display/add151/c10 ),
    .o({\u2_Display/add151/c11 ,\u2_Display/n4946 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u11  (
    .a(\u2_Display/n6090 ),
    .b(1'b1),
    .c(\u2_Display/add151/c11 ),
    .o({\u2_Display/add151/c12 ,\u2_Display/n4946 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u12  (
    .a(\u2_Display/n6089 ),
    .b(1'b1),
    .c(\u2_Display/add151/c12 ),
    .o({\u2_Display/add151/c13 ,\u2_Display/n4946 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u13  (
    .a(\u2_Display/n6088 ),
    .b(1'b1),
    .c(\u2_Display/add151/c13 ),
    .o({\u2_Display/add151/c14 ,\u2_Display/n4946 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u14  (
    .a(\u2_Display/n6087 ),
    .b(1'b1),
    .c(\u2_Display/add151/c14 ),
    .o({\u2_Display/add151/c15 ,\u2_Display/n4946 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u15  (
    .a(\u2_Display/n6086 ),
    .b(1'b1),
    .c(\u2_Display/add151/c15 ),
    .o({\u2_Display/add151/c16 ,\u2_Display/n4946 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u16  (
    .a(\u2_Display/n6085 ),
    .b(1'b1),
    .c(\u2_Display/add151/c16 ),
    .o({\u2_Display/add151/c17 ,\u2_Display/n4946 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u17  (
    .a(\u2_Display/n6084 ),
    .b(1'b1),
    .c(\u2_Display/add151/c17 ),
    .o({\u2_Display/add151/c18 ,\u2_Display/n4946 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u18  (
    .a(\u2_Display/n6083 ),
    .b(1'b1),
    .c(\u2_Display/add151/c18 ),
    .o({\u2_Display/add151/c19 ,\u2_Display/n4946 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u19  (
    .a(\u2_Display/n6082 ),
    .b(1'b1),
    .c(\u2_Display/add151/c19 ),
    .o({\u2_Display/add151/c20 ,\u2_Display/n4946 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u2  (
    .a(\u2_Display/n6099 ),
    .b(1'b1),
    .c(\u2_Display/add151/c2 ),
    .o({\u2_Display/add151/c3 ,\u2_Display/n4946 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u20  (
    .a(\u2_Display/n6081 ),
    .b(1'b1),
    .c(\u2_Display/add151/c20 ),
    .o({\u2_Display/add151/c21 ,\u2_Display/n4946 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u21  (
    .a(\u2_Display/n6080 ),
    .b(1'b1),
    .c(\u2_Display/add151/c21 ),
    .o({\u2_Display/add151/c22 ,\u2_Display/n4946 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u22  (
    .a(\u2_Display/n6079 ),
    .b(1'b1),
    .c(\u2_Display/add151/c22 ),
    .o({\u2_Display/add151/c23 ,\u2_Display/n4946 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u23  (
    .a(\u2_Display/n6078 ),
    .b(1'b1),
    .c(\u2_Display/add151/c23 ),
    .o({\u2_Display/add151/c24 ,\u2_Display/n4946 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u24  (
    .a(\u2_Display/n6077 ),
    .b(1'b1),
    .c(\u2_Display/add151/c24 ),
    .o({\u2_Display/add151/c25 ,\u2_Display/n4946 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u25  (
    .a(\u2_Display/n6076 ),
    .b(1'b1),
    .c(\u2_Display/add151/c25 ),
    .o({\u2_Display/add151/c26 ,\u2_Display/n4946 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u26  (
    .a(\u2_Display/n6075 ),
    .b(1'b1),
    .c(\u2_Display/add151/c26 ),
    .o({\u2_Display/add151/c27 ,\u2_Display/n4946 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u27  (
    .a(\u2_Display/n6074 ),
    .b(1'b1),
    .c(\u2_Display/add151/c27 ),
    .o({\u2_Display/add151/c28 ,\u2_Display/n4946 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u28  (
    .a(\u2_Display/n6073 ),
    .b(1'b0),
    .c(\u2_Display/add151/c28 ),
    .o({\u2_Display/add151/c29 ,\u2_Display/n4946 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u29  (
    .a(\u2_Display/n6072 ),
    .b(1'b1),
    .c(\u2_Display/add151/c29 ),
    .o({\u2_Display/add151/c30 ,\u2_Display/n4946 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u3  (
    .a(\u2_Display/n6098 ),
    .b(1'b1),
    .c(\u2_Display/add151/c3 ),
    .o({\u2_Display/add151/c4 ,\u2_Display/n4946 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u30  (
    .a(\u2_Display/n6071 ),
    .b(1'b0),
    .c(\u2_Display/add151/c30 ),
    .o({\u2_Display/add151/c31 ,\u2_Display/n4946 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u31  (
    .a(\u2_Display/n6070 ),
    .b(1'b1),
    .c(\u2_Display/add151/c31 ),
    .o({open_n1003,\u2_Display/n4946 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u4  (
    .a(\u2_Display/n6097 ),
    .b(1'b1),
    .c(\u2_Display/add151/c4 ),
    .o({\u2_Display/add151/c5 ,\u2_Display/n4946 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u5  (
    .a(\u2_Display/n6096 ),
    .b(1'b1),
    .c(\u2_Display/add151/c5 ),
    .o({\u2_Display/add151/c6 ,\u2_Display/n4946 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u6  (
    .a(\u2_Display/n6095 ),
    .b(1'b1),
    .c(\u2_Display/add151/c6 ),
    .o({\u2_Display/add151/c7 ,\u2_Display/n4946 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u7  (
    .a(\u2_Display/n6094 ),
    .b(1'b1),
    .c(\u2_Display/add151/c7 ),
    .o({\u2_Display/add151/c8 ,\u2_Display/n4946 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u8  (
    .a(\u2_Display/n6093 ),
    .b(1'b1),
    .c(\u2_Display/add151/c8 ),
    .o({\u2_Display/add151/c9 ,\u2_Display/n4946 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add151/u9  (
    .a(\u2_Display/n6092 ),
    .b(1'b1),
    .c(\u2_Display/add151/c9 ),
    .o({\u2_Display/add151/c10 ,\u2_Display/n4946 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add151/ucin  (
    .a(1'b1),
    .o({\u2_Display/add151/c0 ,open_n1006}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u0  (
    .a(\u2_Display/n6136 ),
    .b(1'b1),
    .c(\u2_Display/add152/c0 ),
    .o({\u2_Display/add152/c1 ,\u2_Display/n4981 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u1  (
    .a(\u2_Display/n6135 ),
    .b(1'b1),
    .c(\u2_Display/add152/c1 ),
    .o({\u2_Display/add152/c2 ,\u2_Display/n4981 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u10  (
    .a(\u2_Display/n6126 ),
    .b(1'b1),
    .c(\u2_Display/add152/c10 ),
    .o({\u2_Display/add152/c11 ,\u2_Display/n4981 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u11  (
    .a(\u2_Display/n6125 ),
    .b(1'b1),
    .c(\u2_Display/add152/c11 ),
    .o({\u2_Display/add152/c12 ,\u2_Display/n4981 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u12  (
    .a(\u2_Display/n6124 ),
    .b(1'b1),
    .c(\u2_Display/add152/c12 ),
    .o({\u2_Display/add152/c13 ,\u2_Display/n4981 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u13  (
    .a(\u2_Display/n6123 ),
    .b(1'b1),
    .c(\u2_Display/add152/c13 ),
    .o({\u2_Display/add152/c14 ,\u2_Display/n4981 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u14  (
    .a(\u2_Display/n6122 ),
    .b(1'b1),
    .c(\u2_Display/add152/c14 ),
    .o({\u2_Display/add152/c15 ,\u2_Display/n4981 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u15  (
    .a(\u2_Display/n6121 ),
    .b(1'b1),
    .c(\u2_Display/add152/c15 ),
    .o({\u2_Display/add152/c16 ,\u2_Display/n4981 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u16  (
    .a(\u2_Display/n6120 ),
    .b(1'b1),
    .c(\u2_Display/add152/c16 ),
    .o({\u2_Display/add152/c17 ,\u2_Display/n4981 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u17  (
    .a(\u2_Display/n6119 ),
    .b(1'b1),
    .c(\u2_Display/add152/c17 ),
    .o({\u2_Display/add152/c18 ,\u2_Display/n4981 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u18  (
    .a(\u2_Display/n6118 ),
    .b(1'b1),
    .c(\u2_Display/add152/c18 ),
    .o({\u2_Display/add152/c19 ,\u2_Display/n4981 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u19  (
    .a(\u2_Display/n6117 ),
    .b(1'b1),
    .c(\u2_Display/add152/c19 ),
    .o({\u2_Display/add152/c20 ,\u2_Display/n4981 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u2  (
    .a(\u2_Display/n6134 ),
    .b(1'b1),
    .c(\u2_Display/add152/c2 ),
    .o({\u2_Display/add152/c3 ,\u2_Display/n4981 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u20  (
    .a(\u2_Display/n6116 ),
    .b(1'b1),
    .c(\u2_Display/add152/c20 ),
    .o({\u2_Display/add152/c21 ,\u2_Display/n4981 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u21  (
    .a(\u2_Display/n6115 ),
    .b(1'b1),
    .c(\u2_Display/add152/c21 ),
    .o({\u2_Display/add152/c22 ,\u2_Display/n4981 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u22  (
    .a(\u2_Display/n6114 ),
    .b(1'b1),
    .c(\u2_Display/add152/c22 ),
    .o({\u2_Display/add152/c23 ,\u2_Display/n4981 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u23  (
    .a(\u2_Display/n6113 ),
    .b(1'b1),
    .c(\u2_Display/add152/c23 ),
    .o({\u2_Display/add152/c24 ,\u2_Display/n4981 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u24  (
    .a(\u2_Display/n6112 ),
    .b(1'b1),
    .c(\u2_Display/add152/c24 ),
    .o({\u2_Display/add152/c25 ,\u2_Display/n4981 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u25  (
    .a(\u2_Display/n6111 ),
    .b(1'b1),
    .c(\u2_Display/add152/c25 ),
    .o({\u2_Display/add152/c26 ,\u2_Display/n4981 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u26  (
    .a(\u2_Display/n6110 ),
    .b(1'b1),
    .c(\u2_Display/add152/c26 ),
    .o({\u2_Display/add152/c27 ,\u2_Display/n4981 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u27  (
    .a(\u2_Display/n6109 ),
    .b(1'b0),
    .c(\u2_Display/add152/c27 ),
    .o({\u2_Display/add152/c28 ,\u2_Display/n4981 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u28  (
    .a(\u2_Display/n6108 ),
    .b(1'b1),
    .c(\u2_Display/add152/c28 ),
    .o({\u2_Display/add152/c29 ,\u2_Display/n4981 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u29  (
    .a(\u2_Display/n6107 ),
    .b(1'b0),
    .c(\u2_Display/add152/c29 ),
    .o({\u2_Display/add152/c30 ,\u2_Display/n4981 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u3  (
    .a(\u2_Display/n6133 ),
    .b(1'b1),
    .c(\u2_Display/add152/c3 ),
    .o({\u2_Display/add152/c4 ,\u2_Display/n4981 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u30  (
    .a(\u2_Display/n6106 ),
    .b(1'b1),
    .c(\u2_Display/add152/c30 ),
    .o({\u2_Display/add152/c31 ,\u2_Display/n4981 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u31  (
    .a(\u2_Display/n6105 ),
    .b(1'b1),
    .c(\u2_Display/add152/c31 ),
    .o({open_n1007,\u2_Display/n4981 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u4  (
    .a(\u2_Display/n6132 ),
    .b(1'b1),
    .c(\u2_Display/add152/c4 ),
    .o({\u2_Display/add152/c5 ,\u2_Display/n4981 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u5  (
    .a(\u2_Display/n6131 ),
    .b(1'b1),
    .c(\u2_Display/add152/c5 ),
    .o({\u2_Display/add152/c6 ,\u2_Display/n4981 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u6  (
    .a(\u2_Display/n6130 ),
    .b(1'b1),
    .c(\u2_Display/add152/c6 ),
    .o({\u2_Display/add152/c7 ,\u2_Display/n4981 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u7  (
    .a(\u2_Display/n6129 ),
    .b(1'b1),
    .c(\u2_Display/add152/c7 ),
    .o({\u2_Display/add152/c8 ,\u2_Display/n4981 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u8  (
    .a(\u2_Display/n6128 ),
    .b(1'b1),
    .c(\u2_Display/add152/c8 ),
    .o({\u2_Display/add152/c9 ,\u2_Display/n4981 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add152/u9  (
    .a(\u2_Display/n6127 ),
    .b(1'b1),
    .c(\u2_Display/add152/c9 ),
    .o({\u2_Display/add152/c10 ,\u2_Display/n4981 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add152/ucin  (
    .a(1'b1),
    .o({\u2_Display/add152/c0 ,open_n1010}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u0  (
    .a(\u2_Display/n6171 ),
    .b(1'b1),
    .c(\u2_Display/add153/c0 ),
    .o({\u2_Display/add153/c1 ,\u2_Display/n5016 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u1  (
    .a(\u2_Display/n6170 ),
    .b(1'b1),
    .c(\u2_Display/add153/c1 ),
    .o({\u2_Display/add153/c2 ,\u2_Display/n5016 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u10  (
    .a(\u2_Display/n6161 ),
    .b(1'b1),
    .c(\u2_Display/add153/c10 ),
    .o({\u2_Display/add153/c11 ,\u2_Display/n5016 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u11  (
    .a(\u2_Display/n6160 ),
    .b(1'b1),
    .c(\u2_Display/add153/c11 ),
    .o({\u2_Display/add153/c12 ,\u2_Display/n5016 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u12  (
    .a(\u2_Display/n6159 ),
    .b(1'b1),
    .c(\u2_Display/add153/c12 ),
    .o({\u2_Display/add153/c13 ,\u2_Display/n5016 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u13  (
    .a(\u2_Display/n6158 ),
    .b(1'b1),
    .c(\u2_Display/add153/c13 ),
    .o({\u2_Display/add153/c14 ,\u2_Display/n5016 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u14  (
    .a(\u2_Display/n6157 ),
    .b(1'b1),
    .c(\u2_Display/add153/c14 ),
    .o({\u2_Display/add153/c15 ,\u2_Display/n5016 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u15  (
    .a(\u2_Display/n6156 ),
    .b(1'b1),
    .c(\u2_Display/add153/c15 ),
    .o({\u2_Display/add153/c16 ,\u2_Display/n5016 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u16  (
    .a(\u2_Display/n6155 ),
    .b(1'b1),
    .c(\u2_Display/add153/c16 ),
    .o({\u2_Display/add153/c17 ,\u2_Display/n5016 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u17  (
    .a(\u2_Display/n6154 ),
    .b(1'b1),
    .c(\u2_Display/add153/c17 ),
    .o({\u2_Display/add153/c18 ,\u2_Display/n5016 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u18  (
    .a(\u2_Display/n6153 ),
    .b(1'b1),
    .c(\u2_Display/add153/c18 ),
    .o({\u2_Display/add153/c19 ,\u2_Display/n5016 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u19  (
    .a(\u2_Display/n6152 ),
    .b(1'b1),
    .c(\u2_Display/add153/c19 ),
    .o({\u2_Display/add153/c20 ,\u2_Display/n5016 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u2  (
    .a(\u2_Display/n6169 ),
    .b(1'b1),
    .c(\u2_Display/add153/c2 ),
    .o({\u2_Display/add153/c3 ,\u2_Display/n5016 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u20  (
    .a(\u2_Display/n6151 ),
    .b(1'b1),
    .c(\u2_Display/add153/c20 ),
    .o({\u2_Display/add153/c21 ,\u2_Display/n5016 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u21  (
    .a(\u2_Display/n6150 ),
    .b(1'b1),
    .c(\u2_Display/add153/c21 ),
    .o({\u2_Display/add153/c22 ,\u2_Display/n5016 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u22  (
    .a(\u2_Display/n6149 ),
    .b(1'b1),
    .c(\u2_Display/add153/c22 ),
    .o({\u2_Display/add153/c23 ,\u2_Display/n5016 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u23  (
    .a(\u2_Display/n6148 ),
    .b(1'b1),
    .c(\u2_Display/add153/c23 ),
    .o({\u2_Display/add153/c24 ,\u2_Display/n5016 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u24  (
    .a(\u2_Display/n6147 ),
    .b(1'b1),
    .c(\u2_Display/add153/c24 ),
    .o({\u2_Display/add153/c25 ,\u2_Display/n5016 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u25  (
    .a(\u2_Display/n6146 ),
    .b(1'b1),
    .c(\u2_Display/add153/c25 ),
    .o({\u2_Display/add153/c26 ,\u2_Display/n5016 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u26  (
    .a(\u2_Display/n6145 ),
    .b(1'b0),
    .c(\u2_Display/add153/c26 ),
    .o({\u2_Display/add153/c27 ,\u2_Display/n5016 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u27  (
    .a(\u2_Display/n6144 ),
    .b(1'b1),
    .c(\u2_Display/add153/c27 ),
    .o({\u2_Display/add153/c28 ,\u2_Display/n5016 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u28  (
    .a(\u2_Display/n6143 ),
    .b(1'b0),
    .c(\u2_Display/add153/c28 ),
    .o({\u2_Display/add153/c29 ,\u2_Display/n5016 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u29  (
    .a(\u2_Display/n6142 ),
    .b(1'b1),
    .c(\u2_Display/add153/c29 ),
    .o({\u2_Display/add153/c30 ,\u2_Display/n5016 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u3  (
    .a(\u2_Display/n6168 ),
    .b(1'b1),
    .c(\u2_Display/add153/c3 ),
    .o({\u2_Display/add153/c4 ,\u2_Display/n5016 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u30  (
    .a(\u2_Display/n6141 ),
    .b(1'b1),
    .c(\u2_Display/add153/c30 ),
    .o({\u2_Display/add153/c31 ,\u2_Display/n5016 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u31  (
    .a(\u2_Display/n6140 ),
    .b(1'b1),
    .c(\u2_Display/add153/c31 ),
    .o({open_n1011,\u2_Display/n5016 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u4  (
    .a(\u2_Display/n6167 ),
    .b(1'b1),
    .c(\u2_Display/add153/c4 ),
    .o({\u2_Display/add153/c5 ,\u2_Display/n5016 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u5  (
    .a(\u2_Display/n6166 ),
    .b(1'b1),
    .c(\u2_Display/add153/c5 ),
    .o({\u2_Display/add153/c6 ,\u2_Display/n5016 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u6  (
    .a(\u2_Display/n6165 ),
    .b(1'b1),
    .c(\u2_Display/add153/c6 ),
    .o({\u2_Display/add153/c7 ,\u2_Display/n5016 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u7  (
    .a(\u2_Display/n6164 ),
    .b(1'b1),
    .c(\u2_Display/add153/c7 ),
    .o({\u2_Display/add153/c8 ,\u2_Display/n5016 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u8  (
    .a(\u2_Display/n6163 ),
    .b(1'b1),
    .c(\u2_Display/add153/c8 ),
    .o({\u2_Display/add153/c9 ,\u2_Display/n5016 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add153/u9  (
    .a(\u2_Display/n6162 ),
    .b(1'b1),
    .c(\u2_Display/add153/c9 ),
    .o({\u2_Display/add153/c10 ,\u2_Display/n5016 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add153/ucin  (
    .a(1'b1),
    .o({\u2_Display/add153/c0 ,open_n1014}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u0  (
    .a(\u2_Display/n6206 ),
    .b(1'b1),
    .c(\u2_Display/add154/c0 ),
    .o({\u2_Display/add154/c1 ,\u2_Display/n5051 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u1  (
    .a(\u2_Display/n6205 ),
    .b(1'b1),
    .c(\u2_Display/add154/c1 ),
    .o({\u2_Display/add154/c2 ,\u2_Display/n5051 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u10  (
    .a(\u2_Display/n6196 ),
    .b(1'b1),
    .c(\u2_Display/add154/c10 ),
    .o({\u2_Display/add154/c11 ,\u2_Display/n5051 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u11  (
    .a(\u2_Display/n6195 ),
    .b(1'b1),
    .c(\u2_Display/add154/c11 ),
    .o({\u2_Display/add154/c12 ,\u2_Display/n5051 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u12  (
    .a(\u2_Display/n6194 ),
    .b(1'b1),
    .c(\u2_Display/add154/c12 ),
    .o({\u2_Display/add154/c13 ,\u2_Display/n5051 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u13  (
    .a(\u2_Display/n6193 ),
    .b(1'b1),
    .c(\u2_Display/add154/c13 ),
    .o({\u2_Display/add154/c14 ,\u2_Display/n5051 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u14  (
    .a(\u2_Display/n6192 ),
    .b(1'b1),
    .c(\u2_Display/add154/c14 ),
    .o({\u2_Display/add154/c15 ,\u2_Display/n5051 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u15  (
    .a(\u2_Display/n6191 ),
    .b(1'b1),
    .c(\u2_Display/add154/c15 ),
    .o({\u2_Display/add154/c16 ,\u2_Display/n5051 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u16  (
    .a(\u2_Display/n6190 ),
    .b(1'b1),
    .c(\u2_Display/add154/c16 ),
    .o({\u2_Display/add154/c17 ,\u2_Display/n5051 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u17  (
    .a(\u2_Display/n6189 ),
    .b(1'b1),
    .c(\u2_Display/add154/c17 ),
    .o({\u2_Display/add154/c18 ,\u2_Display/n5051 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u18  (
    .a(\u2_Display/n6188 ),
    .b(1'b1),
    .c(\u2_Display/add154/c18 ),
    .o({\u2_Display/add154/c19 ,\u2_Display/n5051 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u19  (
    .a(\u2_Display/n6187 ),
    .b(1'b1),
    .c(\u2_Display/add154/c19 ),
    .o({\u2_Display/add154/c20 ,\u2_Display/n5051 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u2  (
    .a(\u2_Display/n6204 ),
    .b(1'b1),
    .c(\u2_Display/add154/c2 ),
    .o({\u2_Display/add154/c3 ,\u2_Display/n5051 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u20  (
    .a(\u2_Display/n6186 ),
    .b(1'b1),
    .c(\u2_Display/add154/c20 ),
    .o({\u2_Display/add154/c21 ,\u2_Display/n5051 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u21  (
    .a(\u2_Display/n6185 ),
    .b(1'b1),
    .c(\u2_Display/add154/c21 ),
    .o({\u2_Display/add154/c22 ,\u2_Display/n5051 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u22  (
    .a(\u2_Display/n6184 ),
    .b(1'b1),
    .c(\u2_Display/add154/c22 ),
    .o({\u2_Display/add154/c23 ,\u2_Display/n5051 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u23  (
    .a(\u2_Display/n6183 ),
    .b(1'b1),
    .c(\u2_Display/add154/c23 ),
    .o({\u2_Display/add154/c24 ,\u2_Display/n5051 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u24  (
    .a(\u2_Display/n6182 ),
    .b(1'b1),
    .c(\u2_Display/add154/c24 ),
    .o({\u2_Display/add154/c25 ,\u2_Display/n5051 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u25  (
    .a(\u2_Display/n6181 ),
    .b(1'b0),
    .c(\u2_Display/add154/c25 ),
    .o({\u2_Display/add154/c26 ,\u2_Display/n5051 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u26  (
    .a(\u2_Display/n6180 ),
    .b(1'b1),
    .c(\u2_Display/add154/c26 ),
    .o({\u2_Display/add154/c27 ,\u2_Display/n5051 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u27  (
    .a(\u2_Display/n6179 ),
    .b(1'b0),
    .c(\u2_Display/add154/c27 ),
    .o({\u2_Display/add154/c28 ,\u2_Display/n5051 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u28  (
    .a(\u2_Display/n6178 ),
    .b(1'b1),
    .c(\u2_Display/add154/c28 ),
    .o({\u2_Display/add154/c29 ,\u2_Display/n5051 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u29  (
    .a(\u2_Display/n6177 ),
    .b(1'b1),
    .c(\u2_Display/add154/c29 ),
    .o({\u2_Display/add154/c30 ,\u2_Display/n5051 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u3  (
    .a(\u2_Display/n6203 ),
    .b(1'b1),
    .c(\u2_Display/add154/c3 ),
    .o({\u2_Display/add154/c4 ,\u2_Display/n5051 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u30  (
    .a(\u2_Display/n6176 ),
    .b(1'b1),
    .c(\u2_Display/add154/c30 ),
    .o({\u2_Display/add154/c31 ,\u2_Display/n5051 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u31  (
    .a(\u2_Display/n6175 ),
    .b(1'b1),
    .c(\u2_Display/add154/c31 ),
    .o({open_n1015,\u2_Display/n5051 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u4  (
    .a(\u2_Display/n6202 ),
    .b(1'b1),
    .c(\u2_Display/add154/c4 ),
    .o({\u2_Display/add154/c5 ,\u2_Display/n5051 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u5  (
    .a(\u2_Display/n6201 ),
    .b(1'b1),
    .c(\u2_Display/add154/c5 ),
    .o({\u2_Display/add154/c6 ,\u2_Display/n5051 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u6  (
    .a(\u2_Display/n6200 ),
    .b(1'b1),
    .c(\u2_Display/add154/c6 ),
    .o({\u2_Display/add154/c7 ,\u2_Display/n5051 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u7  (
    .a(\u2_Display/n6199 ),
    .b(1'b1),
    .c(\u2_Display/add154/c7 ),
    .o({\u2_Display/add154/c8 ,\u2_Display/n5051 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u8  (
    .a(\u2_Display/n6198 ),
    .b(1'b1),
    .c(\u2_Display/add154/c8 ),
    .o({\u2_Display/add154/c9 ,\u2_Display/n5051 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add154/u9  (
    .a(\u2_Display/n6197 ),
    .b(1'b1),
    .c(\u2_Display/add154/c9 ),
    .o({\u2_Display/add154/c10 ,\u2_Display/n5051 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add154/ucin  (
    .a(1'b1),
    .o({\u2_Display/add154/c0 ,open_n1018}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u0  (
    .a(\u2_Display/n6241 ),
    .b(1'b1),
    .c(\u2_Display/add155/c0 ),
    .o({\u2_Display/add155/c1 ,\u2_Display/n5086 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u1  (
    .a(\u2_Display/n6240 ),
    .b(1'b1),
    .c(\u2_Display/add155/c1 ),
    .o({\u2_Display/add155/c2 ,\u2_Display/n5086 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u10  (
    .a(\u2_Display/n6231 ),
    .b(1'b1),
    .c(\u2_Display/add155/c10 ),
    .o({\u2_Display/add155/c11 ,\u2_Display/n5086 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u11  (
    .a(\u2_Display/n6230 ),
    .b(1'b1),
    .c(\u2_Display/add155/c11 ),
    .o({\u2_Display/add155/c12 ,\u2_Display/n5086 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u12  (
    .a(\u2_Display/n6229 ),
    .b(1'b1),
    .c(\u2_Display/add155/c12 ),
    .o({\u2_Display/add155/c13 ,\u2_Display/n5086 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u13  (
    .a(\u2_Display/n6228 ),
    .b(1'b1),
    .c(\u2_Display/add155/c13 ),
    .o({\u2_Display/add155/c14 ,\u2_Display/n5086 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u14  (
    .a(\u2_Display/n6227 ),
    .b(1'b1),
    .c(\u2_Display/add155/c14 ),
    .o({\u2_Display/add155/c15 ,\u2_Display/n5086 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u15  (
    .a(\u2_Display/n6226 ),
    .b(1'b1),
    .c(\u2_Display/add155/c15 ),
    .o({\u2_Display/add155/c16 ,\u2_Display/n5086 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u16  (
    .a(\u2_Display/n6225 ),
    .b(1'b1),
    .c(\u2_Display/add155/c16 ),
    .o({\u2_Display/add155/c17 ,\u2_Display/n5086 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u17  (
    .a(\u2_Display/n6224 ),
    .b(1'b1),
    .c(\u2_Display/add155/c17 ),
    .o({\u2_Display/add155/c18 ,\u2_Display/n5086 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u18  (
    .a(\u2_Display/n6223 ),
    .b(1'b1),
    .c(\u2_Display/add155/c18 ),
    .o({\u2_Display/add155/c19 ,\u2_Display/n5086 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u19  (
    .a(\u2_Display/n6222 ),
    .b(1'b1),
    .c(\u2_Display/add155/c19 ),
    .o({\u2_Display/add155/c20 ,\u2_Display/n5086 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u2  (
    .a(\u2_Display/n6239 ),
    .b(1'b1),
    .c(\u2_Display/add155/c2 ),
    .o({\u2_Display/add155/c3 ,\u2_Display/n5086 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u20  (
    .a(\u2_Display/n6221 ),
    .b(1'b1),
    .c(\u2_Display/add155/c20 ),
    .o({\u2_Display/add155/c21 ,\u2_Display/n5086 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u21  (
    .a(\u2_Display/n6220 ),
    .b(1'b1),
    .c(\u2_Display/add155/c21 ),
    .o({\u2_Display/add155/c22 ,\u2_Display/n5086 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u22  (
    .a(\u2_Display/n6219 ),
    .b(1'b1),
    .c(\u2_Display/add155/c22 ),
    .o({\u2_Display/add155/c23 ,\u2_Display/n5086 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u23  (
    .a(\u2_Display/n6218 ),
    .b(1'b1),
    .c(\u2_Display/add155/c23 ),
    .o({\u2_Display/add155/c24 ,\u2_Display/n5086 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u24  (
    .a(\u2_Display/n6217 ),
    .b(1'b0),
    .c(\u2_Display/add155/c24 ),
    .o({\u2_Display/add155/c25 ,\u2_Display/n5086 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u25  (
    .a(\u2_Display/n6216 ),
    .b(1'b1),
    .c(\u2_Display/add155/c25 ),
    .o({\u2_Display/add155/c26 ,\u2_Display/n5086 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u26  (
    .a(\u2_Display/n6215 ),
    .b(1'b0),
    .c(\u2_Display/add155/c26 ),
    .o({\u2_Display/add155/c27 ,\u2_Display/n5086 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u27  (
    .a(\u2_Display/n6214 ),
    .b(1'b1),
    .c(\u2_Display/add155/c27 ),
    .o({\u2_Display/add155/c28 ,\u2_Display/n5086 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u28  (
    .a(\u2_Display/n6213 ),
    .b(1'b1),
    .c(\u2_Display/add155/c28 ),
    .o({\u2_Display/add155/c29 ,\u2_Display/n5086 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u29  (
    .a(\u2_Display/n6212 ),
    .b(1'b1),
    .c(\u2_Display/add155/c29 ),
    .o({\u2_Display/add155/c30 ,\u2_Display/n5086 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u3  (
    .a(\u2_Display/n6238 ),
    .b(1'b1),
    .c(\u2_Display/add155/c3 ),
    .o({\u2_Display/add155/c4 ,\u2_Display/n5086 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u30  (
    .a(\u2_Display/n6211 ),
    .b(1'b1),
    .c(\u2_Display/add155/c30 ),
    .o({\u2_Display/add155/c31 ,\u2_Display/n5086 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u31  (
    .a(\u2_Display/n6210 ),
    .b(1'b1),
    .c(\u2_Display/add155/c31 ),
    .o({open_n1019,\u2_Display/n5086 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u4  (
    .a(\u2_Display/n6237 ),
    .b(1'b1),
    .c(\u2_Display/add155/c4 ),
    .o({\u2_Display/add155/c5 ,\u2_Display/n5086 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u5  (
    .a(\u2_Display/n6236 ),
    .b(1'b1),
    .c(\u2_Display/add155/c5 ),
    .o({\u2_Display/add155/c6 ,\u2_Display/n5086 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u6  (
    .a(\u2_Display/n6235 ),
    .b(1'b1),
    .c(\u2_Display/add155/c6 ),
    .o({\u2_Display/add155/c7 ,\u2_Display/n5086 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u7  (
    .a(\u2_Display/n6234 ),
    .b(1'b1),
    .c(\u2_Display/add155/c7 ),
    .o({\u2_Display/add155/c8 ,\u2_Display/n5086 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u8  (
    .a(\u2_Display/n6233 ),
    .b(1'b1),
    .c(\u2_Display/add155/c8 ),
    .o({\u2_Display/add155/c9 ,\u2_Display/n5086 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add155/u9  (
    .a(\u2_Display/n6232 ),
    .b(1'b1),
    .c(\u2_Display/add155/c9 ),
    .o({\u2_Display/add155/c10 ,\u2_Display/n5086 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add155/ucin  (
    .a(1'b1),
    .o({\u2_Display/add155/c0 ,open_n1022}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u0  (
    .a(\u2_Display/n6276 ),
    .b(1'b1),
    .c(\u2_Display/add156/c0 ),
    .o({\u2_Display/add156/c1 ,\u2_Display/n5121 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u1  (
    .a(\u2_Display/n6275 ),
    .b(1'b1),
    .c(\u2_Display/add156/c1 ),
    .o({\u2_Display/add156/c2 ,\u2_Display/n5121 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u10  (
    .a(\u2_Display/n6266 ),
    .b(1'b1),
    .c(\u2_Display/add156/c10 ),
    .o({\u2_Display/add156/c11 ,\u2_Display/n5121 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u11  (
    .a(\u2_Display/n6265 ),
    .b(1'b1),
    .c(\u2_Display/add156/c11 ),
    .o({\u2_Display/add156/c12 ,\u2_Display/n5121 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u12  (
    .a(\u2_Display/n6264 ),
    .b(1'b1),
    .c(\u2_Display/add156/c12 ),
    .o({\u2_Display/add156/c13 ,\u2_Display/n5121 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u13  (
    .a(\u2_Display/n6263 ),
    .b(1'b1),
    .c(\u2_Display/add156/c13 ),
    .o({\u2_Display/add156/c14 ,\u2_Display/n5121 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u14  (
    .a(\u2_Display/n6262 ),
    .b(1'b1),
    .c(\u2_Display/add156/c14 ),
    .o({\u2_Display/add156/c15 ,\u2_Display/n5121 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u15  (
    .a(\u2_Display/n6261 ),
    .b(1'b1),
    .c(\u2_Display/add156/c15 ),
    .o({\u2_Display/add156/c16 ,\u2_Display/n5121 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u16  (
    .a(\u2_Display/n6260 ),
    .b(1'b1),
    .c(\u2_Display/add156/c16 ),
    .o({\u2_Display/add156/c17 ,\u2_Display/n5121 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u17  (
    .a(\u2_Display/n6259 ),
    .b(1'b1),
    .c(\u2_Display/add156/c17 ),
    .o({\u2_Display/add156/c18 ,\u2_Display/n5121 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u18  (
    .a(\u2_Display/n6258 ),
    .b(1'b1),
    .c(\u2_Display/add156/c18 ),
    .o({\u2_Display/add156/c19 ,\u2_Display/n5121 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u19  (
    .a(\u2_Display/n6257 ),
    .b(1'b1),
    .c(\u2_Display/add156/c19 ),
    .o({\u2_Display/add156/c20 ,\u2_Display/n5121 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u2  (
    .a(\u2_Display/n6274 ),
    .b(1'b1),
    .c(\u2_Display/add156/c2 ),
    .o({\u2_Display/add156/c3 ,\u2_Display/n5121 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u20  (
    .a(\u2_Display/n6256 ),
    .b(1'b1),
    .c(\u2_Display/add156/c20 ),
    .o({\u2_Display/add156/c21 ,\u2_Display/n5121 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u21  (
    .a(\u2_Display/n6255 ),
    .b(1'b1),
    .c(\u2_Display/add156/c21 ),
    .o({\u2_Display/add156/c22 ,\u2_Display/n5121 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u22  (
    .a(\u2_Display/n6254 ),
    .b(1'b1),
    .c(\u2_Display/add156/c22 ),
    .o({\u2_Display/add156/c23 ,\u2_Display/n5121 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u23  (
    .a(\u2_Display/n6253 ),
    .b(1'b0),
    .c(\u2_Display/add156/c23 ),
    .o({\u2_Display/add156/c24 ,\u2_Display/n5121 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u24  (
    .a(\u2_Display/n6252 ),
    .b(1'b1),
    .c(\u2_Display/add156/c24 ),
    .o({\u2_Display/add156/c25 ,\u2_Display/n5121 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u25  (
    .a(\u2_Display/n6251 ),
    .b(1'b0),
    .c(\u2_Display/add156/c25 ),
    .o({\u2_Display/add156/c26 ,\u2_Display/n5121 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u26  (
    .a(\u2_Display/n6250 ),
    .b(1'b1),
    .c(\u2_Display/add156/c26 ),
    .o({\u2_Display/add156/c27 ,\u2_Display/n5121 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u27  (
    .a(\u2_Display/n6249 ),
    .b(1'b1),
    .c(\u2_Display/add156/c27 ),
    .o({\u2_Display/add156/c28 ,\u2_Display/n5121 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u28  (
    .a(\u2_Display/n6248 ),
    .b(1'b1),
    .c(\u2_Display/add156/c28 ),
    .o({\u2_Display/add156/c29 ,\u2_Display/n5121 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u29  (
    .a(\u2_Display/n6247 ),
    .b(1'b1),
    .c(\u2_Display/add156/c29 ),
    .o({\u2_Display/add156/c30 ,\u2_Display/n5121 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u3  (
    .a(\u2_Display/n6273 ),
    .b(1'b1),
    .c(\u2_Display/add156/c3 ),
    .o({\u2_Display/add156/c4 ,\u2_Display/n5121 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u30  (
    .a(\u2_Display/n6246 ),
    .b(1'b1),
    .c(\u2_Display/add156/c30 ),
    .o({\u2_Display/add156/c31 ,\u2_Display/n5121 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u31  (
    .a(\u2_Display/n6245 ),
    .b(1'b1),
    .c(\u2_Display/add156/c31 ),
    .o({open_n1023,\u2_Display/n5121 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u4  (
    .a(\u2_Display/n6272 ),
    .b(1'b1),
    .c(\u2_Display/add156/c4 ),
    .o({\u2_Display/add156/c5 ,\u2_Display/n5121 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u5  (
    .a(\u2_Display/n6271 ),
    .b(1'b1),
    .c(\u2_Display/add156/c5 ),
    .o({\u2_Display/add156/c6 ,\u2_Display/n5121 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u6  (
    .a(\u2_Display/n6270 ),
    .b(1'b1),
    .c(\u2_Display/add156/c6 ),
    .o({\u2_Display/add156/c7 ,\u2_Display/n5121 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u7  (
    .a(\u2_Display/n6269 ),
    .b(1'b1),
    .c(\u2_Display/add156/c7 ),
    .o({\u2_Display/add156/c8 ,\u2_Display/n5121 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u8  (
    .a(\u2_Display/n6268 ),
    .b(1'b1),
    .c(\u2_Display/add156/c8 ),
    .o({\u2_Display/add156/c9 ,\u2_Display/n5121 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add156/u9  (
    .a(\u2_Display/n6267 ),
    .b(1'b1),
    .c(\u2_Display/add156/c9 ),
    .o({\u2_Display/add156/c10 ,\u2_Display/n5121 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add156/ucin  (
    .a(1'b1),
    .o({\u2_Display/add156/c0 ,open_n1026}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u0  (
    .a(\u2_Display/n6311 ),
    .b(1'b1),
    .c(\u2_Display/add157/c0 ),
    .o({\u2_Display/add157/c1 ,\u2_Display/n5156 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u1  (
    .a(\u2_Display/n6310 ),
    .b(1'b1),
    .c(\u2_Display/add157/c1 ),
    .o({\u2_Display/add157/c2 ,\u2_Display/n5156 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u10  (
    .a(\u2_Display/n6301 ),
    .b(1'b1),
    .c(\u2_Display/add157/c10 ),
    .o({\u2_Display/add157/c11 ,\u2_Display/n5156 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u11  (
    .a(\u2_Display/n6300 ),
    .b(1'b1),
    .c(\u2_Display/add157/c11 ),
    .o({\u2_Display/add157/c12 ,\u2_Display/n5156 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u12  (
    .a(\u2_Display/n6299 ),
    .b(1'b1),
    .c(\u2_Display/add157/c12 ),
    .o({\u2_Display/add157/c13 ,\u2_Display/n5156 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u13  (
    .a(\u2_Display/n6298 ),
    .b(1'b1),
    .c(\u2_Display/add157/c13 ),
    .o({\u2_Display/add157/c14 ,\u2_Display/n5156 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u14  (
    .a(\u2_Display/n6297 ),
    .b(1'b1),
    .c(\u2_Display/add157/c14 ),
    .o({\u2_Display/add157/c15 ,\u2_Display/n5156 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u15  (
    .a(\u2_Display/n6296 ),
    .b(1'b1),
    .c(\u2_Display/add157/c15 ),
    .o({\u2_Display/add157/c16 ,\u2_Display/n5156 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u16  (
    .a(\u2_Display/n6295 ),
    .b(1'b1),
    .c(\u2_Display/add157/c16 ),
    .o({\u2_Display/add157/c17 ,\u2_Display/n5156 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u17  (
    .a(\u2_Display/n6294 ),
    .b(1'b1),
    .c(\u2_Display/add157/c17 ),
    .o({\u2_Display/add157/c18 ,\u2_Display/n5156 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u18  (
    .a(\u2_Display/n6293 ),
    .b(1'b1),
    .c(\u2_Display/add157/c18 ),
    .o({\u2_Display/add157/c19 ,\u2_Display/n5156 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u19  (
    .a(\u2_Display/n6292 ),
    .b(1'b1),
    .c(\u2_Display/add157/c19 ),
    .o({\u2_Display/add157/c20 ,\u2_Display/n5156 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u2  (
    .a(\u2_Display/n6309 ),
    .b(1'b1),
    .c(\u2_Display/add157/c2 ),
    .o({\u2_Display/add157/c3 ,\u2_Display/n5156 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u20  (
    .a(\u2_Display/n6291 ),
    .b(1'b1),
    .c(\u2_Display/add157/c20 ),
    .o({\u2_Display/add157/c21 ,\u2_Display/n5156 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u21  (
    .a(\u2_Display/n6290 ),
    .b(1'b1),
    .c(\u2_Display/add157/c21 ),
    .o({\u2_Display/add157/c22 ,\u2_Display/n5156 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u22  (
    .a(\u2_Display/n6289 ),
    .b(1'b0),
    .c(\u2_Display/add157/c22 ),
    .o({\u2_Display/add157/c23 ,\u2_Display/n5156 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u23  (
    .a(\u2_Display/n6288 ),
    .b(1'b1),
    .c(\u2_Display/add157/c23 ),
    .o({\u2_Display/add157/c24 ,\u2_Display/n5156 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u24  (
    .a(\u2_Display/n6287 ),
    .b(1'b0),
    .c(\u2_Display/add157/c24 ),
    .o({\u2_Display/add157/c25 ,\u2_Display/n5156 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u25  (
    .a(\u2_Display/n6286 ),
    .b(1'b1),
    .c(\u2_Display/add157/c25 ),
    .o({\u2_Display/add157/c26 ,\u2_Display/n5156 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u26  (
    .a(\u2_Display/n6285 ),
    .b(1'b1),
    .c(\u2_Display/add157/c26 ),
    .o({\u2_Display/add157/c27 ,\u2_Display/n5156 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u27  (
    .a(\u2_Display/n6284 ),
    .b(1'b1),
    .c(\u2_Display/add157/c27 ),
    .o({\u2_Display/add157/c28 ,\u2_Display/n5156 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u28  (
    .a(\u2_Display/n6283 ),
    .b(1'b1),
    .c(\u2_Display/add157/c28 ),
    .o({\u2_Display/add157/c29 ,\u2_Display/n5156 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u29  (
    .a(\u2_Display/n6282 ),
    .b(1'b1),
    .c(\u2_Display/add157/c29 ),
    .o({\u2_Display/add157/c30 ,\u2_Display/n5156 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u3  (
    .a(\u2_Display/n6308 ),
    .b(1'b1),
    .c(\u2_Display/add157/c3 ),
    .o({\u2_Display/add157/c4 ,\u2_Display/n5156 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u30  (
    .a(\u2_Display/n6281 ),
    .b(1'b1),
    .c(\u2_Display/add157/c30 ),
    .o({\u2_Display/add157/c31 ,\u2_Display/n5156 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u31  (
    .a(\u2_Display/n6280 ),
    .b(1'b1),
    .c(\u2_Display/add157/c31 ),
    .o({open_n1027,\u2_Display/n5156 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u4  (
    .a(\u2_Display/n6307 ),
    .b(1'b1),
    .c(\u2_Display/add157/c4 ),
    .o({\u2_Display/add157/c5 ,\u2_Display/n5156 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u5  (
    .a(\u2_Display/n6306 ),
    .b(1'b1),
    .c(\u2_Display/add157/c5 ),
    .o({\u2_Display/add157/c6 ,\u2_Display/n5156 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u6  (
    .a(\u2_Display/n6305 ),
    .b(1'b1),
    .c(\u2_Display/add157/c6 ),
    .o({\u2_Display/add157/c7 ,\u2_Display/n5156 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u7  (
    .a(\u2_Display/n6304 ),
    .b(1'b1),
    .c(\u2_Display/add157/c7 ),
    .o({\u2_Display/add157/c8 ,\u2_Display/n5156 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u8  (
    .a(\u2_Display/n6303 ),
    .b(1'b1),
    .c(\u2_Display/add157/c8 ),
    .o({\u2_Display/add157/c9 ,\u2_Display/n5156 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add157/u9  (
    .a(\u2_Display/n6302 ),
    .b(1'b1),
    .c(\u2_Display/add157/c9 ),
    .o({\u2_Display/add157/c10 ,\u2_Display/n5156 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add157/ucin  (
    .a(1'b1),
    .o({\u2_Display/add157/c0 ,open_n1030}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u0  (
    .a(\u2_Display/n6346 ),
    .b(1'b1),
    .c(\u2_Display/add158/c0 ),
    .o({\u2_Display/add158/c1 ,\u2_Display/n5191 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u1  (
    .a(\u2_Display/n6345 ),
    .b(1'b1),
    .c(\u2_Display/add158/c1 ),
    .o({\u2_Display/add158/c2 ,\u2_Display/n5191 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u10  (
    .a(\u2_Display/n6336 ),
    .b(1'b1),
    .c(\u2_Display/add158/c10 ),
    .o({\u2_Display/add158/c11 ,\u2_Display/n5191 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u11  (
    .a(\u2_Display/n6335 ),
    .b(1'b1),
    .c(\u2_Display/add158/c11 ),
    .o({\u2_Display/add158/c12 ,\u2_Display/n5191 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u12  (
    .a(\u2_Display/n6334 ),
    .b(1'b1),
    .c(\u2_Display/add158/c12 ),
    .o({\u2_Display/add158/c13 ,\u2_Display/n5191 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u13  (
    .a(\u2_Display/n6333 ),
    .b(1'b1),
    .c(\u2_Display/add158/c13 ),
    .o({\u2_Display/add158/c14 ,\u2_Display/n5191 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u14  (
    .a(\u2_Display/n6332 ),
    .b(1'b1),
    .c(\u2_Display/add158/c14 ),
    .o({\u2_Display/add158/c15 ,\u2_Display/n5191 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u15  (
    .a(\u2_Display/n6331 ),
    .b(1'b1),
    .c(\u2_Display/add158/c15 ),
    .o({\u2_Display/add158/c16 ,\u2_Display/n5191 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u16  (
    .a(\u2_Display/n6330 ),
    .b(1'b1),
    .c(\u2_Display/add158/c16 ),
    .o({\u2_Display/add158/c17 ,\u2_Display/n5191 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u17  (
    .a(\u2_Display/n6329 ),
    .b(1'b1),
    .c(\u2_Display/add158/c17 ),
    .o({\u2_Display/add158/c18 ,\u2_Display/n5191 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u18  (
    .a(\u2_Display/n6328 ),
    .b(1'b1),
    .c(\u2_Display/add158/c18 ),
    .o({\u2_Display/add158/c19 ,\u2_Display/n5191 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u19  (
    .a(\u2_Display/n6327 ),
    .b(1'b1),
    .c(\u2_Display/add158/c19 ),
    .o({\u2_Display/add158/c20 ,\u2_Display/n5191 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u2  (
    .a(\u2_Display/n6344 ),
    .b(1'b1),
    .c(\u2_Display/add158/c2 ),
    .o({\u2_Display/add158/c3 ,\u2_Display/n5191 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u20  (
    .a(\u2_Display/n6326 ),
    .b(1'b1),
    .c(\u2_Display/add158/c20 ),
    .o({\u2_Display/add158/c21 ,\u2_Display/n5191 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u21  (
    .a(\u2_Display/n6325 ),
    .b(1'b0),
    .c(\u2_Display/add158/c21 ),
    .o({\u2_Display/add158/c22 ,\u2_Display/n5191 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u22  (
    .a(\u2_Display/n6324 ),
    .b(1'b1),
    .c(\u2_Display/add158/c22 ),
    .o({\u2_Display/add158/c23 ,\u2_Display/n5191 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u23  (
    .a(\u2_Display/n6323 ),
    .b(1'b0),
    .c(\u2_Display/add158/c23 ),
    .o({\u2_Display/add158/c24 ,\u2_Display/n5191 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u24  (
    .a(\u2_Display/n6322 ),
    .b(1'b1),
    .c(\u2_Display/add158/c24 ),
    .o({\u2_Display/add158/c25 ,\u2_Display/n5191 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u25  (
    .a(\u2_Display/n6321 ),
    .b(1'b1),
    .c(\u2_Display/add158/c25 ),
    .o({\u2_Display/add158/c26 ,\u2_Display/n5191 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u26  (
    .a(\u2_Display/n6320 ),
    .b(1'b1),
    .c(\u2_Display/add158/c26 ),
    .o({\u2_Display/add158/c27 ,\u2_Display/n5191 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u27  (
    .a(\u2_Display/n6319 ),
    .b(1'b1),
    .c(\u2_Display/add158/c27 ),
    .o({\u2_Display/add158/c28 ,\u2_Display/n5191 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u28  (
    .a(\u2_Display/n6318 ),
    .b(1'b1),
    .c(\u2_Display/add158/c28 ),
    .o({\u2_Display/add158/c29 ,\u2_Display/n5191 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u29  (
    .a(\u2_Display/n6317 ),
    .b(1'b1),
    .c(\u2_Display/add158/c29 ),
    .o({\u2_Display/add158/c30 ,\u2_Display/n5191 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u3  (
    .a(\u2_Display/n6343 ),
    .b(1'b1),
    .c(\u2_Display/add158/c3 ),
    .o({\u2_Display/add158/c4 ,\u2_Display/n5191 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u30  (
    .a(\u2_Display/n6316 ),
    .b(1'b1),
    .c(\u2_Display/add158/c30 ),
    .o({\u2_Display/add158/c31 ,\u2_Display/n5191 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u31  (
    .a(\u2_Display/n6315 ),
    .b(1'b1),
    .c(\u2_Display/add158/c31 ),
    .o({open_n1031,\u2_Display/n5191 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u4  (
    .a(\u2_Display/n6342 ),
    .b(1'b1),
    .c(\u2_Display/add158/c4 ),
    .o({\u2_Display/add158/c5 ,\u2_Display/n5191 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u5  (
    .a(\u2_Display/n6341 ),
    .b(1'b1),
    .c(\u2_Display/add158/c5 ),
    .o({\u2_Display/add158/c6 ,\u2_Display/n5191 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u6  (
    .a(\u2_Display/n6340 ),
    .b(1'b1),
    .c(\u2_Display/add158/c6 ),
    .o({\u2_Display/add158/c7 ,\u2_Display/n5191 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u7  (
    .a(\u2_Display/n6339 ),
    .b(1'b1),
    .c(\u2_Display/add158/c7 ),
    .o({\u2_Display/add158/c8 ,\u2_Display/n5191 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u8  (
    .a(\u2_Display/n6338 ),
    .b(1'b1),
    .c(\u2_Display/add158/c8 ),
    .o({\u2_Display/add158/c9 ,\u2_Display/n5191 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add158/u9  (
    .a(\u2_Display/n6337 ),
    .b(1'b1),
    .c(\u2_Display/add158/c9 ),
    .o({\u2_Display/add158/c10 ,\u2_Display/n5191 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add158/ucin  (
    .a(1'b1),
    .o({\u2_Display/add158/c0 ,open_n1034}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u0  (
    .a(\u2_Display/n5223 ),
    .b(1'b1),
    .c(\u2_Display/add159/c0 ),
    .o({\u2_Display/add159/c1 ,\u2_Display/n5226 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u1  (
    .a(\u2_Display/n5222 ),
    .b(1'b1),
    .c(\u2_Display/add159/c1 ),
    .o({\u2_Display/add159/c2 ,\u2_Display/n5226 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u10  (
    .a(\u2_Display/n5213 ),
    .b(1'b1),
    .c(\u2_Display/add159/c10 ),
    .o({\u2_Display/add159/c11 ,\u2_Display/n5226 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u11  (
    .a(\u2_Display/n5212 ),
    .b(1'b1),
    .c(\u2_Display/add159/c11 ),
    .o({\u2_Display/add159/c12 ,\u2_Display/n5226 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u12  (
    .a(\u2_Display/n5211 ),
    .b(1'b1),
    .c(\u2_Display/add159/c12 ),
    .o({\u2_Display/add159/c13 ,\u2_Display/n5226 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u13  (
    .a(\u2_Display/n5210 ),
    .b(1'b1),
    .c(\u2_Display/add159/c13 ),
    .o({\u2_Display/add159/c14 ,\u2_Display/n5226 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u14  (
    .a(\u2_Display/n5209 ),
    .b(1'b1),
    .c(\u2_Display/add159/c14 ),
    .o({\u2_Display/add159/c15 ,\u2_Display/n5226 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u15  (
    .a(\u2_Display/n5208 ),
    .b(1'b1),
    .c(\u2_Display/add159/c15 ),
    .o({\u2_Display/add159/c16 ,\u2_Display/n5226 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u16  (
    .a(\u2_Display/n5207 ),
    .b(1'b1),
    .c(\u2_Display/add159/c16 ),
    .o({\u2_Display/add159/c17 ,\u2_Display/n5226 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u17  (
    .a(\u2_Display/n5206 ),
    .b(1'b1),
    .c(\u2_Display/add159/c17 ),
    .o({\u2_Display/add159/c18 ,\u2_Display/n5226 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u18  (
    .a(\u2_Display/n5205 ),
    .b(1'b1),
    .c(\u2_Display/add159/c18 ),
    .o({\u2_Display/add159/c19 ,\u2_Display/n5226 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u19  (
    .a(\u2_Display/n5204 ),
    .b(1'b1),
    .c(\u2_Display/add159/c19 ),
    .o({\u2_Display/add159/c20 ,\u2_Display/n5226 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u2  (
    .a(\u2_Display/n5221 ),
    .b(1'b1),
    .c(\u2_Display/add159/c2 ),
    .o({\u2_Display/add159/c3 ,\u2_Display/n5226 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u20  (
    .a(\u2_Display/n5203 ),
    .b(1'b0),
    .c(\u2_Display/add159/c20 ),
    .o({\u2_Display/add159/c21 ,\u2_Display/n5226 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u21  (
    .a(\u2_Display/n5202 ),
    .b(1'b1),
    .c(\u2_Display/add159/c21 ),
    .o({\u2_Display/add159/c22 ,\u2_Display/n5226 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u22  (
    .a(\u2_Display/n5201 ),
    .b(1'b0),
    .c(\u2_Display/add159/c22 ),
    .o({\u2_Display/add159/c23 ,\u2_Display/n5226 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u23  (
    .a(\u2_Display/n5200 ),
    .b(1'b1),
    .c(\u2_Display/add159/c23 ),
    .o({\u2_Display/add159/c24 ,\u2_Display/n5226 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u24  (
    .a(\u2_Display/n5199 ),
    .b(1'b1),
    .c(\u2_Display/add159/c24 ),
    .o({\u2_Display/add159/c25 ,\u2_Display/n5226 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u25  (
    .a(\u2_Display/n5198 ),
    .b(1'b1),
    .c(\u2_Display/add159/c25 ),
    .o({\u2_Display/add159/c26 ,\u2_Display/n5226 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u26  (
    .a(\u2_Display/n5197 ),
    .b(1'b1),
    .c(\u2_Display/add159/c26 ),
    .o({\u2_Display/add159/c27 ,\u2_Display/n5226 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u27  (
    .a(\u2_Display/n5196 ),
    .b(1'b1),
    .c(\u2_Display/add159/c27 ),
    .o({\u2_Display/add159/c28 ,\u2_Display/n5226 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u28  (
    .a(\u2_Display/n6353 ),
    .b(1'b1),
    .c(\u2_Display/add159/c28 ),
    .o({\u2_Display/add159/c29 ,\u2_Display/n5226 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u29  (
    .a(\u2_Display/n6352 ),
    .b(1'b1),
    .c(\u2_Display/add159/c29 ),
    .o({\u2_Display/add159/c30 ,\u2_Display/n5226 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u3  (
    .a(\u2_Display/n5220 ),
    .b(1'b1),
    .c(\u2_Display/add159/c3 ),
    .o({\u2_Display/add159/c4 ,\u2_Display/n5226 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u30  (
    .a(\u2_Display/n6351 ),
    .b(1'b1),
    .c(\u2_Display/add159/c30 ),
    .o({\u2_Display/add159/c31 ,\u2_Display/n5226 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u31  (
    .a(\u2_Display/n6350 ),
    .b(1'b1),
    .c(\u2_Display/add159/c31 ),
    .o({open_n1035,\u2_Display/n5226 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u4  (
    .a(\u2_Display/n5219 ),
    .b(1'b1),
    .c(\u2_Display/add159/c4 ),
    .o({\u2_Display/add159/c5 ,\u2_Display/n5226 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u5  (
    .a(\u2_Display/n5218 ),
    .b(1'b1),
    .c(\u2_Display/add159/c5 ),
    .o({\u2_Display/add159/c6 ,\u2_Display/n5226 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u6  (
    .a(\u2_Display/n5217 ),
    .b(1'b1),
    .c(\u2_Display/add159/c6 ),
    .o({\u2_Display/add159/c7 ,\u2_Display/n5226 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u7  (
    .a(\u2_Display/n5216 ),
    .b(1'b1),
    .c(\u2_Display/add159/c7 ),
    .o({\u2_Display/add159/c8 ,\u2_Display/n5226 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u8  (
    .a(\u2_Display/n5215 ),
    .b(1'b1),
    .c(\u2_Display/add159/c8 ),
    .o({\u2_Display/add159/c9 ,\u2_Display/n5226 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add159/u9  (
    .a(\u2_Display/n5214 ),
    .b(1'b1),
    .c(\u2_Display/add159/c9 ),
    .o({\u2_Display/add159/c10 ,\u2_Display/n5226 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add159/ucin  (
    .a(1'b1),
    .o({\u2_Display/add159/c0 ,open_n1038}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u0  (
    .a(\u2_Display/n5258 ),
    .b(1'b1),
    .c(\u2_Display/add160/c0 ),
    .o({\u2_Display/add160/c1 ,\u2_Display/n5261 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u1  (
    .a(\u2_Display/n5257 ),
    .b(1'b1),
    .c(\u2_Display/add160/c1 ),
    .o({\u2_Display/add160/c2 ,\u2_Display/n5261 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u10  (
    .a(\u2_Display/n5248 ),
    .b(1'b1),
    .c(\u2_Display/add160/c10 ),
    .o({\u2_Display/add160/c11 ,\u2_Display/n5261 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u11  (
    .a(\u2_Display/n5247 ),
    .b(1'b1),
    .c(\u2_Display/add160/c11 ),
    .o({\u2_Display/add160/c12 ,\u2_Display/n5261 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u12  (
    .a(\u2_Display/n5246 ),
    .b(1'b1),
    .c(\u2_Display/add160/c12 ),
    .o({\u2_Display/add160/c13 ,\u2_Display/n5261 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u13  (
    .a(\u2_Display/n5245 ),
    .b(1'b1),
    .c(\u2_Display/add160/c13 ),
    .o({\u2_Display/add160/c14 ,\u2_Display/n5261 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u14  (
    .a(\u2_Display/n5244 ),
    .b(1'b1),
    .c(\u2_Display/add160/c14 ),
    .o({\u2_Display/add160/c15 ,\u2_Display/n5261 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u15  (
    .a(\u2_Display/n5243 ),
    .b(1'b1),
    .c(\u2_Display/add160/c15 ),
    .o({\u2_Display/add160/c16 ,\u2_Display/n5261 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u16  (
    .a(\u2_Display/n5242 ),
    .b(1'b1),
    .c(\u2_Display/add160/c16 ),
    .o({\u2_Display/add160/c17 ,\u2_Display/n5261 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u17  (
    .a(\u2_Display/n5241 ),
    .b(1'b1),
    .c(\u2_Display/add160/c17 ),
    .o({\u2_Display/add160/c18 ,\u2_Display/n5261 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u18  (
    .a(\u2_Display/n5240 ),
    .b(1'b1),
    .c(\u2_Display/add160/c18 ),
    .o({\u2_Display/add160/c19 ,\u2_Display/n5261 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u19  (
    .a(\u2_Display/n5239 ),
    .b(1'b0),
    .c(\u2_Display/add160/c19 ),
    .o({\u2_Display/add160/c20 ,\u2_Display/n5261 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u2  (
    .a(\u2_Display/n5256 ),
    .b(1'b1),
    .c(\u2_Display/add160/c2 ),
    .o({\u2_Display/add160/c3 ,\u2_Display/n5261 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u20  (
    .a(\u2_Display/n5238 ),
    .b(1'b1),
    .c(\u2_Display/add160/c20 ),
    .o({\u2_Display/add160/c21 ,\u2_Display/n5261 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u21  (
    .a(\u2_Display/n5237 ),
    .b(1'b0),
    .c(\u2_Display/add160/c21 ),
    .o({\u2_Display/add160/c22 ,\u2_Display/n5261 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u22  (
    .a(\u2_Display/n5236 ),
    .b(1'b1),
    .c(\u2_Display/add160/c22 ),
    .o({\u2_Display/add160/c23 ,\u2_Display/n5261 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u23  (
    .a(\u2_Display/n5235 ),
    .b(1'b1),
    .c(\u2_Display/add160/c23 ),
    .o({\u2_Display/add160/c24 ,\u2_Display/n5261 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u24  (
    .a(\u2_Display/n5234 ),
    .b(1'b1),
    .c(\u2_Display/add160/c24 ),
    .o({\u2_Display/add160/c25 ,\u2_Display/n5261 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u25  (
    .a(\u2_Display/n5233 ),
    .b(1'b1),
    .c(\u2_Display/add160/c25 ),
    .o({\u2_Display/add160/c26 ,\u2_Display/n5261 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u26  (
    .a(\u2_Display/n5232 ),
    .b(1'b1),
    .c(\u2_Display/add160/c26 ),
    .o({\u2_Display/add160/c27 ,\u2_Display/n5261 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u27  (
    .a(\u2_Display/n5231 ),
    .b(1'b1),
    .c(\u2_Display/add160/c27 ),
    .o({\u2_Display/add160/c28 ,\u2_Display/n5261 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u28  (
    .a(\u2_Display/n5230 ),
    .b(1'b1),
    .c(\u2_Display/add160/c28 ),
    .o({\u2_Display/add160/c29 ,\u2_Display/n5261 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u29  (
    .a(\u2_Display/n5229 ),
    .b(1'b1),
    .c(\u2_Display/add160/c29 ),
    .o({\u2_Display/add160/c30 ,\u2_Display/n5261 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u3  (
    .a(\u2_Display/n5255 ),
    .b(1'b1),
    .c(\u2_Display/add160/c3 ),
    .o({\u2_Display/add160/c4 ,\u2_Display/n5261 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u30  (
    .a(\u2_Display/n5228 ),
    .b(1'b1),
    .c(\u2_Display/add160/c30 ),
    .o({\u2_Display/add160/c31 ,\u2_Display/n5261 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u31  (
    .a(\u2_Display/n5227 ),
    .b(1'b1),
    .c(\u2_Display/add160/c31 ),
    .o({open_n1039,\u2_Display/n5261 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u4  (
    .a(\u2_Display/n5254 ),
    .b(1'b1),
    .c(\u2_Display/add160/c4 ),
    .o({\u2_Display/add160/c5 ,\u2_Display/n5261 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u5  (
    .a(\u2_Display/n5253 ),
    .b(1'b1),
    .c(\u2_Display/add160/c5 ),
    .o({\u2_Display/add160/c6 ,\u2_Display/n5261 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u6  (
    .a(\u2_Display/n5252 ),
    .b(1'b1),
    .c(\u2_Display/add160/c6 ),
    .o({\u2_Display/add160/c7 ,\u2_Display/n5261 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u7  (
    .a(\u2_Display/n5251 ),
    .b(1'b1),
    .c(\u2_Display/add160/c7 ),
    .o({\u2_Display/add160/c8 ,\u2_Display/n5261 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u8  (
    .a(\u2_Display/n5250 ),
    .b(1'b1),
    .c(\u2_Display/add160/c8 ),
    .o({\u2_Display/add160/c9 ,\u2_Display/n5261 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add160/u9  (
    .a(\u2_Display/n5249 ),
    .b(1'b1),
    .c(\u2_Display/add160/c9 ),
    .o({\u2_Display/add160/c10 ,\u2_Display/n5261 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add160/ucin  (
    .a(1'b1),
    .o({\u2_Display/add160/c0 ,open_n1042}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u0  (
    .a(\u2_Display/n5293 ),
    .b(1'b1),
    .c(\u2_Display/add161/c0 ),
    .o({\u2_Display/add161/c1 ,\u2_Display/n5296 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u1  (
    .a(\u2_Display/n5292 ),
    .b(1'b1),
    .c(\u2_Display/add161/c1 ),
    .o({\u2_Display/add161/c2 ,\u2_Display/n5296 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u10  (
    .a(\u2_Display/n5283 ),
    .b(1'b1),
    .c(\u2_Display/add161/c10 ),
    .o({\u2_Display/add161/c11 ,\u2_Display/n5296 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u11  (
    .a(\u2_Display/n5282 ),
    .b(1'b1),
    .c(\u2_Display/add161/c11 ),
    .o({\u2_Display/add161/c12 ,\u2_Display/n5296 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u12  (
    .a(\u2_Display/n5281 ),
    .b(1'b1),
    .c(\u2_Display/add161/c12 ),
    .o({\u2_Display/add161/c13 ,\u2_Display/n5296 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u13  (
    .a(\u2_Display/n5280 ),
    .b(1'b1),
    .c(\u2_Display/add161/c13 ),
    .o({\u2_Display/add161/c14 ,\u2_Display/n5296 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u14  (
    .a(\u2_Display/n5279 ),
    .b(1'b1),
    .c(\u2_Display/add161/c14 ),
    .o({\u2_Display/add161/c15 ,\u2_Display/n5296 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u15  (
    .a(\u2_Display/n5278 ),
    .b(1'b1),
    .c(\u2_Display/add161/c15 ),
    .o({\u2_Display/add161/c16 ,\u2_Display/n5296 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u16  (
    .a(\u2_Display/n5277 ),
    .b(1'b1),
    .c(\u2_Display/add161/c16 ),
    .o({\u2_Display/add161/c17 ,\u2_Display/n5296 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u17  (
    .a(\u2_Display/n5276 ),
    .b(1'b1),
    .c(\u2_Display/add161/c17 ),
    .o({\u2_Display/add161/c18 ,\u2_Display/n5296 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u18  (
    .a(\u2_Display/n5275 ),
    .b(1'b0),
    .c(\u2_Display/add161/c18 ),
    .o({\u2_Display/add161/c19 ,\u2_Display/n5296 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u19  (
    .a(\u2_Display/n5274 ),
    .b(1'b1),
    .c(\u2_Display/add161/c19 ),
    .o({\u2_Display/add161/c20 ,\u2_Display/n5296 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u2  (
    .a(\u2_Display/n5291 ),
    .b(1'b1),
    .c(\u2_Display/add161/c2 ),
    .o({\u2_Display/add161/c3 ,\u2_Display/n5296 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u20  (
    .a(\u2_Display/n5273 ),
    .b(1'b0),
    .c(\u2_Display/add161/c20 ),
    .o({\u2_Display/add161/c21 ,\u2_Display/n5296 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u21  (
    .a(\u2_Display/n5272 ),
    .b(1'b1),
    .c(\u2_Display/add161/c21 ),
    .o({\u2_Display/add161/c22 ,\u2_Display/n5296 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u22  (
    .a(\u2_Display/n5271 ),
    .b(1'b1),
    .c(\u2_Display/add161/c22 ),
    .o({\u2_Display/add161/c23 ,\u2_Display/n5296 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u23  (
    .a(\u2_Display/n5270 ),
    .b(1'b1),
    .c(\u2_Display/add161/c23 ),
    .o({\u2_Display/add161/c24 ,\u2_Display/n5296 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u24  (
    .a(\u2_Display/n5269 ),
    .b(1'b1),
    .c(\u2_Display/add161/c24 ),
    .o({\u2_Display/add161/c25 ,\u2_Display/n5296 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u25  (
    .a(\u2_Display/n5268 ),
    .b(1'b1),
    .c(\u2_Display/add161/c25 ),
    .o({\u2_Display/add161/c26 ,\u2_Display/n5296 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u26  (
    .a(\u2_Display/n5267 ),
    .b(1'b1),
    .c(\u2_Display/add161/c26 ),
    .o({\u2_Display/add161/c27 ,\u2_Display/n5296 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u27  (
    .a(\u2_Display/n5266 ),
    .b(1'b1),
    .c(\u2_Display/add161/c27 ),
    .o({\u2_Display/add161/c28 ,\u2_Display/n5296 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u28  (
    .a(\u2_Display/n5265 ),
    .b(1'b1),
    .c(\u2_Display/add161/c28 ),
    .o({\u2_Display/add161/c29 ,\u2_Display/n5296 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u29  (
    .a(\u2_Display/n5264 ),
    .b(1'b1),
    .c(\u2_Display/add161/c29 ),
    .o({\u2_Display/add161/c30 ,\u2_Display/n5296 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u3  (
    .a(\u2_Display/n5290 ),
    .b(1'b1),
    .c(\u2_Display/add161/c3 ),
    .o({\u2_Display/add161/c4 ,\u2_Display/n5296 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u30  (
    .a(\u2_Display/n5263 ),
    .b(1'b1),
    .c(\u2_Display/add161/c30 ),
    .o({\u2_Display/add161/c31 ,\u2_Display/n5296 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u31  (
    .a(\u2_Display/n5262 ),
    .b(1'b1),
    .c(\u2_Display/add161/c31 ),
    .o({open_n1043,\u2_Display/n5296 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u4  (
    .a(\u2_Display/n5289 ),
    .b(1'b1),
    .c(\u2_Display/add161/c4 ),
    .o({\u2_Display/add161/c5 ,\u2_Display/n5296 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u5  (
    .a(\u2_Display/n5288 ),
    .b(1'b1),
    .c(\u2_Display/add161/c5 ),
    .o({\u2_Display/add161/c6 ,\u2_Display/n5296 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u6  (
    .a(\u2_Display/n5287 ),
    .b(1'b1),
    .c(\u2_Display/add161/c6 ),
    .o({\u2_Display/add161/c7 ,\u2_Display/n5296 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u7  (
    .a(\u2_Display/n5286 ),
    .b(1'b1),
    .c(\u2_Display/add161/c7 ),
    .o({\u2_Display/add161/c8 ,\u2_Display/n5296 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u8  (
    .a(\u2_Display/n5285 ),
    .b(1'b1),
    .c(\u2_Display/add161/c8 ),
    .o({\u2_Display/add161/c9 ,\u2_Display/n5296 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add161/u9  (
    .a(\u2_Display/n5284 ),
    .b(1'b1),
    .c(\u2_Display/add161/c9 ),
    .o({\u2_Display/add161/c10 ,\u2_Display/n5296 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add161/ucin  (
    .a(1'b1),
    .o({\u2_Display/add161/c0 ,open_n1046}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u0  (
    .a(\u2_Display/n5328 ),
    .b(1'b1),
    .c(\u2_Display/add162/c0 ),
    .o({\u2_Display/add162/c1 ,\u2_Display/n5331 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u1  (
    .a(\u2_Display/n5327 ),
    .b(1'b1),
    .c(\u2_Display/add162/c1 ),
    .o({\u2_Display/add162/c2 ,\u2_Display/n5331 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u10  (
    .a(\u2_Display/n5318 ),
    .b(1'b1),
    .c(\u2_Display/add162/c10 ),
    .o({\u2_Display/add162/c11 ,\u2_Display/n5331 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u11  (
    .a(\u2_Display/n5317 ),
    .b(1'b1),
    .c(\u2_Display/add162/c11 ),
    .o({\u2_Display/add162/c12 ,\u2_Display/n5331 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u12  (
    .a(\u2_Display/n5316 ),
    .b(1'b1),
    .c(\u2_Display/add162/c12 ),
    .o({\u2_Display/add162/c13 ,\u2_Display/n5331 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u13  (
    .a(\u2_Display/n5315 ),
    .b(1'b1),
    .c(\u2_Display/add162/c13 ),
    .o({\u2_Display/add162/c14 ,\u2_Display/n5331 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u14  (
    .a(\u2_Display/n5314 ),
    .b(1'b1),
    .c(\u2_Display/add162/c14 ),
    .o({\u2_Display/add162/c15 ,\u2_Display/n5331 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u15  (
    .a(\u2_Display/n5313 ),
    .b(1'b1),
    .c(\u2_Display/add162/c15 ),
    .o({\u2_Display/add162/c16 ,\u2_Display/n5331 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u16  (
    .a(\u2_Display/n5312 ),
    .b(1'b1),
    .c(\u2_Display/add162/c16 ),
    .o({\u2_Display/add162/c17 ,\u2_Display/n5331 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u17  (
    .a(\u2_Display/n5311 ),
    .b(1'b0),
    .c(\u2_Display/add162/c17 ),
    .o({\u2_Display/add162/c18 ,\u2_Display/n5331 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u18  (
    .a(\u2_Display/n5310 ),
    .b(1'b1),
    .c(\u2_Display/add162/c18 ),
    .o({\u2_Display/add162/c19 ,\u2_Display/n5331 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u19  (
    .a(\u2_Display/n5309 ),
    .b(1'b0),
    .c(\u2_Display/add162/c19 ),
    .o({\u2_Display/add162/c20 ,\u2_Display/n5331 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u2  (
    .a(\u2_Display/n5326 ),
    .b(1'b1),
    .c(\u2_Display/add162/c2 ),
    .o({\u2_Display/add162/c3 ,\u2_Display/n5331 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u20  (
    .a(\u2_Display/n5308 ),
    .b(1'b1),
    .c(\u2_Display/add162/c20 ),
    .o({\u2_Display/add162/c21 ,\u2_Display/n5331 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u21  (
    .a(\u2_Display/n5307 ),
    .b(1'b1),
    .c(\u2_Display/add162/c21 ),
    .o({\u2_Display/add162/c22 ,\u2_Display/n5331 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u22  (
    .a(\u2_Display/n5306 ),
    .b(1'b1),
    .c(\u2_Display/add162/c22 ),
    .o({\u2_Display/add162/c23 ,\u2_Display/n5331 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u23  (
    .a(\u2_Display/n5305 ),
    .b(1'b1),
    .c(\u2_Display/add162/c23 ),
    .o({\u2_Display/add162/c24 ,\u2_Display/n5331 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u24  (
    .a(\u2_Display/n5304 ),
    .b(1'b1),
    .c(\u2_Display/add162/c24 ),
    .o({\u2_Display/add162/c25 ,\u2_Display/n5331 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u25  (
    .a(\u2_Display/n5303 ),
    .b(1'b1),
    .c(\u2_Display/add162/c25 ),
    .o({\u2_Display/add162/c26 ,\u2_Display/n5331 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u26  (
    .a(\u2_Display/n5302 ),
    .b(1'b1),
    .c(\u2_Display/add162/c26 ),
    .o({\u2_Display/add162/c27 ,\u2_Display/n5331 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u27  (
    .a(\u2_Display/n5301 ),
    .b(1'b1),
    .c(\u2_Display/add162/c27 ),
    .o({\u2_Display/add162/c28 ,\u2_Display/n5331 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u28  (
    .a(\u2_Display/n5300 ),
    .b(1'b1),
    .c(\u2_Display/add162/c28 ),
    .o({\u2_Display/add162/c29 ,\u2_Display/n5331 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u29  (
    .a(\u2_Display/n5299 ),
    .b(1'b1),
    .c(\u2_Display/add162/c29 ),
    .o({\u2_Display/add162/c30 ,\u2_Display/n5331 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u3  (
    .a(\u2_Display/n5325 ),
    .b(1'b1),
    .c(\u2_Display/add162/c3 ),
    .o({\u2_Display/add162/c4 ,\u2_Display/n5331 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u30  (
    .a(\u2_Display/n5298 ),
    .b(1'b1),
    .c(\u2_Display/add162/c30 ),
    .o({\u2_Display/add162/c31 ,\u2_Display/n5331 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u31  (
    .a(\u2_Display/n5297 ),
    .b(1'b1),
    .c(\u2_Display/add162/c31 ),
    .o({open_n1047,\u2_Display/n5331 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u4  (
    .a(\u2_Display/n5324 ),
    .b(1'b1),
    .c(\u2_Display/add162/c4 ),
    .o({\u2_Display/add162/c5 ,\u2_Display/n5331 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u5  (
    .a(\u2_Display/n5323 ),
    .b(1'b1),
    .c(\u2_Display/add162/c5 ),
    .o({\u2_Display/add162/c6 ,\u2_Display/n5331 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u6  (
    .a(\u2_Display/n5322 ),
    .b(1'b1),
    .c(\u2_Display/add162/c6 ),
    .o({\u2_Display/add162/c7 ,\u2_Display/n5331 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u7  (
    .a(\u2_Display/n5321 ),
    .b(1'b1),
    .c(\u2_Display/add162/c7 ),
    .o({\u2_Display/add162/c8 ,\u2_Display/n5331 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u8  (
    .a(\u2_Display/n5320 ),
    .b(1'b1),
    .c(\u2_Display/add162/c8 ),
    .o({\u2_Display/add162/c9 ,\u2_Display/n5331 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add162/u9  (
    .a(\u2_Display/n5319 ),
    .b(1'b1),
    .c(\u2_Display/add162/c9 ),
    .o({\u2_Display/add162/c10 ,\u2_Display/n5331 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add162/ucin  (
    .a(1'b1),
    .o({\u2_Display/add162/c0 ,open_n1050}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u0  (
    .a(\u2_Display/n5363 ),
    .b(1'b1),
    .c(\u2_Display/add163/c0 ),
    .o({\u2_Display/add163/c1 ,\u2_Display/n5366 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u1  (
    .a(\u2_Display/n5362 ),
    .b(1'b1),
    .c(\u2_Display/add163/c1 ),
    .o({\u2_Display/add163/c2 ,\u2_Display/n5366 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u10  (
    .a(\u2_Display/n5353 ),
    .b(1'b1),
    .c(\u2_Display/add163/c10 ),
    .o({\u2_Display/add163/c11 ,\u2_Display/n5366 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u11  (
    .a(\u2_Display/n5352 ),
    .b(1'b1),
    .c(\u2_Display/add163/c11 ),
    .o({\u2_Display/add163/c12 ,\u2_Display/n5366 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u12  (
    .a(\u2_Display/n5351 ),
    .b(1'b1),
    .c(\u2_Display/add163/c12 ),
    .o({\u2_Display/add163/c13 ,\u2_Display/n5366 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u13  (
    .a(\u2_Display/n5350 ),
    .b(1'b1),
    .c(\u2_Display/add163/c13 ),
    .o({\u2_Display/add163/c14 ,\u2_Display/n5366 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u14  (
    .a(\u2_Display/n5349 ),
    .b(1'b1),
    .c(\u2_Display/add163/c14 ),
    .o({\u2_Display/add163/c15 ,\u2_Display/n5366 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u15  (
    .a(\u2_Display/n5348 ),
    .b(1'b1),
    .c(\u2_Display/add163/c15 ),
    .o({\u2_Display/add163/c16 ,\u2_Display/n5366 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u16  (
    .a(\u2_Display/n5347 ),
    .b(1'b0),
    .c(\u2_Display/add163/c16 ),
    .o({\u2_Display/add163/c17 ,\u2_Display/n5366 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u17  (
    .a(\u2_Display/n5346 ),
    .b(1'b1),
    .c(\u2_Display/add163/c17 ),
    .o({\u2_Display/add163/c18 ,\u2_Display/n5366 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u18  (
    .a(\u2_Display/n5345 ),
    .b(1'b0),
    .c(\u2_Display/add163/c18 ),
    .o({\u2_Display/add163/c19 ,\u2_Display/n5366 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u19  (
    .a(\u2_Display/n5344 ),
    .b(1'b1),
    .c(\u2_Display/add163/c19 ),
    .o({\u2_Display/add163/c20 ,\u2_Display/n5366 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u2  (
    .a(\u2_Display/n5361 ),
    .b(1'b1),
    .c(\u2_Display/add163/c2 ),
    .o({\u2_Display/add163/c3 ,\u2_Display/n5366 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u20  (
    .a(\u2_Display/n5343 ),
    .b(1'b1),
    .c(\u2_Display/add163/c20 ),
    .o({\u2_Display/add163/c21 ,\u2_Display/n5366 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u21  (
    .a(\u2_Display/n5342 ),
    .b(1'b1),
    .c(\u2_Display/add163/c21 ),
    .o({\u2_Display/add163/c22 ,\u2_Display/n5366 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u22  (
    .a(\u2_Display/n5341 ),
    .b(1'b1),
    .c(\u2_Display/add163/c22 ),
    .o({\u2_Display/add163/c23 ,\u2_Display/n5366 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u23  (
    .a(\u2_Display/n5340 ),
    .b(1'b1),
    .c(\u2_Display/add163/c23 ),
    .o({\u2_Display/add163/c24 ,\u2_Display/n5366 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u24  (
    .a(\u2_Display/n5339 ),
    .b(1'b1),
    .c(\u2_Display/add163/c24 ),
    .o({\u2_Display/add163/c25 ,\u2_Display/n5366 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u25  (
    .a(\u2_Display/n5338 ),
    .b(1'b1),
    .c(\u2_Display/add163/c25 ),
    .o({\u2_Display/add163/c26 ,\u2_Display/n5366 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u26  (
    .a(\u2_Display/n5337 ),
    .b(1'b1),
    .c(\u2_Display/add163/c26 ),
    .o({\u2_Display/add163/c27 ,\u2_Display/n5366 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u27  (
    .a(\u2_Display/n5336 ),
    .b(1'b1),
    .c(\u2_Display/add163/c27 ),
    .o({\u2_Display/add163/c28 ,\u2_Display/n5366 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u28  (
    .a(\u2_Display/n5335 ),
    .b(1'b1),
    .c(\u2_Display/add163/c28 ),
    .o({\u2_Display/add163/c29 ,\u2_Display/n5366 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u29  (
    .a(\u2_Display/n5334 ),
    .b(1'b1),
    .c(\u2_Display/add163/c29 ),
    .o({\u2_Display/add163/c30 ,\u2_Display/n5366 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u3  (
    .a(\u2_Display/n5360 ),
    .b(1'b1),
    .c(\u2_Display/add163/c3 ),
    .o({\u2_Display/add163/c4 ,\u2_Display/n5366 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u30  (
    .a(\u2_Display/n5333 ),
    .b(1'b1),
    .c(\u2_Display/add163/c30 ),
    .o({\u2_Display/add163/c31 ,\u2_Display/n5366 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u31  (
    .a(\u2_Display/n5332 ),
    .b(1'b1),
    .c(\u2_Display/add163/c31 ),
    .o({open_n1051,\u2_Display/n5366 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u4  (
    .a(\u2_Display/n5359 ),
    .b(1'b1),
    .c(\u2_Display/add163/c4 ),
    .o({\u2_Display/add163/c5 ,\u2_Display/n5366 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u5  (
    .a(\u2_Display/n5358 ),
    .b(1'b1),
    .c(\u2_Display/add163/c5 ),
    .o({\u2_Display/add163/c6 ,\u2_Display/n5366 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u6  (
    .a(\u2_Display/n5357 ),
    .b(1'b1),
    .c(\u2_Display/add163/c6 ),
    .o({\u2_Display/add163/c7 ,\u2_Display/n5366 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u7  (
    .a(\u2_Display/n5356 ),
    .b(1'b1),
    .c(\u2_Display/add163/c7 ),
    .o({\u2_Display/add163/c8 ,\u2_Display/n5366 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u8  (
    .a(\u2_Display/n5355 ),
    .b(1'b1),
    .c(\u2_Display/add163/c8 ),
    .o({\u2_Display/add163/c9 ,\u2_Display/n5366 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add163/u9  (
    .a(\u2_Display/n5354 ),
    .b(1'b1),
    .c(\u2_Display/add163/c9 ),
    .o({\u2_Display/add163/c10 ,\u2_Display/n5366 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add163/ucin  (
    .a(1'b1),
    .o({\u2_Display/add163/c0 ,open_n1054}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u0  (
    .a(\u2_Display/n5398 ),
    .b(1'b1),
    .c(\u2_Display/add164/c0 ),
    .o({\u2_Display/add164/c1 ,\u2_Display/n5401 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u1  (
    .a(\u2_Display/n5397 ),
    .b(1'b1),
    .c(\u2_Display/add164/c1 ),
    .o({\u2_Display/add164/c2 ,\u2_Display/n5401 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u10  (
    .a(\u2_Display/n5388 ),
    .b(1'b1),
    .c(\u2_Display/add164/c10 ),
    .o({\u2_Display/add164/c11 ,\u2_Display/n5401 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u11  (
    .a(\u2_Display/n5387 ),
    .b(1'b1),
    .c(\u2_Display/add164/c11 ),
    .o({\u2_Display/add164/c12 ,\u2_Display/n5401 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u12  (
    .a(\u2_Display/n5386 ),
    .b(1'b1),
    .c(\u2_Display/add164/c12 ),
    .o({\u2_Display/add164/c13 ,\u2_Display/n5401 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u13  (
    .a(\u2_Display/n5385 ),
    .b(1'b1),
    .c(\u2_Display/add164/c13 ),
    .o({\u2_Display/add164/c14 ,\u2_Display/n5401 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u14  (
    .a(\u2_Display/n5384 ),
    .b(1'b1),
    .c(\u2_Display/add164/c14 ),
    .o({\u2_Display/add164/c15 ,\u2_Display/n5401 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u15  (
    .a(\u2_Display/n5383 ),
    .b(1'b0),
    .c(\u2_Display/add164/c15 ),
    .o({\u2_Display/add164/c16 ,\u2_Display/n5401 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u16  (
    .a(\u2_Display/n5382 ),
    .b(1'b1),
    .c(\u2_Display/add164/c16 ),
    .o({\u2_Display/add164/c17 ,\u2_Display/n5401 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u17  (
    .a(\u2_Display/n5381 ),
    .b(1'b0),
    .c(\u2_Display/add164/c17 ),
    .o({\u2_Display/add164/c18 ,\u2_Display/n5401 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u18  (
    .a(\u2_Display/n5380 ),
    .b(1'b1),
    .c(\u2_Display/add164/c18 ),
    .o({\u2_Display/add164/c19 ,\u2_Display/n5401 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u19  (
    .a(\u2_Display/n5379 ),
    .b(1'b1),
    .c(\u2_Display/add164/c19 ),
    .o({\u2_Display/add164/c20 ,\u2_Display/n5401 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u2  (
    .a(\u2_Display/n5396 ),
    .b(1'b1),
    .c(\u2_Display/add164/c2 ),
    .o({\u2_Display/add164/c3 ,\u2_Display/n5401 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u20  (
    .a(\u2_Display/n5378 ),
    .b(1'b1),
    .c(\u2_Display/add164/c20 ),
    .o({\u2_Display/add164/c21 ,\u2_Display/n5401 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u21  (
    .a(\u2_Display/n5377 ),
    .b(1'b1),
    .c(\u2_Display/add164/c21 ),
    .o({\u2_Display/add164/c22 ,\u2_Display/n5401 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u22  (
    .a(\u2_Display/n5376 ),
    .b(1'b1),
    .c(\u2_Display/add164/c22 ),
    .o({\u2_Display/add164/c23 ,\u2_Display/n5401 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u23  (
    .a(\u2_Display/n5375 ),
    .b(1'b1),
    .c(\u2_Display/add164/c23 ),
    .o({\u2_Display/add164/c24 ,\u2_Display/n5401 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u24  (
    .a(\u2_Display/n5374 ),
    .b(1'b1),
    .c(\u2_Display/add164/c24 ),
    .o({\u2_Display/add164/c25 ,\u2_Display/n5401 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u25  (
    .a(\u2_Display/n5373 ),
    .b(1'b1),
    .c(\u2_Display/add164/c25 ),
    .o({\u2_Display/add164/c26 ,\u2_Display/n5401 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u26  (
    .a(\u2_Display/n5372 ),
    .b(1'b1),
    .c(\u2_Display/add164/c26 ),
    .o({\u2_Display/add164/c27 ,\u2_Display/n5401 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u27  (
    .a(\u2_Display/n5371 ),
    .b(1'b1),
    .c(\u2_Display/add164/c27 ),
    .o({\u2_Display/add164/c28 ,\u2_Display/n5401 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u28  (
    .a(\u2_Display/n5370 ),
    .b(1'b1),
    .c(\u2_Display/add164/c28 ),
    .o({\u2_Display/add164/c29 ,\u2_Display/n5401 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u29  (
    .a(\u2_Display/n5369 ),
    .b(1'b1),
    .c(\u2_Display/add164/c29 ),
    .o({\u2_Display/add164/c30 ,\u2_Display/n5401 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u3  (
    .a(\u2_Display/n5395 ),
    .b(1'b1),
    .c(\u2_Display/add164/c3 ),
    .o({\u2_Display/add164/c4 ,\u2_Display/n5401 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u30  (
    .a(\u2_Display/n5368 ),
    .b(1'b1),
    .c(\u2_Display/add164/c30 ),
    .o({\u2_Display/add164/c31 ,\u2_Display/n5401 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u31  (
    .a(\u2_Display/n5367 ),
    .b(1'b1),
    .c(\u2_Display/add164/c31 ),
    .o({open_n1055,\u2_Display/n5401 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u4  (
    .a(\u2_Display/n5394 ),
    .b(1'b1),
    .c(\u2_Display/add164/c4 ),
    .o({\u2_Display/add164/c5 ,\u2_Display/n5401 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u5  (
    .a(\u2_Display/n5393 ),
    .b(1'b1),
    .c(\u2_Display/add164/c5 ),
    .o({\u2_Display/add164/c6 ,\u2_Display/n5401 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u6  (
    .a(\u2_Display/n5392 ),
    .b(1'b1),
    .c(\u2_Display/add164/c6 ),
    .o({\u2_Display/add164/c7 ,\u2_Display/n5401 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u7  (
    .a(\u2_Display/n5391 ),
    .b(1'b1),
    .c(\u2_Display/add164/c7 ),
    .o({\u2_Display/add164/c8 ,\u2_Display/n5401 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u8  (
    .a(\u2_Display/n5390 ),
    .b(1'b1),
    .c(\u2_Display/add164/c8 ),
    .o({\u2_Display/add164/c9 ,\u2_Display/n5401 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add164/u9  (
    .a(\u2_Display/n5389 ),
    .b(1'b1),
    .c(\u2_Display/add164/c9 ),
    .o({\u2_Display/add164/c10 ,\u2_Display/n5401 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add164/ucin  (
    .a(1'b1),
    .o({\u2_Display/add164/c0 ,open_n1058}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u0  (
    .a(\u2_Display/n5433 ),
    .b(1'b1),
    .c(\u2_Display/add165/c0 ),
    .o({\u2_Display/add165/c1 ,\u2_Display/n5436 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u1  (
    .a(\u2_Display/n5432 ),
    .b(1'b1),
    .c(\u2_Display/add165/c1 ),
    .o({\u2_Display/add165/c2 ,\u2_Display/n5436 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u10  (
    .a(\u2_Display/n5423 ),
    .b(1'b1),
    .c(\u2_Display/add165/c10 ),
    .o({\u2_Display/add165/c11 ,\u2_Display/n5436 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u11  (
    .a(\u2_Display/n5422 ),
    .b(1'b1),
    .c(\u2_Display/add165/c11 ),
    .o({\u2_Display/add165/c12 ,\u2_Display/n5436 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u12  (
    .a(\u2_Display/n5421 ),
    .b(1'b1),
    .c(\u2_Display/add165/c12 ),
    .o({\u2_Display/add165/c13 ,\u2_Display/n5436 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u13  (
    .a(\u2_Display/n5420 ),
    .b(1'b1),
    .c(\u2_Display/add165/c13 ),
    .o({\u2_Display/add165/c14 ,\u2_Display/n5436 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u14  (
    .a(\u2_Display/n5419 ),
    .b(1'b0),
    .c(\u2_Display/add165/c14 ),
    .o({\u2_Display/add165/c15 ,\u2_Display/n5436 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u15  (
    .a(\u2_Display/n5418 ),
    .b(1'b1),
    .c(\u2_Display/add165/c15 ),
    .o({\u2_Display/add165/c16 ,\u2_Display/n5436 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u16  (
    .a(\u2_Display/n5417 ),
    .b(1'b0),
    .c(\u2_Display/add165/c16 ),
    .o({\u2_Display/add165/c17 ,\u2_Display/n5436 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u17  (
    .a(\u2_Display/n5416 ),
    .b(1'b1),
    .c(\u2_Display/add165/c17 ),
    .o({\u2_Display/add165/c18 ,\u2_Display/n5436 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u18  (
    .a(\u2_Display/n5415 ),
    .b(1'b1),
    .c(\u2_Display/add165/c18 ),
    .o({\u2_Display/add165/c19 ,\u2_Display/n5436 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u19  (
    .a(\u2_Display/n5414 ),
    .b(1'b1),
    .c(\u2_Display/add165/c19 ),
    .o({\u2_Display/add165/c20 ,\u2_Display/n5436 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u2  (
    .a(\u2_Display/n5431 ),
    .b(1'b1),
    .c(\u2_Display/add165/c2 ),
    .o({\u2_Display/add165/c3 ,\u2_Display/n5436 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u20  (
    .a(\u2_Display/n5413 ),
    .b(1'b1),
    .c(\u2_Display/add165/c20 ),
    .o({\u2_Display/add165/c21 ,\u2_Display/n5436 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u21  (
    .a(\u2_Display/n5412 ),
    .b(1'b1),
    .c(\u2_Display/add165/c21 ),
    .o({\u2_Display/add165/c22 ,\u2_Display/n5436 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u22  (
    .a(\u2_Display/n5411 ),
    .b(1'b1),
    .c(\u2_Display/add165/c22 ),
    .o({\u2_Display/add165/c23 ,\u2_Display/n5436 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u23  (
    .a(\u2_Display/n5410 ),
    .b(1'b1),
    .c(\u2_Display/add165/c23 ),
    .o({\u2_Display/add165/c24 ,\u2_Display/n5436 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u24  (
    .a(\u2_Display/n5409 ),
    .b(1'b1),
    .c(\u2_Display/add165/c24 ),
    .o({\u2_Display/add165/c25 ,\u2_Display/n5436 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u25  (
    .a(\u2_Display/n5408 ),
    .b(1'b1),
    .c(\u2_Display/add165/c25 ),
    .o({\u2_Display/add165/c26 ,\u2_Display/n5436 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u26  (
    .a(\u2_Display/n5407 ),
    .b(1'b1),
    .c(\u2_Display/add165/c26 ),
    .o({\u2_Display/add165/c27 ,\u2_Display/n5436 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u27  (
    .a(\u2_Display/n5406 ),
    .b(1'b1),
    .c(\u2_Display/add165/c27 ),
    .o({\u2_Display/add165/c28 ,\u2_Display/n5436 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u28  (
    .a(\u2_Display/n5405 ),
    .b(1'b1),
    .c(\u2_Display/add165/c28 ),
    .o({\u2_Display/add165/c29 ,\u2_Display/n5436 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u29  (
    .a(\u2_Display/n5404 ),
    .b(1'b1),
    .c(\u2_Display/add165/c29 ),
    .o({\u2_Display/add165/c30 ,\u2_Display/n5436 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u3  (
    .a(\u2_Display/n5430 ),
    .b(1'b1),
    .c(\u2_Display/add165/c3 ),
    .o({\u2_Display/add165/c4 ,\u2_Display/n5436 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u30  (
    .a(\u2_Display/n5403 ),
    .b(1'b1),
    .c(\u2_Display/add165/c30 ),
    .o({\u2_Display/add165/c31 ,\u2_Display/n5436 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u31  (
    .a(\u2_Display/n5402 ),
    .b(1'b1),
    .c(\u2_Display/add165/c31 ),
    .o({open_n1059,\u2_Display/n5436 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u4  (
    .a(\u2_Display/n5429 ),
    .b(1'b1),
    .c(\u2_Display/add165/c4 ),
    .o({\u2_Display/add165/c5 ,\u2_Display/n5436 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u5  (
    .a(\u2_Display/n5428 ),
    .b(1'b1),
    .c(\u2_Display/add165/c5 ),
    .o({\u2_Display/add165/c6 ,\u2_Display/n5436 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u6  (
    .a(\u2_Display/n5427 ),
    .b(1'b1),
    .c(\u2_Display/add165/c6 ),
    .o({\u2_Display/add165/c7 ,\u2_Display/n5436 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u7  (
    .a(\u2_Display/n5426 ),
    .b(1'b1),
    .c(\u2_Display/add165/c7 ),
    .o({\u2_Display/add165/c8 ,\u2_Display/n5436 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u8  (
    .a(\u2_Display/n5425 ),
    .b(1'b1),
    .c(\u2_Display/add165/c8 ),
    .o({\u2_Display/add165/c9 ,\u2_Display/n5436 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add165/u9  (
    .a(\u2_Display/n5424 ),
    .b(1'b1),
    .c(\u2_Display/add165/c9 ),
    .o({\u2_Display/add165/c10 ,\u2_Display/n5436 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add165/ucin  (
    .a(1'b1),
    .o({\u2_Display/add165/c0 ,open_n1062}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u0  (
    .a(\u2_Display/n5468 ),
    .b(1'b1),
    .c(\u2_Display/add166/c0 ),
    .o({\u2_Display/add166/c1 ,\u2_Display/n5471 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u1  (
    .a(\u2_Display/n5467 ),
    .b(1'b1),
    .c(\u2_Display/add166/c1 ),
    .o({\u2_Display/add166/c2 ,\u2_Display/n5471 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u10  (
    .a(\u2_Display/n5458 ),
    .b(1'b1),
    .c(\u2_Display/add166/c10 ),
    .o({\u2_Display/add166/c11 ,\u2_Display/n5471 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u11  (
    .a(\u2_Display/n5457 ),
    .b(1'b1),
    .c(\u2_Display/add166/c11 ),
    .o({\u2_Display/add166/c12 ,\u2_Display/n5471 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u12  (
    .a(\u2_Display/n5456 ),
    .b(1'b1),
    .c(\u2_Display/add166/c12 ),
    .o({\u2_Display/add166/c13 ,\u2_Display/n5471 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u13  (
    .a(\u2_Display/n5455 ),
    .b(1'b0),
    .c(\u2_Display/add166/c13 ),
    .o({\u2_Display/add166/c14 ,\u2_Display/n5471 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u14  (
    .a(\u2_Display/n5454 ),
    .b(1'b1),
    .c(\u2_Display/add166/c14 ),
    .o({\u2_Display/add166/c15 ,\u2_Display/n5471 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u15  (
    .a(\u2_Display/n5453 ),
    .b(1'b0),
    .c(\u2_Display/add166/c15 ),
    .o({\u2_Display/add166/c16 ,\u2_Display/n5471 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u16  (
    .a(\u2_Display/n5452 ),
    .b(1'b1),
    .c(\u2_Display/add166/c16 ),
    .o({\u2_Display/add166/c17 ,\u2_Display/n5471 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u17  (
    .a(\u2_Display/n5451 ),
    .b(1'b1),
    .c(\u2_Display/add166/c17 ),
    .o({\u2_Display/add166/c18 ,\u2_Display/n5471 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u18  (
    .a(\u2_Display/n5450 ),
    .b(1'b1),
    .c(\u2_Display/add166/c18 ),
    .o({\u2_Display/add166/c19 ,\u2_Display/n5471 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u19  (
    .a(\u2_Display/n5449 ),
    .b(1'b1),
    .c(\u2_Display/add166/c19 ),
    .o({\u2_Display/add166/c20 ,\u2_Display/n5471 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u2  (
    .a(\u2_Display/n5466 ),
    .b(1'b1),
    .c(\u2_Display/add166/c2 ),
    .o({\u2_Display/add166/c3 ,\u2_Display/n5471 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u20  (
    .a(\u2_Display/n5448 ),
    .b(1'b1),
    .c(\u2_Display/add166/c20 ),
    .o({\u2_Display/add166/c21 ,\u2_Display/n5471 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u21  (
    .a(\u2_Display/n5447 ),
    .b(1'b1),
    .c(\u2_Display/add166/c21 ),
    .o({\u2_Display/add166/c22 ,\u2_Display/n5471 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u22  (
    .a(\u2_Display/n5446 ),
    .b(1'b1),
    .c(\u2_Display/add166/c22 ),
    .o({\u2_Display/add166/c23 ,\u2_Display/n5471 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u23  (
    .a(\u2_Display/n5445 ),
    .b(1'b1),
    .c(\u2_Display/add166/c23 ),
    .o({\u2_Display/add166/c24 ,\u2_Display/n5471 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u24  (
    .a(\u2_Display/n5444 ),
    .b(1'b1),
    .c(\u2_Display/add166/c24 ),
    .o({\u2_Display/add166/c25 ,\u2_Display/n5471 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u25  (
    .a(\u2_Display/n5443 ),
    .b(1'b1),
    .c(\u2_Display/add166/c25 ),
    .o({\u2_Display/add166/c26 ,\u2_Display/n5471 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u26  (
    .a(\u2_Display/n5442 ),
    .b(1'b1),
    .c(\u2_Display/add166/c26 ),
    .o({\u2_Display/add166/c27 ,\u2_Display/n5471 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u27  (
    .a(\u2_Display/n5441 ),
    .b(1'b1),
    .c(\u2_Display/add166/c27 ),
    .o({\u2_Display/add166/c28 ,\u2_Display/n5471 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u28  (
    .a(\u2_Display/n5440 ),
    .b(1'b1),
    .c(\u2_Display/add166/c28 ),
    .o({\u2_Display/add166/c29 ,\u2_Display/n5471 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u29  (
    .a(\u2_Display/n5439 ),
    .b(1'b1),
    .c(\u2_Display/add166/c29 ),
    .o({\u2_Display/add166/c30 ,\u2_Display/n5471 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u3  (
    .a(\u2_Display/n5465 ),
    .b(1'b1),
    .c(\u2_Display/add166/c3 ),
    .o({\u2_Display/add166/c4 ,\u2_Display/n5471 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u30  (
    .a(\u2_Display/n5438 ),
    .b(1'b1),
    .c(\u2_Display/add166/c30 ),
    .o({\u2_Display/add166/c31 ,\u2_Display/n5471 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u31  (
    .a(\u2_Display/n5437 ),
    .b(1'b1),
    .c(\u2_Display/add166/c31 ),
    .o({open_n1063,\u2_Display/n5471 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u4  (
    .a(\u2_Display/n5464 ),
    .b(1'b1),
    .c(\u2_Display/add166/c4 ),
    .o({\u2_Display/add166/c5 ,\u2_Display/n5471 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u5  (
    .a(\u2_Display/n5463 ),
    .b(1'b1),
    .c(\u2_Display/add166/c5 ),
    .o({\u2_Display/add166/c6 ,\u2_Display/n5471 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u6  (
    .a(\u2_Display/n5462 ),
    .b(1'b1),
    .c(\u2_Display/add166/c6 ),
    .o({\u2_Display/add166/c7 ,\u2_Display/n5471 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u7  (
    .a(\u2_Display/n5461 ),
    .b(1'b1),
    .c(\u2_Display/add166/c7 ),
    .o({\u2_Display/add166/c8 ,\u2_Display/n5471 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u8  (
    .a(\u2_Display/n5460 ),
    .b(1'b1),
    .c(\u2_Display/add166/c8 ),
    .o({\u2_Display/add166/c9 ,\u2_Display/n5471 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add166/u9  (
    .a(\u2_Display/n5459 ),
    .b(1'b1),
    .c(\u2_Display/add166/c9 ),
    .o({\u2_Display/add166/c10 ,\u2_Display/n5471 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add166/ucin  (
    .a(1'b1),
    .o({\u2_Display/add166/c0 ,open_n1066}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u0  (
    .a(\u2_Display/n5503 ),
    .b(1'b1),
    .c(\u2_Display/add167/c0 ),
    .o({\u2_Display/add167/c1 ,\u2_Display/n5506 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u1  (
    .a(\u2_Display/n5502 ),
    .b(1'b1),
    .c(\u2_Display/add167/c1 ),
    .o({\u2_Display/add167/c2 ,\u2_Display/n5506 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u10  (
    .a(\u2_Display/n5493 ),
    .b(1'b1),
    .c(\u2_Display/add167/c10 ),
    .o({\u2_Display/add167/c11 ,\u2_Display/n5506 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u11  (
    .a(\u2_Display/n5492 ),
    .b(1'b1),
    .c(\u2_Display/add167/c11 ),
    .o({\u2_Display/add167/c12 ,\u2_Display/n5506 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u12  (
    .a(\u2_Display/n5491 ),
    .b(1'b0),
    .c(\u2_Display/add167/c12 ),
    .o({\u2_Display/add167/c13 ,\u2_Display/n5506 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u13  (
    .a(\u2_Display/n5490 ),
    .b(1'b1),
    .c(\u2_Display/add167/c13 ),
    .o({\u2_Display/add167/c14 ,\u2_Display/n5506 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u14  (
    .a(\u2_Display/n5489 ),
    .b(1'b0),
    .c(\u2_Display/add167/c14 ),
    .o({\u2_Display/add167/c15 ,\u2_Display/n5506 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u15  (
    .a(\u2_Display/n5488 ),
    .b(1'b1),
    .c(\u2_Display/add167/c15 ),
    .o({\u2_Display/add167/c16 ,\u2_Display/n5506 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u16  (
    .a(\u2_Display/n5487 ),
    .b(1'b1),
    .c(\u2_Display/add167/c16 ),
    .o({\u2_Display/add167/c17 ,\u2_Display/n5506 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u17  (
    .a(\u2_Display/n5486 ),
    .b(1'b1),
    .c(\u2_Display/add167/c17 ),
    .o({\u2_Display/add167/c18 ,\u2_Display/n5506 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u18  (
    .a(\u2_Display/n5485 ),
    .b(1'b1),
    .c(\u2_Display/add167/c18 ),
    .o({\u2_Display/add167/c19 ,\u2_Display/n5506 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u19  (
    .a(\u2_Display/n5484 ),
    .b(1'b1),
    .c(\u2_Display/add167/c19 ),
    .o({\u2_Display/add167/c20 ,\u2_Display/n5506 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u2  (
    .a(\u2_Display/n5501 ),
    .b(1'b1),
    .c(\u2_Display/add167/c2 ),
    .o({\u2_Display/add167/c3 ,\u2_Display/n5506 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u20  (
    .a(\u2_Display/n5483 ),
    .b(1'b1),
    .c(\u2_Display/add167/c20 ),
    .o({\u2_Display/add167/c21 ,\u2_Display/n5506 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u21  (
    .a(\u2_Display/n5482 ),
    .b(1'b1),
    .c(\u2_Display/add167/c21 ),
    .o({\u2_Display/add167/c22 ,\u2_Display/n5506 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u22  (
    .a(\u2_Display/n5481 ),
    .b(1'b1),
    .c(\u2_Display/add167/c22 ),
    .o({\u2_Display/add167/c23 ,\u2_Display/n5506 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u23  (
    .a(\u2_Display/n5480 ),
    .b(1'b1),
    .c(\u2_Display/add167/c23 ),
    .o({\u2_Display/add167/c24 ,\u2_Display/n5506 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u24  (
    .a(\u2_Display/n5479 ),
    .b(1'b1),
    .c(\u2_Display/add167/c24 ),
    .o({\u2_Display/add167/c25 ,\u2_Display/n5506 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u25  (
    .a(\u2_Display/n5478 ),
    .b(1'b1),
    .c(\u2_Display/add167/c25 ),
    .o({\u2_Display/add167/c26 ,\u2_Display/n5506 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u26  (
    .a(\u2_Display/n5477 ),
    .b(1'b1),
    .c(\u2_Display/add167/c26 ),
    .o({\u2_Display/add167/c27 ,\u2_Display/n5506 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u27  (
    .a(\u2_Display/n5476 ),
    .b(1'b1),
    .c(\u2_Display/add167/c27 ),
    .o({\u2_Display/add167/c28 ,\u2_Display/n5506 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u28  (
    .a(\u2_Display/n5475 ),
    .b(1'b1),
    .c(\u2_Display/add167/c28 ),
    .o({\u2_Display/add167/c29 ,\u2_Display/n5506 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u29  (
    .a(\u2_Display/n5474 ),
    .b(1'b1),
    .c(\u2_Display/add167/c29 ),
    .o({\u2_Display/add167/c30 ,\u2_Display/n5506 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u3  (
    .a(\u2_Display/n5500 ),
    .b(1'b1),
    .c(\u2_Display/add167/c3 ),
    .o({\u2_Display/add167/c4 ,\u2_Display/n5506 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u30  (
    .a(\u2_Display/n5473 ),
    .b(1'b1),
    .c(\u2_Display/add167/c30 ),
    .o({\u2_Display/add167/c31 ,\u2_Display/n5506 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u31  (
    .a(\u2_Display/n5472 ),
    .b(1'b1),
    .c(\u2_Display/add167/c31 ),
    .o({open_n1067,\u2_Display/n5506 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u4  (
    .a(\u2_Display/n5499 ),
    .b(1'b1),
    .c(\u2_Display/add167/c4 ),
    .o({\u2_Display/add167/c5 ,\u2_Display/n5506 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u5  (
    .a(\u2_Display/n5498 ),
    .b(1'b1),
    .c(\u2_Display/add167/c5 ),
    .o({\u2_Display/add167/c6 ,\u2_Display/n5506 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u6  (
    .a(\u2_Display/n5497 ),
    .b(1'b1),
    .c(\u2_Display/add167/c6 ),
    .o({\u2_Display/add167/c7 ,\u2_Display/n5506 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u7  (
    .a(\u2_Display/n5496 ),
    .b(1'b1),
    .c(\u2_Display/add167/c7 ),
    .o({\u2_Display/add167/c8 ,\u2_Display/n5506 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u8  (
    .a(\u2_Display/n5495 ),
    .b(1'b1),
    .c(\u2_Display/add167/c8 ),
    .o({\u2_Display/add167/c9 ,\u2_Display/n5506 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add167/u9  (
    .a(\u2_Display/n5494 ),
    .b(1'b1),
    .c(\u2_Display/add167/c9 ),
    .o({\u2_Display/add167/c10 ,\u2_Display/n5506 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add167/ucin  (
    .a(1'b1),
    .o({\u2_Display/add167/c0 ,open_n1070}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u0  (
    .a(\u2_Display/n5538 ),
    .b(1'b1),
    .c(\u2_Display/add168/c0 ),
    .o({\u2_Display/add168/c1 ,\u2_Display/n5541 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u1  (
    .a(\u2_Display/n5537 ),
    .b(1'b1),
    .c(\u2_Display/add168/c1 ),
    .o({\u2_Display/add168/c2 ,\u2_Display/n5541 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u10  (
    .a(\u2_Display/n5528 ),
    .b(1'b1),
    .c(\u2_Display/add168/c10 ),
    .o({\u2_Display/add168/c11 ,\u2_Display/n5541 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u11  (
    .a(\u2_Display/n5527 ),
    .b(1'b0),
    .c(\u2_Display/add168/c11 ),
    .o({\u2_Display/add168/c12 ,\u2_Display/n5541 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u12  (
    .a(\u2_Display/n5526 ),
    .b(1'b1),
    .c(\u2_Display/add168/c12 ),
    .o({\u2_Display/add168/c13 ,\u2_Display/n5541 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u13  (
    .a(\u2_Display/n5525 ),
    .b(1'b0),
    .c(\u2_Display/add168/c13 ),
    .o({\u2_Display/add168/c14 ,\u2_Display/n5541 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u14  (
    .a(\u2_Display/n5524 ),
    .b(1'b1),
    .c(\u2_Display/add168/c14 ),
    .o({\u2_Display/add168/c15 ,\u2_Display/n5541 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u15  (
    .a(\u2_Display/n5523 ),
    .b(1'b1),
    .c(\u2_Display/add168/c15 ),
    .o({\u2_Display/add168/c16 ,\u2_Display/n5541 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u16  (
    .a(\u2_Display/n5522 ),
    .b(1'b1),
    .c(\u2_Display/add168/c16 ),
    .o({\u2_Display/add168/c17 ,\u2_Display/n5541 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u17  (
    .a(\u2_Display/n5521 ),
    .b(1'b1),
    .c(\u2_Display/add168/c17 ),
    .o({\u2_Display/add168/c18 ,\u2_Display/n5541 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u18  (
    .a(\u2_Display/n5520 ),
    .b(1'b1),
    .c(\u2_Display/add168/c18 ),
    .o({\u2_Display/add168/c19 ,\u2_Display/n5541 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u19  (
    .a(\u2_Display/n5519 ),
    .b(1'b1),
    .c(\u2_Display/add168/c19 ),
    .o({\u2_Display/add168/c20 ,\u2_Display/n5541 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u2  (
    .a(\u2_Display/n5536 ),
    .b(1'b1),
    .c(\u2_Display/add168/c2 ),
    .o({\u2_Display/add168/c3 ,\u2_Display/n5541 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u20  (
    .a(\u2_Display/n5518 ),
    .b(1'b1),
    .c(\u2_Display/add168/c20 ),
    .o({\u2_Display/add168/c21 ,\u2_Display/n5541 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u21  (
    .a(\u2_Display/n5517 ),
    .b(1'b1),
    .c(\u2_Display/add168/c21 ),
    .o({\u2_Display/add168/c22 ,\u2_Display/n5541 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u22  (
    .a(\u2_Display/n5516 ),
    .b(1'b1),
    .c(\u2_Display/add168/c22 ),
    .o({\u2_Display/add168/c23 ,\u2_Display/n5541 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u23  (
    .a(\u2_Display/n5515 ),
    .b(1'b1),
    .c(\u2_Display/add168/c23 ),
    .o({\u2_Display/add168/c24 ,\u2_Display/n5541 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u24  (
    .a(\u2_Display/n5514 ),
    .b(1'b1),
    .c(\u2_Display/add168/c24 ),
    .o({\u2_Display/add168/c25 ,\u2_Display/n5541 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u25  (
    .a(\u2_Display/n5513 ),
    .b(1'b1),
    .c(\u2_Display/add168/c25 ),
    .o({\u2_Display/add168/c26 ,\u2_Display/n5541 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u26  (
    .a(\u2_Display/n5512 ),
    .b(1'b1),
    .c(\u2_Display/add168/c26 ),
    .o({\u2_Display/add168/c27 ,\u2_Display/n5541 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u27  (
    .a(\u2_Display/n5511 ),
    .b(1'b1),
    .c(\u2_Display/add168/c27 ),
    .o({\u2_Display/add168/c28 ,\u2_Display/n5541 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u28  (
    .a(\u2_Display/n5510 ),
    .b(1'b1),
    .c(\u2_Display/add168/c28 ),
    .o({\u2_Display/add168/c29 ,\u2_Display/n5541 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u29  (
    .a(\u2_Display/n5509 ),
    .b(1'b1),
    .c(\u2_Display/add168/c29 ),
    .o({\u2_Display/add168/c30 ,\u2_Display/n5541 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u3  (
    .a(\u2_Display/n5535 ),
    .b(1'b1),
    .c(\u2_Display/add168/c3 ),
    .o({\u2_Display/add168/c4 ,\u2_Display/n5541 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u30  (
    .a(\u2_Display/n5508 ),
    .b(1'b1),
    .c(\u2_Display/add168/c30 ),
    .o({\u2_Display/add168/c31 ,\u2_Display/n5541 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u31  (
    .a(\u2_Display/n5507 ),
    .b(1'b1),
    .c(\u2_Display/add168/c31 ),
    .o({open_n1071,\u2_Display/n5541 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u4  (
    .a(\u2_Display/n5534 ),
    .b(1'b1),
    .c(\u2_Display/add168/c4 ),
    .o({\u2_Display/add168/c5 ,\u2_Display/n5541 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u5  (
    .a(\u2_Display/n5533 ),
    .b(1'b1),
    .c(\u2_Display/add168/c5 ),
    .o({\u2_Display/add168/c6 ,\u2_Display/n5541 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u6  (
    .a(\u2_Display/n5532 ),
    .b(1'b1),
    .c(\u2_Display/add168/c6 ),
    .o({\u2_Display/add168/c7 ,\u2_Display/n5541 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u7  (
    .a(\u2_Display/n5531 ),
    .b(1'b1),
    .c(\u2_Display/add168/c7 ),
    .o({\u2_Display/add168/c8 ,\u2_Display/n5541 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u8  (
    .a(\u2_Display/n5530 ),
    .b(1'b1),
    .c(\u2_Display/add168/c8 ),
    .o({\u2_Display/add168/c9 ,\u2_Display/n5541 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add168/u9  (
    .a(\u2_Display/n5529 ),
    .b(1'b1),
    .c(\u2_Display/add168/c9 ),
    .o({\u2_Display/add168/c10 ,\u2_Display/n5541 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add168/ucin  (
    .a(1'b1),
    .o({\u2_Display/add168/c0 ,open_n1074}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u0  (
    .a(\u2_Display/n5573 ),
    .b(1'b1),
    .c(\u2_Display/add169/c0 ),
    .o({\u2_Display/add169/c1 ,\u2_Display/n5576 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u1  (
    .a(\u2_Display/n5572 ),
    .b(1'b1),
    .c(\u2_Display/add169/c1 ),
    .o({\u2_Display/add169/c2 ,\u2_Display/n5576 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u10  (
    .a(\u2_Display/n5563 ),
    .b(1'b0),
    .c(\u2_Display/add169/c10 ),
    .o({\u2_Display/add169/c11 ,\u2_Display/n5576 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u11  (
    .a(\u2_Display/n5562 ),
    .b(1'b1),
    .c(\u2_Display/add169/c11 ),
    .o({\u2_Display/add169/c12 ,\u2_Display/n5576 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u12  (
    .a(\u2_Display/n5561 ),
    .b(1'b0),
    .c(\u2_Display/add169/c12 ),
    .o({\u2_Display/add169/c13 ,\u2_Display/n5576 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u13  (
    .a(\u2_Display/n5560 ),
    .b(1'b1),
    .c(\u2_Display/add169/c13 ),
    .o({\u2_Display/add169/c14 ,\u2_Display/n5576 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u14  (
    .a(\u2_Display/n5559 ),
    .b(1'b1),
    .c(\u2_Display/add169/c14 ),
    .o({\u2_Display/add169/c15 ,\u2_Display/n5576 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u15  (
    .a(\u2_Display/n5558 ),
    .b(1'b1),
    .c(\u2_Display/add169/c15 ),
    .o({\u2_Display/add169/c16 ,\u2_Display/n5576 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u16  (
    .a(\u2_Display/n5557 ),
    .b(1'b1),
    .c(\u2_Display/add169/c16 ),
    .o({\u2_Display/add169/c17 ,\u2_Display/n5576 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u17  (
    .a(\u2_Display/n5556 ),
    .b(1'b1),
    .c(\u2_Display/add169/c17 ),
    .o({\u2_Display/add169/c18 ,\u2_Display/n5576 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u18  (
    .a(\u2_Display/n5555 ),
    .b(1'b1),
    .c(\u2_Display/add169/c18 ),
    .o({\u2_Display/add169/c19 ,\u2_Display/n5576 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u19  (
    .a(\u2_Display/n5554 ),
    .b(1'b1),
    .c(\u2_Display/add169/c19 ),
    .o({\u2_Display/add169/c20 ,\u2_Display/n5576 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u2  (
    .a(\u2_Display/n5571 ),
    .b(1'b1),
    .c(\u2_Display/add169/c2 ),
    .o({\u2_Display/add169/c3 ,\u2_Display/n5576 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u20  (
    .a(\u2_Display/n5553 ),
    .b(1'b1),
    .c(\u2_Display/add169/c20 ),
    .o({\u2_Display/add169/c21 ,\u2_Display/n5576 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u21  (
    .a(\u2_Display/n5552 ),
    .b(1'b1),
    .c(\u2_Display/add169/c21 ),
    .o({\u2_Display/add169/c22 ,\u2_Display/n5576 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u22  (
    .a(\u2_Display/n5551 ),
    .b(1'b1),
    .c(\u2_Display/add169/c22 ),
    .o({\u2_Display/add169/c23 ,\u2_Display/n5576 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u23  (
    .a(\u2_Display/n5550 ),
    .b(1'b1),
    .c(\u2_Display/add169/c23 ),
    .o({\u2_Display/add169/c24 ,\u2_Display/n5576 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u24  (
    .a(\u2_Display/n5549 ),
    .b(1'b1),
    .c(\u2_Display/add169/c24 ),
    .o({\u2_Display/add169/c25 ,\u2_Display/n5576 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u25  (
    .a(\u2_Display/n5548 ),
    .b(1'b1),
    .c(\u2_Display/add169/c25 ),
    .o({\u2_Display/add169/c26 ,\u2_Display/n5576 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u26  (
    .a(\u2_Display/n5547 ),
    .b(1'b1),
    .c(\u2_Display/add169/c26 ),
    .o({\u2_Display/add169/c27 ,\u2_Display/n5576 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u27  (
    .a(\u2_Display/n5546 ),
    .b(1'b1),
    .c(\u2_Display/add169/c27 ),
    .o({\u2_Display/add169/c28 ,\u2_Display/n5576 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u28  (
    .a(\u2_Display/n5545 ),
    .b(1'b1),
    .c(\u2_Display/add169/c28 ),
    .o({\u2_Display/add169/c29 ,\u2_Display/n5576 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u29  (
    .a(\u2_Display/n5544 ),
    .b(1'b1),
    .c(\u2_Display/add169/c29 ),
    .o({\u2_Display/add169/c30 ,\u2_Display/n5576 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u3  (
    .a(\u2_Display/n5570 ),
    .b(1'b1),
    .c(\u2_Display/add169/c3 ),
    .o({\u2_Display/add169/c4 ,\u2_Display/n5576 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u30  (
    .a(\u2_Display/n5543 ),
    .b(1'b1),
    .c(\u2_Display/add169/c30 ),
    .o({\u2_Display/add169/c31 ,\u2_Display/n5576 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u31  (
    .a(\u2_Display/n5542 ),
    .b(1'b1),
    .c(\u2_Display/add169/c31 ),
    .o({open_n1075,\u2_Display/n5576 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u4  (
    .a(\u2_Display/n5569 ),
    .b(1'b1),
    .c(\u2_Display/add169/c4 ),
    .o({\u2_Display/add169/c5 ,\u2_Display/n5576 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u5  (
    .a(\u2_Display/n5568 ),
    .b(1'b1),
    .c(\u2_Display/add169/c5 ),
    .o({\u2_Display/add169/c6 ,\u2_Display/n5576 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u6  (
    .a(\u2_Display/n5567 ),
    .b(1'b1),
    .c(\u2_Display/add169/c6 ),
    .o({\u2_Display/add169/c7 ,\u2_Display/n5576 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u7  (
    .a(\u2_Display/n5566 ),
    .b(1'b1),
    .c(\u2_Display/add169/c7 ),
    .o({\u2_Display/add169/c8 ,\u2_Display/n5576 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u8  (
    .a(\u2_Display/n5565 ),
    .b(1'b1),
    .c(\u2_Display/add169/c8 ),
    .o({\u2_Display/add169/c9 ,\u2_Display/n5576 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add169/u9  (
    .a(\u2_Display/n5564 ),
    .b(1'b1),
    .c(\u2_Display/add169/c9 ),
    .o({\u2_Display/add169/c10 ,\u2_Display/n5576 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add169/ucin  (
    .a(1'b1),
    .o({\u2_Display/add169/c0 ,open_n1078}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u0  (
    .a(\u2_Display/n5608 ),
    .b(1'b1),
    .c(\u2_Display/add170/c0 ),
    .o({\u2_Display/add170/c1 ,\u2_Display/n5611 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u1  (
    .a(\u2_Display/n5607 ),
    .b(1'b1),
    .c(\u2_Display/add170/c1 ),
    .o({\u2_Display/add170/c2 ,\u2_Display/n5611 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u10  (
    .a(\u2_Display/n5598 ),
    .b(1'b1),
    .c(\u2_Display/add170/c10 ),
    .o({\u2_Display/add170/c11 ,\u2_Display/n5611 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u11  (
    .a(\u2_Display/n5597 ),
    .b(1'b0),
    .c(\u2_Display/add170/c11 ),
    .o({\u2_Display/add170/c12 ,\u2_Display/n5611 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u12  (
    .a(\u2_Display/n5596 ),
    .b(1'b1),
    .c(\u2_Display/add170/c12 ),
    .o({\u2_Display/add170/c13 ,\u2_Display/n5611 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u13  (
    .a(\u2_Display/n5595 ),
    .b(1'b1),
    .c(\u2_Display/add170/c13 ),
    .o({\u2_Display/add170/c14 ,\u2_Display/n5611 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u14  (
    .a(\u2_Display/n5594 ),
    .b(1'b1),
    .c(\u2_Display/add170/c14 ),
    .o({\u2_Display/add170/c15 ,\u2_Display/n5611 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u15  (
    .a(\u2_Display/n5593 ),
    .b(1'b1),
    .c(\u2_Display/add170/c15 ),
    .o({\u2_Display/add170/c16 ,\u2_Display/n5611 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u16  (
    .a(\u2_Display/n5592 ),
    .b(1'b1),
    .c(\u2_Display/add170/c16 ),
    .o({\u2_Display/add170/c17 ,\u2_Display/n5611 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u17  (
    .a(\u2_Display/n5591 ),
    .b(1'b1),
    .c(\u2_Display/add170/c17 ),
    .o({\u2_Display/add170/c18 ,\u2_Display/n5611 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u18  (
    .a(\u2_Display/n5590 ),
    .b(1'b1),
    .c(\u2_Display/add170/c18 ),
    .o({\u2_Display/add170/c19 ,\u2_Display/n5611 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u19  (
    .a(\u2_Display/n5589 ),
    .b(1'b1),
    .c(\u2_Display/add170/c19 ),
    .o({\u2_Display/add170/c20 ,\u2_Display/n5611 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u2  (
    .a(\u2_Display/n5606 ),
    .b(1'b1),
    .c(\u2_Display/add170/c2 ),
    .o({\u2_Display/add170/c3 ,\u2_Display/n5611 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u20  (
    .a(\u2_Display/n5588 ),
    .b(1'b1),
    .c(\u2_Display/add170/c20 ),
    .o({\u2_Display/add170/c21 ,\u2_Display/n5611 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u21  (
    .a(\u2_Display/n5587 ),
    .b(1'b1),
    .c(\u2_Display/add170/c21 ),
    .o({\u2_Display/add170/c22 ,\u2_Display/n5611 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u22  (
    .a(\u2_Display/n5586 ),
    .b(1'b1),
    .c(\u2_Display/add170/c22 ),
    .o({\u2_Display/add170/c23 ,\u2_Display/n5611 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u23  (
    .a(\u2_Display/n5585 ),
    .b(1'b1),
    .c(\u2_Display/add170/c23 ),
    .o({\u2_Display/add170/c24 ,\u2_Display/n5611 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u24  (
    .a(\u2_Display/n5584 ),
    .b(1'b1),
    .c(\u2_Display/add170/c24 ),
    .o({\u2_Display/add170/c25 ,\u2_Display/n5611 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u25  (
    .a(\u2_Display/n5583 ),
    .b(1'b1),
    .c(\u2_Display/add170/c25 ),
    .o({\u2_Display/add170/c26 ,\u2_Display/n5611 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u26  (
    .a(\u2_Display/n5582 ),
    .b(1'b1),
    .c(\u2_Display/add170/c26 ),
    .o({\u2_Display/add170/c27 ,\u2_Display/n5611 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u27  (
    .a(\u2_Display/n5581 ),
    .b(1'b1),
    .c(\u2_Display/add170/c27 ),
    .o({\u2_Display/add170/c28 ,\u2_Display/n5611 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u28  (
    .a(\u2_Display/n5580 ),
    .b(1'b1),
    .c(\u2_Display/add170/c28 ),
    .o({\u2_Display/add170/c29 ,\u2_Display/n5611 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u29  (
    .a(\u2_Display/n5579 ),
    .b(1'b1),
    .c(\u2_Display/add170/c29 ),
    .o({\u2_Display/add170/c30 ,\u2_Display/n5611 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u3  (
    .a(\u2_Display/n5605 ),
    .b(1'b1),
    .c(\u2_Display/add170/c3 ),
    .o({\u2_Display/add170/c4 ,\u2_Display/n5611 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u30  (
    .a(\u2_Display/n5578 ),
    .b(1'b1),
    .c(\u2_Display/add170/c30 ),
    .o({\u2_Display/add170/c31 ,\u2_Display/n5611 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u31  (
    .a(\u2_Display/n5577 ),
    .b(1'b1),
    .c(\u2_Display/add170/c31 ),
    .o({open_n1079,\u2_Display/n5611 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u4  (
    .a(\u2_Display/n5604 ),
    .b(1'b1),
    .c(\u2_Display/add170/c4 ),
    .o({\u2_Display/add170/c5 ,\u2_Display/n5611 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u5  (
    .a(\u2_Display/n5603 ),
    .b(1'b1),
    .c(\u2_Display/add170/c5 ),
    .o({\u2_Display/add170/c6 ,\u2_Display/n5611 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u6  (
    .a(\u2_Display/n5602 ),
    .b(1'b1),
    .c(\u2_Display/add170/c6 ),
    .o({\u2_Display/add170/c7 ,\u2_Display/n5611 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u7  (
    .a(\u2_Display/n5601 ),
    .b(1'b1),
    .c(\u2_Display/add170/c7 ),
    .o({\u2_Display/add170/c8 ,\u2_Display/n5611 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u8  (
    .a(\u2_Display/n5600 ),
    .b(1'b1),
    .c(\u2_Display/add170/c8 ),
    .o({\u2_Display/add170/c9 ,\u2_Display/n5611 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add170/u9  (
    .a(\u2_Display/n5599 ),
    .b(1'b0),
    .c(\u2_Display/add170/c9 ),
    .o({\u2_Display/add170/c10 ,\u2_Display/n5611 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add170/ucin  (
    .a(1'b1),
    .o({\u2_Display/add170/c0 ,open_n1082}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u0  (
    .a(\u2_Display/n5643 ),
    .b(1'b1),
    .c(\u2_Display/add171/c0 ),
    .o({\u2_Display/add171/c1 ,\u2_Display/n5646 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u1  (
    .a(\u2_Display/n5642 ),
    .b(1'b1),
    .c(\u2_Display/add171/c1 ),
    .o({\u2_Display/add171/c2 ,\u2_Display/n5646 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u10  (
    .a(\u2_Display/n5633 ),
    .b(1'b0),
    .c(\u2_Display/add171/c10 ),
    .o({\u2_Display/add171/c11 ,\u2_Display/n5646 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u11  (
    .a(\u2_Display/n5632 ),
    .b(1'b1),
    .c(\u2_Display/add171/c11 ),
    .o({\u2_Display/add171/c12 ,\u2_Display/n5646 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u12  (
    .a(\u2_Display/n5631 ),
    .b(1'b1),
    .c(\u2_Display/add171/c12 ),
    .o({\u2_Display/add171/c13 ,\u2_Display/n5646 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u13  (
    .a(\u2_Display/n5630 ),
    .b(1'b1),
    .c(\u2_Display/add171/c13 ),
    .o({\u2_Display/add171/c14 ,\u2_Display/n5646 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u14  (
    .a(\u2_Display/n5629 ),
    .b(1'b1),
    .c(\u2_Display/add171/c14 ),
    .o({\u2_Display/add171/c15 ,\u2_Display/n5646 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u15  (
    .a(\u2_Display/n5628 ),
    .b(1'b1),
    .c(\u2_Display/add171/c15 ),
    .o({\u2_Display/add171/c16 ,\u2_Display/n5646 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u16  (
    .a(\u2_Display/n5627 ),
    .b(1'b1),
    .c(\u2_Display/add171/c16 ),
    .o({\u2_Display/add171/c17 ,\u2_Display/n5646 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u17  (
    .a(\u2_Display/n5626 ),
    .b(1'b1),
    .c(\u2_Display/add171/c17 ),
    .o({\u2_Display/add171/c18 ,\u2_Display/n5646 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u18  (
    .a(\u2_Display/n5625 ),
    .b(1'b1),
    .c(\u2_Display/add171/c18 ),
    .o({\u2_Display/add171/c19 ,\u2_Display/n5646 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u19  (
    .a(\u2_Display/n5624 ),
    .b(1'b1),
    .c(\u2_Display/add171/c19 ),
    .o({\u2_Display/add171/c20 ,\u2_Display/n5646 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u2  (
    .a(\u2_Display/n5641 ),
    .b(1'b1),
    .c(\u2_Display/add171/c2 ),
    .o({\u2_Display/add171/c3 ,\u2_Display/n5646 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u20  (
    .a(\u2_Display/n5623 ),
    .b(1'b1),
    .c(\u2_Display/add171/c20 ),
    .o({\u2_Display/add171/c21 ,\u2_Display/n5646 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u21  (
    .a(\u2_Display/n5622 ),
    .b(1'b1),
    .c(\u2_Display/add171/c21 ),
    .o({\u2_Display/add171/c22 ,\u2_Display/n5646 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u22  (
    .a(\u2_Display/n5621 ),
    .b(1'b1),
    .c(\u2_Display/add171/c22 ),
    .o({\u2_Display/add171/c23 ,\u2_Display/n5646 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u23  (
    .a(\u2_Display/n5620 ),
    .b(1'b1),
    .c(\u2_Display/add171/c23 ),
    .o({\u2_Display/add171/c24 ,\u2_Display/n5646 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u24  (
    .a(\u2_Display/n5619 ),
    .b(1'b1),
    .c(\u2_Display/add171/c24 ),
    .o({\u2_Display/add171/c25 ,\u2_Display/n5646 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u25  (
    .a(\u2_Display/n5618 ),
    .b(1'b1),
    .c(\u2_Display/add171/c25 ),
    .o({\u2_Display/add171/c26 ,\u2_Display/n5646 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u26  (
    .a(\u2_Display/n5617 ),
    .b(1'b1),
    .c(\u2_Display/add171/c26 ),
    .o({\u2_Display/add171/c27 ,\u2_Display/n5646 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u27  (
    .a(\u2_Display/n5616 ),
    .b(1'b1),
    .c(\u2_Display/add171/c27 ),
    .o({\u2_Display/add171/c28 ,\u2_Display/n5646 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u28  (
    .a(\u2_Display/n5615 ),
    .b(1'b1),
    .c(\u2_Display/add171/c28 ),
    .o({\u2_Display/add171/c29 ,\u2_Display/n5646 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u29  (
    .a(\u2_Display/n5614 ),
    .b(1'b1),
    .c(\u2_Display/add171/c29 ),
    .o({\u2_Display/add171/c30 ,\u2_Display/n5646 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u3  (
    .a(\u2_Display/n5640 ),
    .b(1'b1),
    .c(\u2_Display/add171/c3 ),
    .o({\u2_Display/add171/c4 ,\u2_Display/n5646 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u30  (
    .a(\u2_Display/n5613 ),
    .b(1'b1),
    .c(\u2_Display/add171/c30 ),
    .o({\u2_Display/add171/c31 ,\u2_Display/n5646 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u31  (
    .a(\u2_Display/n5612 ),
    .b(1'b1),
    .c(\u2_Display/add171/c31 ),
    .o({open_n1083,\u2_Display/n5646 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u4  (
    .a(\u2_Display/n5639 ),
    .b(1'b1),
    .c(\u2_Display/add171/c4 ),
    .o({\u2_Display/add171/c5 ,\u2_Display/n5646 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u5  (
    .a(\u2_Display/n5638 ),
    .b(1'b1),
    .c(\u2_Display/add171/c5 ),
    .o({\u2_Display/add171/c6 ,\u2_Display/n5646 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u6  (
    .a(\u2_Display/n5637 ),
    .b(1'b1),
    .c(\u2_Display/add171/c6 ),
    .o({\u2_Display/add171/c7 ,\u2_Display/n5646 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u7  (
    .a(\u2_Display/n5636 ),
    .b(1'b1),
    .c(\u2_Display/add171/c7 ),
    .o({\u2_Display/add171/c8 ,\u2_Display/n5646 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u8  (
    .a(\u2_Display/n5635 ),
    .b(1'b0),
    .c(\u2_Display/add171/c8 ),
    .o({\u2_Display/add171/c9 ,\u2_Display/n5646 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add171/u9  (
    .a(\u2_Display/n5634 ),
    .b(1'b1),
    .c(\u2_Display/add171/c9 ),
    .o({\u2_Display/add171/c10 ,\u2_Display/n5646 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add171/ucin  (
    .a(1'b1),
    .o({\u2_Display/add171/c0 ,open_n1086}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add172/u0  (
    .a(\u2_Display/n5678 ),
    .b(1'b1),
    .c(\u2_Display/add172/c0 ),
    .o({\u2_Display/add172/c1 ,\u2_Display/n5681 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add172/u1  (
    .a(\u2_Display/n5677 ),
    .b(1'b1),
    .c(\u2_Display/add172/c1 ),
    .o({\u2_Display/add172/c2 ,\u2_Display/n5681 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add172/u2  (
    .a(\u2_Display/n5676 ),
    .b(1'b1),
    .c(\u2_Display/add172/c2 ),
    .o({\u2_Display/add172/c3 ,\u2_Display/n5681 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add172/u3  (
    .a(\u2_Display/n5675 ),
    .b(1'b1),
    .c(\u2_Display/add172/c3 ),
    .o({\u2_Display/add172/c4 ,\u2_Display/n5681 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add172/u4  (
    .a(\u2_Display/n5674 ),
    .b(1'b1),
    .c(\u2_Display/add172/c4 ),
    .o({\u2_Display/add172/c5 ,\u2_Display/n5681 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add172/u5  (
    .a(\u2_Display/n5673 ),
    .b(1'b1),
    .c(\u2_Display/add172/c5 ),
    .o({\u2_Display/add172/c6 ,\u2_Display/n5681 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add172/u6  (
    .a(\u2_Display/n5672 ),
    .b(1'b1),
    .c(\u2_Display/add172/c6 ),
    .o({\u2_Display/add172/c7 ,\u2_Display/n5681 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add172/u7  (
    .a(\u2_Display/n5671 ),
    .b(1'b0),
    .c(\u2_Display/add172/c7 ),
    .o({\u2_Display/add172/c8 ,\u2_Display/n5681 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add172/u8  (
    .a(\u2_Display/n5670 ),
    .b(1'b1),
    .c(\u2_Display/add172/c8 ),
    .o({\u2_Display/add172/c9 ,\u2_Display/n5681 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add172/u9  (
    .a(\u2_Display/n5669 ),
    .b(1'b0),
    .c(\u2_Display/add172/c9 ),
    .o({open_n1087,\u2_Display/n5681 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add172/ucin  (
    .a(1'b1),
    .o({\u2_Display/add172/c0 ,open_n1090}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u0  (
    .a(\u2_Display/counta [0]),
    .b(1'b1),
    .c(\u2_Display/add18/c0 ),
    .o({\u2_Display/add18/c1 ,\u2_Display/n419 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u1  (
    .a(\u2_Display/counta [1]),
    .b(1'b1),
    .c(\u2_Display/add18/c1 ),
    .o({\u2_Display/add18/c2 ,\u2_Display/n419 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u10  (
    .a(\u2_Display/counta [10]),
    .b(1'b1),
    .c(\u2_Display/add18/c10 ),
    .o({\u2_Display/add18/c11 ,\u2_Display/n419 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u11  (
    .a(\u2_Display/counta [11]),
    .b(1'b1),
    .c(\u2_Display/add18/c11 ),
    .o({\u2_Display/add18/c12 ,\u2_Display/n419 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u12  (
    .a(\u2_Display/counta [12]),
    .b(1'b1),
    .c(\u2_Display/add18/c12 ),
    .o({\u2_Display/add18/c13 ,\u2_Display/n419 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u13  (
    .a(\u2_Display/counta [13]),
    .b(1'b1),
    .c(\u2_Display/add18/c13 ),
    .o({\u2_Display/add18/c14 ,\u2_Display/n419 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u14  (
    .a(\u2_Display/counta [14]),
    .b(1'b1),
    .c(\u2_Display/add18/c14 ),
    .o({\u2_Display/add18/c15 ,\u2_Display/n419 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u15  (
    .a(\u2_Display/counta [15]),
    .b(1'b1),
    .c(\u2_Display/add18/c15 ),
    .o({\u2_Display/add18/c16 ,\u2_Display/n419 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u16  (
    .a(\u2_Display/counta [16]),
    .b(1'b1),
    .c(\u2_Display/add18/c16 ),
    .o({\u2_Display/add18/c17 ,\u2_Display/n419 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u17  (
    .a(\u2_Display/counta [17]),
    .b(1'b1),
    .c(\u2_Display/add18/c17 ),
    .o({\u2_Display/add18/c18 ,\u2_Display/n419 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u18  (
    .a(\u2_Display/counta [18]),
    .b(1'b1),
    .c(\u2_Display/add18/c18 ),
    .o({\u2_Display/add18/c19 ,\u2_Display/n419 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u19  (
    .a(\u2_Display/counta [19]),
    .b(1'b1),
    .c(\u2_Display/add18/c19 ),
    .o({\u2_Display/add18/c20 ,\u2_Display/n419 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u2  (
    .a(\u2_Display/counta [2]),
    .b(1'b1),
    .c(\u2_Display/add18/c2 ),
    .o({\u2_Display/add18/c3 ,\u2_Display/n419 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u20  (
    .a(\u2_Display/counta [20]),
    .b(1'b1),
    .c(\u2_Display/add18/c20 ),
    .o({\u2_Display/add18/c21 ,\u2_Display/n419 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u21  (
    .a(\u2_Display/counta [21]),
    .b(1'b1),
    .c(\u2_Display/add18/c21 ),
    .o({\u2_Display/add18/c22 ,\u2_Display/n419 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u22  (
    .a(\u2_Display/counta [22]),
    .b(1'b1),
    .c(\u2_Display/add18/c22 ),
    .o({\u2_Display/add18/c23 ,\u2_Display/n419 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u23  (
    .a(\u2_Display/counta [23]),
    .b(1'b1),
    .c(\u2_Display/add18/c23 ),
    .o({\u2_Display/add18/c24 ,\u2_Display/n419 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u24  (
    .a(\u2_Display/counta [24]),
    .b(1'b1),
    .c(\u2_Display/add18/c24 ),
    .o({\u2_Display/add18/c25 ,\u2_Display/n419 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u25  (
    .a(\u2_Display/counta [25]),
    .b(1'b0),
    .c(\u2_Display/add18/c25 ),
    .o({\u2_Display/add18/c26 ,\u2_Display/n419 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u26  (
    .a(\u2_Display/counta [26]),
    .b(1'b1),
    .c(\u2_Display/add18/c26 ),
    .o({\u2_Display/add18/c27 ,\u2_Display/n419 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u27  (
    .a(\u2_Display/counta [27]),
    .b(1'b0),
    .c(\u2_Display/add18/c27 ),
    .o({\u2_Display/add18/c28 ,\u2_Display/n419 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u28  (
    .a(\u2_Display/counta [28]),
    .b(1'b0),
    .c(\u2_Display/add18/c28 ),
    .o({\u2_Display/add18/c29 ,\u2_Display/n419 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u29  (
    .a(\u2_Display/counta [29]),
    .b(1'b0),
    .c(\u2_Display/add18/c29 ),
    .o({\u2_Display/add18/c30 ,\u2_Display/n419 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u3  (
    .a(\u2_Display/counta [3]),
    .b(1'b1),
    .c(\u2_Display/add18/c3 ),
    .o({\u2_Display/add18/c4 ,\u2_Display/n419 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u30  (
    .a(\u2_Display/counta [30]),
    .b(1'b0),
    .c(\u2_Display/add18/c30 ),
    .o({\u2_Display/add18/c31 ,\u2_Display/n419 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u31  (
    .a(\u2_Display/counta [31]),
    .b(1'b0),
    .c(\u2_Display/add18/c31 ),
    .o({open_n1091,\u2_Display/n419 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u4  (
    .a(\u2_Display/counta [4]),
    .b(1'b1),
    .c(\u2_Display/add18/c4 ),
    .o({\u2_Display/add18/c5 ,\u2_Display/n419 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u5  (
    .a(\u2_Display/counta [5]),
    .b(1'b1),
    .c(\u2_Display/add18/c5 ),
    .o({\u2_Display/add18/c6 ,\u2_Display/n419 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u6  (
    .a(\u2_Display/counta [6]),
    .b(1'b1),
    .c(\u2_Display/add18/c6 ),
    .o({\u2_Display/add18/c7 ,\u2_Display/n419 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u7  (
    .a(\u2_Display/counta [7]),
    .b(1'b1),
    .c(\u2_Display/add18/c7 ),
    .o({\u2_Display/add18/c8 ,\u2_Display/n419 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u8  (
    .a(\u2_Display/counta [8]),
    .b(1'b1),
    .c(\u2_Display/add18/c8 ),
    .o({\u2_Display/add18/c9 ,\u2_Display/n419 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add18/u9  (
    .a(\u2_Display/counta [9]),
    .b(1'b1),
    .c(\u2_Display/add18/c9 ),
    .o({\u2_Display/add18/c10 ,\u2_Display/n419 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add18/ucin  (
    .a(1'b1),
    .o({\u2_Display/add18/c0 ,open_n1094}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u0  (
    .a(\u2_Display/n451 ),
    .b(1'b1),
    .c(\u2_Display/add19/c0 ),
    .o({\u2_Display/add19/c1 ,\u2_Display/n454 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u1  (
    .a(\u2_Display/n450 ),
    .b(1'b1),
    .c(\u2_Display/add19/c1 ),
    .o({\u2_Display/add19/c2 ,\u2_Display/n454 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u10  (
    .a(\u2_Display/n441 ),
    .b(1'b1),
    .c(\u2_Display/add19/c10 ),
    .o({\u2_Display/add19/c11 ,\u2_Display/n454 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u11  (
    .a(\u2_Display/n440 ),
    .b(1'b1),
    .c(\u2_Display/add19/c11 ),
    .o({\u2_Display/add19/c12 ,\u2_Display/n454 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u12  (
    .a(\u2_Display/n439 ),
    .b(1'b1),
    .c(\u2_Display/add19/c12 ),
    .o({\u2_Display/add19/c13 ,\u2_Display/n454 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u13  (
    .a(\u2_Display/n438 ),
    .b(1'b1),
    .c(\u2_Display/add19/c13 ),
    .o({\u2_Display/add19/c14 ,\u2_Display/n454 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u14  (
    .a(\u2_Display/n437 ),
    .b(1'b1),
    .c(\u2_Display/add19/c14 ),
    .o({\u2_Display/add19/c15 ,\u2_Display/n454 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u15  (
    .a(\u2_Display/n436 ),
    .b(1'b1),
    .c(\u2_Display/add19/c15 ),
    .o({\u2_Display/add19/c16 ,\u2_Display/n454 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u16  (
    .a(\u2_Display/n435 ),
    .b(1'b1),
    .c(\u2_Display/add19/c16 ),
    .o({\u2_Display/add19/c17 ,\u2_Display/n454 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u17  (
    .a(\u2_Display/n434 ),
    .b(1'b1),
    .c(\u2_Display/add19/c17 ),
    .o({\u2_Display/add19/c18 ,\u2_Display/n454 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u18  (
    .a(\u2_Display/n433 ),
    .b(1'b1),
    .c(\u2_Display/add19/c18 ),
    .o({\u2_Display/add19/c19 ,\u2_Display/n454 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u19  (
    .a(\u2_Display/n432 ),
    .b(1'b1),
    .c(\u2_Display/add19/c19 ),
    .o({\u2_Display/add19/c20 ,\u2_Display/n454 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u2  (
    .a(\u2_Display/n449 ),
    .b(1'b1),
    .c(\u2_Display/add19/c2 ),
    .o({\u2_Display/add19/c3 ,\u2_Display/n454 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u20  (
    .a(\u2_Display/n431 ),
    .b(1'b1),
    .c(\u2_Display/add19/c20 ),
    .o({\u2_Display/add19/c21 ,\u2_Display/n454 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u21  (
    .a(\u2_Display/n430 ),
    .b(1'b1),
    .c(\u2_Display/add19/c21 ),
    .o({\u2_Display/add19/c22 ,\u2_Display/n454 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u22  (
    .a(\u2_Display/n429 ),
    .b(1'b1),
    .c(\u2_Display/add19/c22 ),
    .o({\u2_Display/add19/c23 ,\u2_Display/n454 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u23  (
    .a(\u2_Display/n428 ),
    .b(1'b1),
    .c(\u2_Display/add19/c23 ),
    .o({\u2_Display/add19/c24 ,\u2_Display/n454 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u24  (
    .a(\u2_Display/n427 ),
    .b(1'b0),
    .c(\u2_Display/add19/c24 ),
    .o({\u2_Display/add19/c25 ,\u2_Display/n454 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u25  (
    .a(\u2_Display/n426 ),
    .b(1'b1),
    .c(\u2_Display/add19/c25 ),
    .o({\u2_Display/add19/c26 ,\u2_Display/n454 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u26  (
    .a(\u2_Display/n425 ),
    .b(1'b0),
    .c(\u2_Display/add19/c26 ),
    .o({\u2_Display/add19/c27 ,\u2_Display/n454 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u27  (
    .a(\u2_Display/n424 ),
    .b(1'b0),
    .c(\u2_Display/add19/c27 ),
    .o({\u2_Display/add19/c28 ,\u2_Display/n454 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u28  (
    .a(\u2_Display/n423 ),
    .b(1'b0),
    .c(\u2_Display/add19/c28 ),
    .o({\u2_Display/add19/c29 ,\u2_Display/n454 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u29  (
    .a(\u2_Display/n422 ),
    .b(1'b0),
    .c(\u2_Display/add19/c29 ),
    .o({\u2_Display/add19/c30 ,\u2_Display/n454 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u3  (
    .a(\u2_Display/n448 ),
    .b(1'b1),
    .c(\u2_Display/add19/c3 ),
    .o({\u2_Display/add19/c4 ,\u2_Display/n454 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u30  (
    .a(\u2_Display/n421 ),
    .b(1'b0),
    .c(\u2_Display/add19/c30 ),
    .o({\u2_Display/add19/c31 ,\u2_Display/n454 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u31  (
    .a(\u2_Display/n420 ),
    .b(1'b1),
    .c(\u2_Display/add19/c31 ),
    .o({open_n1095,\u2_Display/n454 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u4  (
    .a(\u2_Display/n447 ),
    .b(1'b1),
    .c(\u2_Display/add19/c4 ),
    .o({\u2_Display/add19/c5 ,\u2_Display/n454 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u5  (
    .a(\u2_Display/n446 ),
    .b(1'b1),
    .c(\u2_Display/add19/c5 ),
    .o({\u2_Display/add19/c6 ,\u2_Display/n454 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u6  (
    .a(\u2_Display/n445 ),
    .b(1'b1),
    .c(\u2_Display/add19/c6 ),
    .o({\u2_Display/add19/c7 ,\u2_Display/n454 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u7  (
    .a(\u2_Display/n444 ),
    .b(1'b1),
    .c(\u2_Display/add19/c7 ),
    .o({\u2_Display/add19/c8 ,\u2_Display/n454 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u8  (
    .a(\u2_Display/n443 ),
    .b(1'b1),
    .c(\u2_Display/add19/c8 ),
    .o({\u2_Display/add19/c9 ,\u2_Display/n454 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add19/u9  (
    .a(\u2_Display/n442 ),
    .b(1'b1),
    .c(\u2_Display/add19/c9 ),
    .o({\u2_Display/add19/c10 ,\u2_Display/n454 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add19/ucin  (
    .a(1'b1),
    .o({\u2_Display/add19/c0 ,open_n1098}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u0  (
    .a(\u2_Display/n486 ),
    .b(1'b1),
    .c(\u2_Display/add20/c0 ),
    .o({\u2_Display/add20/c1 ,\u2_Display/n489 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u1  (
    .a(\u2_Display/n485 ),
    .b(1'b1),
    .c(\u2_Display/add20/c1 ),
    .o({\u2_Display/add20/c2 ,\u2_Display/n489 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u10  (
    .a(\u2_Display/n476 ),
    .b(1'b1),
    .c(\u2_Display/add20/c10 ),
    .o({\u2_Display/add20/c11 ,\u2_Display/n489 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u11  (
    .a(\u2_Display/n475 ),
    .b(1'b1),
    .c(\u2_Display/add20/c11 ),
    .o({\u2_Display/add20/c12 ,\u2_Display/n489 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u12  (
    .a(\u2_Display/n474 ),
    .b(1'b1),
    .c(\u2_Display/add20/c12 ),
    .o({\u2_Display/add20/c13 ,\u2_Display/n489 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u13  (
    .a(\u2_Display/n473 ),
    .b(1'b1),
    .c(\u2_Display/add20/c13 ),
    .o({\u2_Display/add20/c14 ,\u2_Display/n489 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u14  (
    .a(\u2_Display/n472 ),
    .b(1'b1),
    .c(\u2_Display/add20/c14 ),
    .o({\u2_Display/add20/c15 ,\u2_Display/n489 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u15  (
    .a(\u2_Display/n471 ),
    .b(1'b1),
    .c(\u2_Display/add20/c15 ),
    .o({\u2_Display/add20/c16 ,\u2_Display/n489 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u16  (
    .a(\u2_Display/n470 ),
    .b(1'b1),
    .c(\u2_Display/add20/c16 ),
    .o({\u2_Display/add20/c17 ,\u2_Display/n489 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u17  (
    .a(\u2_Display/n469 ),
    .b(1'b1),
    .c(\u2_Display/add20/c17 ),
    .o({\u2_Display/add20/c18 ,\u2_Display/n489 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u18  (
    .a(\u2_Display/n468 ),
    .b(1'b1),
    .c(\u2_Display/add20/c18 ),
    .o({\u2_Display/add20/c19 ,\u2_Display/n489 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u19  (
    .a(\u2_Display/n467 ),
    .b(1'b1),
    .c(\u2_Display/add20/c19 ),
    .o({\u2_Display/add20/c20 ,\u2_Display/n489 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u2  (
    .a(\u2_Display/n484 ),
    .b(1'b1),
    .c(\u2_Display/add20/c2 ),
    .o({\u2_Display/add20/c3 ,\u2_Display/n489 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u20  (
    .a(\u2_Display/n466 ),
    .b(1'b1),
    .c(\u2_Display/add20/c20 ),
    .o({\u2_Display/add20/c21 ,\u2_Display/n489 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u21  (
    .a(\u2_Display/n465 ),
    .b(1'b1),
    .c(\u2_Display/add20/c21 ),
    .o({\u2_Display/add20/c22 ,\u2_Display/n489 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u22  (
    .a(\u2_Display/n464 ),
    .b(1'b1),
    .c(\u2_Display/add20/c22 ),
    .o({\u2_Display/add20/c23 ,\u2_Display/n489 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u23  (
    .a(\u2_Display/n463 ),
    .b(1'b0),
    .c(\u2_Display/add20/c23 ),
    .o({\u2_Display/add20/c24 ,\u2_Display/n489 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u24  (
    .a(\u2_Display/n462 ),
    .b(1'b1),
    .c(\u2_Display/add20/c24 ),
    .o({\u2_Display/add20/c25 ,\u2_Display/n489 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u25  (
    .a(\u2_Display/n461 ),
    .b(1'b0),
    .c(\u2_Display/add20/c25 ),
    .o({\u2_Display/add20/c26 ,\u2_Display/n489 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u26  (
    .a(\u2_Display/n460 ),
    .b(1'b0),
    .c(\u2_Display/add20/c26 ),
    .o({\u2_Display/add20/c27 ,\u2_Display/n489 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u27  (
    .a(\u2_Display/n459 ),
    .b(1'b0),
    .c(\u2_Display/add20/c27 ),
    .o({\u2_Display/add20/c28 ,\u2_Display/n489 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u28  (
    .a(\u2_Display/n458 ),
    .b(1'b0),
    .c(\u2_Display/add20/c28 ),
    .o({\u2_Display/add20/c29 ,\u2_Display/n489 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u29  (
    .a(\u2_Display/n457 ),
    .b(1'b0),
    .c(\u2_Display/add20/c29 ),
    .o({\u2_Display/add20/c30 ,\u2_Display/n489 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u3  (
    .a(\u2_Display/n483 ),
    .b(1'b1),
    .c(\u2_Display/add20/c3 ),
    .o({\u2_Display/add20/c4 ,\u2_Display/n489 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u30  (
    .a(\u2_Display/n456 ),
    .b(1'b1),
    .c(\u2_Display/add20/c30 ),
    .o({\u2_Display/add20/c31 ,\u2_Display/n489 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u31  (
    .a(\u2_Display/n455 ),
    .b(1'b1),
    .c(\u2_Display/add20/c31 ),
    .o({open_n1099,\u2_Display/n489 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u4  (
    .a(\u2_Display/n482 ),
    .b(1'b1),
    .c(\u2_Display/add20/c4 ),
    .o({\u2_Display/add20/c5 ,\u2_Display/n489 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u5  (
    .a(\u2_Display/n481 ),
    .b(1'b1),
    .c(\u2_Display/add20/c5 ),
    .o({\u2_Display/add20/c6 ,\u2_Display/n489 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u6  (
    .a(\u2_Display/n480 ),
    .b(1'b1),
    .c(\u2_Display/add20/c6 ),
    .o({\u2_Display/add20/c7 ,\u2_Display/n489 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u7  (
    .a(\u2_Display/n479 ),
    .b(1'b1),
    .c(\u2_Display/add20/c7 ),
    .o({\u2_Display/add20/c8 ,\u2_Display/n489 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u8  (
    .a(\u2_Display/n478 ),
    .b(1'b1),
    .c(\u2_Display/add20/c8 ),
    .o({\u2_Display/add20/c9 ,\u2_Display/n489 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add20/u9  (
    .a(\u2_Display/n477 ),
    .b(1'b1),
    .c(\u2_Display/add20/c9 ),
    .o({\u2_Display/add20/c10 ,\u2_Display/n489 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add20/ucin  (
    .a(1'b1),
    .o({\u2_Display/add20/c0 ,open_n1102}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u0  (
    .a(\u2_Display/n521 ),
    .b(1'b1),
    .c(\u2_Display/add21/c0 ),
    .o({\u2_Display/add21/c1 ,\u2_Display/n524 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u1  (
    .a(\u2_Display/n520 ),
    .b(1'b1),
    .c(\u2_Display/add21/c1 ),
    .o({\u2_Display/add21/c2 ,\u2_Display/n524 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u10  (
    .a(\u2_Display/n511 ),
    .b(1'b1),
    .c(\u2_Display/add21/c10 ),
    .o({\u2_Display/add21/c11 ,\u2_Display/n524 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u11  (
    .a(\u2_Display/n510 ),
    .b(1'b1),
    .c(\u2_Display/add21/c11 ),
    .o({\u2_Display/add21/c12 ,\u2_Display/n524 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u12  (
    .a(\u2_Display/n509 ),
    .b(1'b1),
    .c(\u2_Display/add21/c12 ),
    .o({\u2_Display/add21/c13 ,\u2_Display/n524 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u13  (
    .a(\u2_Display/n508 ),
    .b(1'b1),
    .c(\u2_Display/add21/c13 ),
    .o({\u2_Display/add21/c14 ,\u2_Display/n524 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u14  (
    .a(\u2_Display/n507 ),
    .b(1'b1),
    .c(\u2_Display/add21/c14 ),
    .o({\u2_Display/add21/c15 ,\u2_Display/n524 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u15  (
    .a(\u2_Display/n506 ),
    .b(1'b1),
    .c(\u2_Display/add21/c15 ),
    .o({\u2_Display/add21/c16 ,\u2_Display/n524 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u16  (
    .a(\u2_Display/n505 ),
    .b(1'b1),
    .c(\u2_Display/add21/c16 ),
    .o({\u2_Display/add21/c17 ,\u2_Display/n524 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u17  (
    .a(\u2_Display/n504 ),
    .b(1'b1),
    .c(\u2_Display/add21/c17 ),
    .o({\u2_Display/add21/c18 ,\u2_Display/n524 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u18  (
    .a(\u2_Display/n503 ),
    .b(1'b1),
    .c(\u2_Display/add21/c18 ),
    .o({\u2_Display/add21/c19 ,\u2_Display/n524 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u19  (
    .a(\u2_Display/n502 ),
    .b(1'b1),
    .c(\u2_Display/add21/c19 ),
    .o({\u2_Display/add21/c20 ,\u2_Display/n524 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u2  (
    .a(\u2_Display/n519 ),
    .b(1'b1),
    .c(\u2_Display/add21/c2 ),
    .o({\u2_Display/add21/c3 ,\u2_Display/n524 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u20  (
    .a(\u2_Display/n501 ),
    .b(1'b1),
    .c(\u2_Display/add21/c20 ),
    .o({\u2_Display/add21/c21 ,\u2_Display/n524 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u21  (
    .a(\u2_Display/n500 ),
    .b(1'b1),
    .c(\u2_Display/add21/c21 ),
    .o({\u2_Display/add21/c22 ,\u2_Display/n524 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u22  (
    .a(\u2_Display/n499 ),
    .b(1'b0),
    .c(\u2_Display/add21/c22 ),
    .o({\u2_Display/add21/c23 ,\u2_Display/n524 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u23  (
    .a(\u2_Display/n498 ),
    .b(1'b1),
    .c(\u2_Display/add21/c23 ),
    .o({\u2_Display/add21/c24 ,\u2_Display/n524 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u24  (
    .a(\u2_Display/n497 ),
    .b(1'b0),
    .c(\u2_Display/add21/c24 ),
    .o({\u2_Display/add21/c25 ,\u2_Display/n524 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u25  (
    .a(\u2_Display/n496 ),
    .b(1'b0),
    .c(\u2_Display/add21/c25 ),
    .o({\u2_Display/add21/c26 ,\u2_Display/n524 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u26  (
    .a(\u2_Display/n495 ),
    .b(1'b0),
    .c(\u2_Display/add21/c26 ),
    .o({\u2_Display/add21/c27 ,\u2_Display/n524 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u27  (
    .a(\u2_Display/n494 ),
    .b(1'b0),
    .c(\u2_Display/add21/c27 ),
    .o({\u2_Display/add21/c28 ,\u2_Display/n524 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u28  (
    .a(\u2_Display/n493 ),
    .b(1'b0),
    .c(\u2_Display/add21/c28 ),
    .o({\u2_Display/add21/c29 ,\u2_Display/n524 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u29  (
    .a(\u2_Display/n492 ),
    .b(1'b1),
    .c(\u2_Display/add21/c29 ),
    .o({\u2_Display/add21/c30 ,\u2_Display/n524 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u3  (
    .a(\u2_Display/n518 ),
    .b(1'b1),
    .c(\u2_Display/add21/c3 ),
    .o({\u2_Display/add21/c4 ,\u2_Display/n524 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u30  (
    .a(\u2_Display/n491 ),
    .b(1'b1),
    .c(\u2_Display/add21/c30 ),
    .o({\u2_Display/add21/c31 ,\u2_Display/n524 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u31  (
    .a(\u2_Display/n490 ),
    .b(1'b1),
    .c(\u2_Display/add21/c31 ),
    .o({open_n1103,\u2_Display/n524 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u4  (
    .a(\u2_Display/n517 ),
    .b(1'b1),
    .c(\u2_Display/add21/c4 ),
    .o({\u2_Display/add21/c5 ,\u2_Display/n524 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u5  (
    .a(\u2_Display/n516 ),
    .b(1'b1),
    .c(\u2_Display/add21/c5 ),
    .o({\u2_Display/add21/c6 ,\u2_Display/n524 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u6  (
    .a(\u2_Display/n515 ),
    .b(1'b1),
    .c(\u2_Display/add21/c6 ),
    .o({\u2_Display/add21/c7 ,\u2_Display/n524 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u7  (
    .a(\u2_Display/n514 ),
    .b(1'b1),
    .c(\u2_Display/add21/c7 ),
    .o({\u2_Display/add21/c8 ,\u2_Display/n524 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u8  (
    .a(\u2_Display/n513 ),
    .b(1'b1),
    .c(\u2_Display/add21/c8 ),
    .o({\u2_Display/add21/c9 ,\u2_Display/n524 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add21/u9  (
    .a(\u2_Display/n512 ),
    .b(1'b1),
    .c(\u2_Display/add21/c9 ),
    .o({\u2_Display/add21/c10 ,\u2_Display/n524 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add21/ucin  (
    .a(1'b1),
    .o({\u2_Display/add21/c0 ,open_n1106}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u0  (
    .a(\u2_Display/n556 ),
    .b(1'b1),
    .c(\u2_Display/add22/c0 ),
    .o({\u2_Display/add22/c1 ,\u2_Display/n559 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u1  (
    .a(\u2_Display/n555 ),
    .b(1'b1),
    .c(\u2_Display/add22/c1 ),
    .o({\u2_Display/add22/c2 ,\u2_Display/n559 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u10  (
    .a(\u2_Display/n546 ),
    .b(1'b1),
    .c(\u2_Display/add22/c10 ),
    .o({\u2_Display/add22/c11 ,\u2_Display/n559 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u11  (
    .a(\u2_Display/n545 ),
    .b(1'b1),
    .c(\u2_Display/add22/c11 ),
    .o({\u2_Display/add22/c12 ,\u2_Display/n559 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u12  (
    .a(\u2_Display/n544 ),
    .b(1'b1),
    .c(\u2_Display/add22/c12 ),
    .o({\u2_Display/add22/c13 ,\u2_Display/n559 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u13  (
    .a(\u2_Display/n543 ),
    .b(1'b1),
    .c(\u2_Display/add22/c13 ),
    .o({\u2_Display/add22/c14 ,\u2_Display/n559 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u14  (
    .a(\u2_Display/n542 ),
    .b(1'b1),
    .c(\u2_Display/add22/c14 ),
    .o({\u2_Display/add22/c15 ,\u2_Display/n559 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u15  (
    .a(\u2_Display/n541 ),
    .b(1'b1),
    .c(\u2_Display/add22/c15 ),
    .o({\u2_Display/add22/c16 ,\u2_Display/n559 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u16  (
    .a(\u2_Display/n540 ),
    .b(1'b1),
    .c(\u2_Display/add22/c16 ),
    .o({\u2_Display/add22/c17 ,\u2_Display/n559 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u17  (
    .a(\u2_Display/n539 ),
    .b(1'b1),
    .c(\u2_Display/add22/c17 ),
    .o({\u2_Display/add22/c18 ,\u2_Display/n559 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u18  (
    .a(\u2_Display/n538 ),
    .b(1'b1),
    .c(\u2_Display/add22/c18 ),
    .o({\u2_Display/add22/c19 ,\u2_Display/n559 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u19  (
    .a(\u2_Display/n537 ),
    .b(1'b1),
    .c(\u2_Display/add22/c19 ),
    .o({\u2_Display/add22/c20 ,\u2_Display/n559 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u2  (
    .a(\u2_Display/n554 ),
    .b(1'b1),
    .c(\u2_Display/add22/c2 ),
    .o({\u2_Display/add22/c3 ,\u2_Display/n559 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u20  (
    .a(\u2_Display/n536 ),
    .b(1'b1),
    .c(\u2_Display/add22/c20 ),
    .o({\u2_Display/add22/c21 ,\u2_Display/n559 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u21  (
    .a(\u2_Display/n535 ),
    .b(1'b0),
    .c(\u2_Display/add22/c21 ),
    .o({\u2_Display/add22/c22 ,\u2_Display/n559 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u22  (
    .a(\u2_Display/n534 ),
    .b(1'b1),
    .c(\u2_Display/add22/c22 ),
    .o({\u2_Display/add22/c23 ,\u2_Display/n559 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u23  (
    .a(\u2_Display/n533 ),
    .b(1'b0),
    .c(\u2_Display/add22/c23 ),
    .o({\u2_Display/add22/c24 ,\u2_Display/n559 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u24  (
    .a(\u2_Display/n532 ),
    .b(1'b0),
    .c(\u2_Display/add22/c24 ),
    .o({\u2_Display/add22/c25 ,\u2_Display/n559 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u25  (
    .a(\u2_Display/n531 ),
    .b(1'b0),
    .c(\u2_Display/add22/c25 ),
    .o({\u2_Display/add22/c26 ,\u2_Display/n559 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u26  (
    .a(\u2_Display/n530 ),
    .b(1'b0),
    .c(\u2_Display/add22/c26 ),
    .o({\u2_Display/add22/c27 ,\u2_Display/n559 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u27  (
    .a(\u2_Display/n529 ),
    .b(1'b0),
    .c(\u2_Display/add22/c27 ),
    .o({\u2_Display/add22/c28 ,\u2_Display/n559 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u28  (
    .a(\u2_Display/n528 ),
    .b(1'b1),
    .c(\u2_Display/add22/c28 ),
    .o({\u2_Display/add22/c29 ,\u2_Display/n559 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u29  (
    .a(\u2_Display/n527 ),
    .b(1'b1),
    .c(\u2_Display/add22/c29 ),
    .o({\u2_Display/add22/c30 ,\u2_Display/n559 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u3  (
    .a(\u2_Display/n553 ),
    .b(1'b1),
    .c(\u2_Display/add22/c3 ),
    .o({\u2_Display/add22/c4 ,\u2_Display/n559 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u30  (
    .a(\u2_Display/n526 ),
    .b(1'b1),
    .c(\u2_Display/add22/c30 ),
    .o({\u2_Display/add22/c31 ,\u2_Display/n559 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u31  (
    .a(\u2_Display/n525 ),
    .b(1'b1),
    .c(\u2_Display/add22/c31 ),
    .o({open_n1107,\u2_Display/n559 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u4  (
    .a(\u2_Display/n552 ),
    .b(1'b1),
    .c(\u2_Display/add22/c4 ),
    .o({\u2_Display/add22/c5 ,\u2_Display/n559 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u5  (
    .a(\u2_Display/n551 ),
    .b(1'b1),
    .c(\u2_Display/add22/c5 ),
    .o({\u2_Display/add22/c6 ,\u2_Display/n559 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u6  (
    .a(\u2_Display/n550 ),
    .b(1'b1),
    .c(\u2_Display/add22/c6 ),
    .o({\u2_Display/add22/c7 ,\u2_Display/n559 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u7  (
    .a(\u2_Display/n549 ),
    .b(1'b1),
    .c(\u2_Display/add22/c7 ),
    .o({\u2_Display/add22/c8 ,\u2_Display/n559 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u8  (
    .a(\u2_Display/n548 ),
    .b(1'b1),
    .c(\u2_Display/add22/c8 ),
    .o({\u2_Display/add22/c9 ,\u2_Display/n559 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add22/u9  (
    .a(\u2_Display/n547 ),
    .b(1'b1),
    .c(\u2_Display/add22/c9 ),
    .o({\u2_Display/add22/c10 ,\u2_Display/n559 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add22/ucin  (
    .a(1'b1),
    .o({\u2_Display/add22/c0 ,open_n1110}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u0  (
    .a(\u2_Display/n591 ),
    .b(1'b1),
    .c(\u2_Display/add23/c0 ),
    .o({\u2_Display/add23/c1 ,\u2_Display/n594 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u1  (
    .a(\u2_Display/n590 ),
    .b(1'b1),
    .c(\u2_Display/add23/c1 ),
    .o({\u2_Display/add23/c2 ,\u2_Display/n594 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u10  (
    .a(\u2_Display/n581 ),
    .b(1'b1),
    .c(\u2_Display/add23/c10 ),
    .o({\u2_Display/add23/c11 ,\u2_Display/n594 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u11  (
    .a(\u2_Display/n580 ),
    .b(1'b1),
    .c(\u2_Display/add23/c11 ),
    .o({\u2_Display/add23/c12 ,\u2_Display/n594 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u12  (
    .a(\u2_Display/n579 ),
    .b(1'b1),
    .c(\u2_Display/add23/c12 ),
    .o({\u2_Display/add23/c13 ,\u2_Display/n594 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u13  (
    .a(\u2_Display/n578 ),
    .b(1'b1),
    .c(\u2_Display/add23/c13 ),
    .o({\u2_Display/add23/c14 ,\u2_Display/n594 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u14  (
    .a(\u2_Display/n577 ),
    .b(1'b1),
    .c(\u2_Display/add23/c14 ),
    .o({\u2_Display/add23/c15 ,\u2_Display/n594 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u15  (
    .a(\u2_Display/n576 ),
    .b(1'b1),
    .c(\u2_Display/add23/c15 ),
    .o({\u2_Display/add23/c16 ,\u2_Display/n594 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u16  (
    .a(\u2_Display/n575 ),
    .b(1'b1),
    .c(\u2_Display/add23/c16 ),
    .o({\u2_Display/add23/c17 ,\u2_Display/n594 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u17  (
    .a(\u2_Display/n574 ),
    .b(1'b1),
    .c(\u2_Display/add23/c17 ),
    .o({\u2_Display/add23/c18 ,\u2_Display/n594 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u18  (
    .a(\u2_Display/n573 ),
    .b(1'b1),
    .c(\u2_Display/add23/c18 ),
    .o({\u2_Display/add23/c19 ,\u2_Display/n594 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u19  (
    .a(\u2_Display/n572 ),
    .b(1'b1),
    .c(\u2_Display/add23/c19 ),
    .o({\u2_Display/add23/c20 ,\u2_Display/n594 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u2  (
    .a(\u2_Display/n589 ),
    .b(1'b1),
    .c(\u2_Display/add23/c2 ),
    .o({\u2_Display/add23/c3 ,\u2_Display/n594 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u20  (
    .a(\u2_Display/n571 ),
    .b(1'b0),
    .c(\u2_Display/add23/c20 ),
    .o({\u2_Display/add23/c21 ,\u2_Display/n594 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u21  (
    .a(\u2_Display/n570 ),
    .b(1'b1),
    .c(\u2_Display/add23/c21 ),
    .o({\u2_Display/add23/c22 ,\u2_Display/n594 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u22  (
    .a(\u2_Display/n569 ),
    .b(1'b0),
    .c(\u2_Display/add23/c22 ),
    .o({\u2_Display/add23/c23 ,\u2_Display/n594 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u23  (
    .a(\u2_Display/n568 ),
    .b(1'b0),
    .c(\u2_Display/add23/c23 ),
    .o({\u2_Display/add23/c24 ,\u2_Display/n594 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u24  (
    .a(\u2_Display/n567 ),
    .b(1'b0),
    .c(\u2_Display/add23/c24 ),
    .o({\u2_Display/add23/c25 ,\u2_Display/n594 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u25  (
    .a(\u2_Display/n566 ),
    .b(1'b0),
    .c(\u2_Display/add23/c25 ),
    .o({\u2_Display/add23/c26 ,\u2_Display/n594 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u26  (
    .a(\u2_Display/n565 ),
    .b(1'b0),
    .c(\u2_Display/add23/c26 ),
    .o({\u2_Display/add23/c27 ,\u2_Display/n594 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u27  (
    .a(\u2_Display/n564 ),
    .b(1'b1),
    .c(\u2_Display/add23/c27 ),
    .o({\u2_Display/add23/c28 ,\u2_Display/n594 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u28  (
    .a(\u2_Display/n563 ),
    .b(1'b1),
    .c(\u2_Display/add23/c28 ),
    .o({\u2_Display/add23/c29 ,\u2_Display/n594 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u29  (
    .a(\u2_Display/n562 ),
    .b(1'b1),
    .c(\u2_Display/add23/c29 ),
    .o({\u2_Display/add23/c30 ,\u2_Display/n594 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u3  (
    .a(\u2_Display/n588 ),
    .b(1'b1),
    .c(\u2_Display/add23/c3 ),
    .o({\u2_Display/add23/c4 ,\u2_Display/n594 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u30  (
    .a(\u2_Display/n561 ),
    .b(1'b1),
    .c(\u2_Display/add23/c30 ),
    .o({\u2_Display/add23/c31 ,\u2_Display/n594 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u31  (
    .a(\u2_Display/n560 ),
    .b(1'b1),
    .c(\u2_Display/add23/c31 ),
    .o({open_n1111,\u2_Display/n594 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u4  (
    .a(\u2_Display/n587 ),
    .b(1'b1),
    .c(\u2_Display/add23/c4 ),
    .o({\u2_Display/add23/c5 ,\u2_Display/n594 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u5  (
    .a(\u2_Display/n586 ),
    .b(1'b1),
    .c(\u2_Display/add23/c5 ),
    .o({\u2_Display/add23/c6 ,\u2_Display/n594 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u6  (
    .a(\u2_Display/n585 ),
    .b(1'b1),
    .c(\u2_Display/add23/c6 ),
    .o({\u2_Display/add23/c7 ,\u2_Display/n594 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u7  (
    .a(\u2_Display/n584 ),
    .b(1'b1),
    .c(\u2_Display/add23/c7 ),
    .o({\u2_Display/add23/c8 ,\u2_Display/n594 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u8  (
    .a(\u2_Display/n583 ),
    .b(1'b1),
    .c(\u2_Display/add23/c8 ),
    .o({\u2_Display/add23/c9 ,\u2_Display/n594 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add23/u9  (
    .a(\u2_Display/n582 ),
    .b(1'b1),
    .c(\u2_Display/add23/c9 ),
    .o({\u2_Display/add23/c10 ,\u2_Display/n594 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add23/ucin  (
    .a(1'b1),
    .o({\u2_Display/add23/c0 ,open_n1114}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u0  (
    .a(\u2_Display/n626 ),
    .b(1'b1),
    .c(\u2_Display/add24/c0 ),
    .o({\u2_Display/add24/c1 ,\u2_Display/n629 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u1  (
    .a(\u2_Display/n625 ),
    .b(1'b1),
    .c(\u2_Display/add24/c1 ),
    .o({\u2_Display/add24/c2 ,\u2_Display/n629 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u10  (
    .a(\u2_Display/n616 ),
    .b(1'b1),
    .c(\u2_Display/add24/c10 ),
    .o({\u2_Display/add24/c11 ,\u2_Display/n629 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u11  (
    .a(\u2_Display/n615 ),
    .b(1'b1),
    .c(\u2_Display/add24/c11 ),
    .o({\u2_Display/add24/c12 ,\u2_Display/n629 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u12  (
    .a(\u2_Display/n614 ),
    .b(1'b1),
    .c(\u2_Display/add24/c12 ),
    .o({\u2_Display/add24/c13 ,\u2_Display/n629 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u13  (
    .a(\u2_Display/n613 ),
    .b(1'b1),
    .c(\u2_Display/add24/c13 ),
    .o({\u2_Display/add24/c14 ,\u2_Display/n629 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u14  (
    .a(\u2_Display/n612 ),
    .b(1'b1),
    .c(\u2_Display/add24/c14 ),
    .o({\u2_Display/add24/c15 ,\u2_Display/n629 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u15  (
    .a(\u2_Display/n611 ),
    .b(1'b1),
    .c(\u2_Display/add24/c15 ),
    .o({\u2_Display/add24/c16 ,\u2_Display/n629 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u16  (
    .a(\u2_Display/n610 ),
    .b(1'b1),
    .c(\u2_Display/add24/c16 ),
    .o({\u2_Display/add24/c17 ,\u2_Display/n629 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u17  (
    .a(\u2_Display/n609 ),
    .b(1'b1),
    .c(\u2_Display/add24/c17 ),
    .o({\u2_Display/add24/c18 ,\u2_Display/n629 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u18  (
    .a(\u2_Display/n608 ),
    .b(1'b1),
    .c(\u2_Display/add24/c18 ),
    .o({\u2_Display/add24/c19 ,\u2_Display/n629 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u19  (
    .a(\u2_Display/n607 ),
    .b(1'b0),
    .c(\u2_Display/add24/c19 ),
    .o({\u2_Display/add24/c20 ,\u2_Display/n629 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u2  (
    .a(\u2_Display/n624 ),
    .b(1'b1),
    .c(\u2_Display/add24/c2 ),
    .o({\u2_Display/add24/c3 ,\u2_Display/n629 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u20  (
    .a(\u2_Display/n606 ),
    .b(1'b1),
    .c(\u2_Display/add24/c20 ),
    .o({\u2_Display/add24/c21 ,\u2_Display/n629 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u21  (
    .a(\u2_Display/n605 ),
    .b(1'b0),
    .c(\u2_Display/add24/c21 ),
    .o({\u2_Display/add24/c22 ,\u2_Display/n629 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u22  (
    .a(\u2_Display/n604 ),
    .b(1'b0),
    .c(\u2_Display/add24/c22 ),
    .o({\u2_Display/add24/c23 ,\u2_Display/n629 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u23  (
    .a(\u2_Display/n603 ),
    .b(1'b0),
    .c(\u2_Display/add24/c23 ),
    .o({\u2_Display/add24/c24 ,\u2_Display/n629 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u24  (
    .a(\u2_Display/n602 ),
    .b(1'b0),
    .c(\u2_Display/add24/c24 ),
    .o({\u2_Display/add24/c25 ,\u2_Display/n629 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u25  (
    .a(\u2_Display/n601 ),
    .b(1'b0),
    .c(\u2_Display/add24/c25 ),
    .o({\u2_Display/add24/c26 ,\u2_Display/n629 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u26  (
    .a(\u2_Display/n600 ),
    .b(1'b1),
    .c(\u2_Display/add24/c26 ),
    .o({\u2_Display/add24/c27 ,\u2_Display/n629 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u27  (
    .a(\u2_Display/n599 ),
    .b(1'b1),
    .c(\u2_Display/add24/c27 ),
    .o({\u2_Display/add24/c28 ,\u2_Display/n629 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u28  (
    .a(\u2_Display/n598 ),
    .b(1'b1),
    .c(\u2_Display/add24/c28 ),
    .o({\u2_Display/add24/c29 ,\u2_Display/n629 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u29  (
    .a(\u2_Display/n597 ),
    .b(1'b1),
    .c(\u2_Display/add24/c29 ),
    .o({\u2_Display/add24/c30 ,\u2_Display/n629 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u3  (
    .a(\u2_Display/n623 ),
    .b(1'b1),
    .c(\u2_Display/add24/c3 ),
    .o({\u2_Display/add24/c4 ,\u2_Display/n629 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u30  (
    .a(\u2_Display/n596 ),
    .b(1'b1),
    .c(\u2_Display/add24/c30 ),
    .o({\u2_Display/add24/c31 ,\u2_Display/n629 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u31  (
    .a(\u2_Display/n595 ),
    .b(1'b1),
    .c(\u2_Display/add24/c31 ),
    .o({open_n1115,\u2_Display/n629 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u4  (
    .a(\u2_Display/n622 ),
    .b(1'b1),
    .c(\u2_Display/add24/c4 ),
    .o({\u2_Display/add24/c5 ,\u2_Display/n629 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u5  (
    .a(\u2_Display/n621 ),
    .b(1'b1),
    .c(\u2_Display/add24/c5 ),
    .o({\u2_Display/add24/c6 ,\u2_Display/n629 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u6  (
    .a(\u2_Display/n620 ),
    .b(1'b1),
    .c(\u2_Display/add24/c6 ),
    .o({\u2_Display/add24/c7 ,\u2_Display/n629 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u7  (
    .a(\u2_Display/n619 ),
    .b(1'b1),
    .c(\u2_Display/add24/c7 ),
    .o({\u2_Display/add24/c8 ,\u2_Display/n629 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u8  (
    .a(\u2_Display/n618 ),
    .b(1'b1),
    .c(\u2_Display/add24/c8 ),
    .o({\u2_Display/add24/c9 ,\u2_Display/n629 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add24/u9  (
    .a(\u2_Display/n617 ),
    .b(1'b1),
    .c(\u2_Display/add24/c9 ),
    .o({\u2_Display/add24/c10 ,\u2_Display/n629 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add24/ucin  (
    .a(1'b1),
    .o({\u2_Display/add24/c0 ,open_n1118}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u0  (
    .a(\u2_Display/n661 ),
    .b(1'b1),
    .c(\u2_Display/add25/c0 ),
    .o({\u2_Display/add25/c1 ,\u2_Display/n664 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u1  (
    .a(\u2_Display/n660 ),
    .b(1'b1),
    .c(\u2_Display/add25/c1 ),
    .o({\u2_Display/add25/c2 ,\u2_Display/n664 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u10  (
    .a(\u2_Display/n651 ),
    .b(1'b1),
    .c(\u2_Display/add25/c10 ),
    .o({\u2_Display/add25/c11 ,\u2_Display/n664 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u11  (
    .a(\u2_Display/n650 ),
    .b(1'b1),
    .c(\u2_Display/add25/c11 ),
    .o({\u2_Display/add25/c12 ,\u2_Display/n664 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u12  (
    .a(\u2_Display/n649 ),
    .b(1'b1),
    .c(\u2_Display/add25/c12 ),
    .o({\u2_Display/add25/c13 ,\u2_Display/n664 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u13  (
    .a(\u2_Display/n648 ),
    .b(1'b1),
    .c(\u2_Display/add25/c13 ),
    .o({\u2_Display/add25/c14 ,\u2_Display/n664 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u14  (
    .a(\u2_Display/n647 ),
    .b(1'b1),
    .c(\u2_Display/add25/c14 ),
    .o({\u2_Display/add25/c15 ,\u2_Display/n664 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u15  (
    .a(\u2_Display/n646 ),
    .b(1'b1),
    .c(\u2_Display/add25/c15 ),
    .o({\u2_Display/add25/c16 ,\u2_Display/n664 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u16  (
    .a(\u2_Display/n645 ),
    .b(1'b1),
    .c(\u2_Display/add25/c16 ),
    .o({\u2_Display/add25/c17 ,\u2_Display/n664 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u17  (
    .a(\u2_Display/n644 ),
    .b(1'b1),
    .c(\u2_Display/add25/c17 ),
    .o({\u2_Display/add25/c18 ,\u2_Display/n664 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u18  (
    .a(\u2_Display/n643 ),
    .b(1'b0),
    .c(\u2_Display/add25/c18 ),
    .o({\u2_Display/add25/c19 ,\u2_Display/n664 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u19  (
    .a(\u2_Display/n642 ),
    .b(1'b1),
    .c(\u2_Display/add25/c19 ),
    .o({\u2_Display/add25/c20 ,\u2_Display/n664 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u2  (
    .a(\u2_Display/n659 ),
    .b(1'b1),
    .c(\u2_Display/add25/c2 ),
    .o({\u2_Display/add25/c3 ,\u2_Display/n664 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u20  (
    .a(\u2_Display/n641 ),
    .b(1'b0),
    .c(\u2_Display/add25/c20 ),
    .o({\u2_Display/add25/c21 ,\u2_Display/n664 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u21  (
    .a(\u2_Display/n640 ),
    .b(1'b0),
    .c(\u2_Display/add25/c21 ),
    .o({\u2_Display/add25/c22 ,\u2_Display/n664 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u22  (
    .a(\u2_Display/n639 ),
    .b(1'b0),
    .c(\u2_Display/add25/c22 ),
    .o({\u2_Display/add25/c23 ,\u2_Display/n664 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u23  (
    .a(\u2_Display/n638 ),
    .b(1'b0),
    .c(\u2_Display/add25/c23 ),
    .o({\u2_Display/add25/c24 ,\u2_Display/n664 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u24  (
    .a(\u2_Display/n637 ),
    .b(1'b0),
    .c(\u2_Display/add25/c24 ),
    .o({\u2_Display/add25/c25 ,\u2_Display/n664 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u25  (
    .a(\u2_Display/n636 ),
    .b(1'b1),
    .c(\u2_Display/add25/c25 ),
    .o({\u2_Display/add25/c26 ,\u2_Display/n664 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u26  (
    .a(\u2_Display/n635 ),
    .b(1'b1),
    .c(\u2_Display/add25/c26 ),
    .o({\u2_Display/add25/c27 ,\u2_Display/n664 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u27  (
    .a(\u2_Display/n634 ),
    .b(1'b1),
    .c(\u2_Display/add25/c27 ),
    .o({\u2_Display/add25/c28 ,\u2_Display/n664 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u28  (
    .a(\u2_Display/n633 ),
    .b(1'b1),
    .c(\u2_Display/add25/c28 ),
    .o({\u2_Display/add25/c29 ,\u2_Display/n664 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u29  (
    .a(\u2_Display/n632 ),
    .b(1'b1),
    .c(\u2_Display/add25/c29 ),
    .o({\u2_Display/add25/c30 ,\u2_Display/n664 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u3  (
    .a(\u2_Display/n658 ),
    .b(1'b1),
    .c(\u2_Display/add25/c3 ),
    .o({\u2_Display/add25/c4 ,\u2_Display/n664 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u30  (
    .a(\u2_Display/n631 ),
    .b(1'b1),
    .c(\u2_Display/add25/c30 ),
    .o({\u2_Display/add25/c31 ,\u2_Display/n664 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u31  (
    .a(\u2_Display/n630 ),
    .b(1'b1),
    .c(\u2_Display/add25/c31 ),
    .o({open_n1119,\u2_Display/n664 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u4  (
    .a(\u2_Display/n657 ),
    .b(1'b1),
    .c(\u2_Display/add25/c4 ),
    .o({\u2_Display/add25/c5 ,\u2_Display/n664 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u5  (
    .a(\u2_Display/n656 ),
    .b(1'b1),
    .c(\u2_Display/add25/c5 ),
    .o({\u2_Display/add25/c6 ,\u2_Display/n664 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u6  (
    .a(\u2_Display/n655 ),
    .b(1'b1),
    .c(\u2_Display/add25/c6 ),
    .o({\u2_Display/add25/c7 ,\u2_Display/n664 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u7  (
    .a(\u2_Display/n654 ),
    .b(1'b1),
    .c(\u2_Display/add25/c7 ),
    .o({\u2_Display/add25/c8 ,\u2_Display/n664 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u8  (
    .a(\u2_Display/n653 ),
    .b(1'b1),
    .c(\u2_Display/add25/c8 ),
    .o({\u2_Display/add25/c9 ,\u2_Display/n664 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add25/u9  (
    .a(\u2_Display/n652 ),
    .b(1'b1),
    .c(\u2_Display/add25/c9 ),
    .o({\u2_Display/add25/c10 ,\u2_Display/n664 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add25/ucin  (
    .a(1'b1),
    .o({\u2_Display/add25/c0 ,open_n1122}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u0  (
    .a(\u2_Display/n696 ),
    .b(1'b1),
    .c(\u2_Display/add26/c0 ),
    .o({\u2_Display/add26/c1 ,\u2_Display/n699 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u1  (
    .a(\u2_Display/n695 ),
    .b(1'b1),
    .c(\u2_Display/add26/c1 ),
    .o({\u2_Display/add26/c2 ,\u2_Display/n699 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u10  (
    .a(\u2_Display/n686 ),
    .b(1'b1),
    .c(\u2_Display/add26/c10 ),
    .o({\u2_Display/add26/c11 ,\u2_Display/n699 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u11  (
    .a(\u2_Display/n685 ),
    .b(1'b1),
    .c(\u2_Display/add26/c11 ),
    .o({\u2_Display/add26/c12 ,\u2_Display/n699 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u12  (
    .a(\u2_Display/n684 ),
    .b(1'b1),
    .c(\u2_Display/add26/c12 ),
    .o({\u2_Display/add26/c13 ,\u2_Display/n699 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u13  (
    .a(\u2_Display/n683 ),
    .b(1'b1),
    .c(\u2_Display/add26/c13 ),
    .o({\u2_Display/add26/c14 ,\u2_Display/n699 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u14  (
    .a(\u2_Display/n682 ),
    .b(1'b1),
    .c(\u2_Display/add26/c14 ),
    .o({\u2_Display/add26/c15 ,\u2_Display/n699 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u15  (
    .a(\u2_Display/n681 ),
    .b(1'b1),
    .c(\u2_Display/add26/c15 ),
    .o({\u2_Display/add26/c16 ,\u2_Display/n699 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u16  (
    .a(\u2_Display/n680 ),
    .b(1'b1),
    .c(\u2_Display/add26/c16 ),
    .o({\u2_Display/add26/c17 ,\u2_Display/n699 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u17  (
    .a(\u2_Display/n679 ),
    .b(1'b0),
    .c(\u2_Display/add26/c17 ),
    .o({\u2_Display/add26/c18 ,\u2_Display/n699 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u18  (
    .a(\u2_Display/n678 ),
    .b(1'b1),
    .c(\u2_Display/add26/c18 ),
    .o({\u2_Display/add26/c19 ,\u2_Display/n699 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u19  (
    .a(\u2_Display/n677 ),
    .b(1'b0),
    .c(\u2_Display/add26/c19 ),
    .o({\u2_Display/add26/c20 ,\u2_Display/n699 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u2  (
    .a(\u2_Display/n694 ),
    .b(1'b1),
    .c(\u2_Display/add26/c2 ),
    .o({\u2_Display/add26/c3 ,\u2_Display/n699 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u20  (
    .a(\u2_Display/n676 ),
    .b(1'b0),
    .c(\u2_Display/add26/c20 ),
    .o({\u2_Display/add26/c21 ,\u2_Display/n699 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u21  (
    .a(\u2_Display/n675 ),
    .b(1'b0),
    .c(\u2_Display/add26/c21 ),
    .o({\u2_Display/add26/c22 ,\u2_Display/n699 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u22  (
    .a(\u2_Display/n674 ),
    .b(1'b0),
    .c(\u2_Display/add26/c22 ),
    .o({\u2_Display/add26/c23 ,\u2_Display/n699 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u23  (
    .a(\u2_Display/n673 ),
    .b(1'b0),
    .c(\u2_Display/add26/c23 ),
    .o({\u2_Display/add26/c24 ,\u2_Display/n699 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u24  (
    .a(\u2_Display/n672 ),
    .b(1'b1),
    .c(\u2_Display/add26/c24 ),
    .o({\u2_Display/add26/c25 ,\u2_Display/n699 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u25  (
    .a(\u2_Display/n671 ),
    .b(1'b1),
    .c(\u2_Display/add26/c25 ),
    .o({\u2_Display/add26/c26 ,\u2_Display/n699 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u26  (
    .a(\u2_Display/n670 ),
    .b(1'b1),
    .c(\u2_Display/add26/c26 ),
    .o({\u2_Display/add26/c27 ,\u2_Display/n699 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u27  (
    .a(\u2_Display/n669 ),
    .b(1'b1),
    .c(\u2_Display/add26/c27 ),
    .o({\u2_Display/add26/c28 ,\u2_Display/n699 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u28  (
    .a(\u2_Display/n668 ),
    .b(1'b1),
    .c(\u2_Display/add26/c28 ),
    .o({\u2_Display/add26/c29 ,\u2_Display/n699 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u29  (
    .a(\u2_Display/n667 ),
    .b(1'b1),
    .c(\u2_Display/add26/c29 ),
    .o({\u2_Display/add26/c30 ,\u2_Display/n699 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u3  (
    .a(\u2_Display/n693 ),
    .b(1'b1),
    .c(\u2_Display/add26/c3 ),
    .o({\u2_Display/add26/c4 ,\u2_Display/n699 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u30  (
    .a(\u2_Display/n666 ),
    .b(1'b1),
    .c(\u2_Display/add26/c30 ),
    .o({\u2_Display/add26/c31 ,\u2_Display/n699 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u31  (
    .a(\u2_Display/n665 ),
    .b(1'b1),
    .c(\u2_Display/add26/c31 ),
    .o({open_n1123,\u2_Display/n699 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u4  (
    .a(\u2_Display/n692 ),
    .b(1'b1),
    .c(\u2_Display/add26/c4 ),
    .o({\u2_Display/add26/c5 ,\u2_Display/n699 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u5  (
    .a(\u2_Display/n691 ),
    .b(1'b1),
    .c(\u2_Display/add26/c5 ),
    .o({\u2_Display/add26/c6 ,\u2_Display/n699 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u6  (
    .a(\u2_Display/n690 ),
    .b(1'b1),
    .c(\u2_Display/add26/c6 ),
    .o({\u2_Display/add26/c7 ,\u2_Display/n699 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u7  (
    .a(\u2_Display/n689 ),
    .b(1'b1),
    .c(\u2_Display/add26/c7 ),
    .o({\u2_Display/add26/c8 ,\u2_Display/n699 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u8  (
    .a(\u2_Display/n688 ),
    .b(1'b1),
    .c(\u2_Display/add26/c8 ),
    .o({\u2_Display/add26/c9 ,\u2_Display/n699 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add26/u9  (
    .a(\u2_Display/n687 ),
    .b(1'b1),
    .c(\u2_Display/add26/c9 ),
    .o({\u2_Display/add26/c10 ,\u2_Display/n699 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add26/ucin  (
    .a(1'b1),
    .o({\u2_Display/add26/c0 ,open_n1126}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u0  (
    .a(\u2_Display/n731 ),
    .b(1'b1),
    .c(\u2_Display/add27/c0 ),
    .o({\u2_Display/add27/c1 ,\u2_Display/n734 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u1  (
    .a(\u2_Display/n730 ),
    .b(1'b1),
    .c(\u2_Display/add27/c1 ),
    .o({\u2_Display/add27/c2 ,\u2_Display/n734 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u10  (
    .a(\u2_Display/n721 ),
    .b(1'b1),
    .c(\u2_Display/add27/c10 ),
    .o({\u2_Display/add27/c11 ,\u2_Display/n734 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u11  (
    .a(\u2_Display/n720 ),
    .b(1'b1),
    .c(\u2_Display/add27/c11 ),
    .o({\u2_Display/add27/c12 ,\u2_Display/n734 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u12  (
    .a(\u2_Display/n719 ),
    .b(1'b1),
    .c(\u2_Display/add27/c12 ),
    .o({\u2_Display/add27/c13 ,\u2_Display/n734 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u13  (
    .a(\u2_Display/n718 ),
    .b(1'b1),
    .c(\u2_Display/add27/c13 ),
    .o({\u2_Display/add27/c14 ,\u2_Display/n734 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u14  (
    .a(\u2_Display/n717 ),
    .b(1'b1),
    .c(\u2_Display/add27/c14 ),
    .o({\u2_Display/add27/c15 ,\u2_Display/n734 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u15  (
    .a(\u2_Display/n716 ),
    .b(1'b1),
    .c(\u2_Display/add27/c15 ),
    .o({\u2_Display/add27/c16 ,\u2_Display/n734 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u16  (
    .a(\u2_Display/n715 ),
    .b(1'b0),
    .c(\u2_Display/add27/c16 ),
    .o({\u2_Display/add27/c17 ,\u2_Display/n734 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u17  (
    .a(\u2_Display/n714 ),
    .b(1'b1),
    .c(\u2_Display/add27/c17 ),
    .o({\u2_Display/add27/c18 ,\u2_Display/n734 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u18  (
    .a(\u2_Display/n713 ),
    .b(1'b0),
    .c(\u2_Display/add27/c18 ),
    .o({\u2_Display/add27/c19 ,\u2_Display/n734 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u19  (
    .a(\u2_Display/n712 ),
    .b(1'b0),
    .c(\u2_Display/add27/c19 ),
    .o({\u2_Display/add27/c20 ,\u2_Display/n734 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u2  (
    .a(\u2_Display/n729 ),
    .b(1'b1),
    .c(\u2_Display/add27/c2 ),
    .o({\u2_Display/add27/c3 ,\u2_Display/n734 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u20  (
    .a(\u2_Display/n711 ),
    .b(1'b0),
    .c(\u2_Display/add27/c20 ),
    .o({\u2_Display/add27/c21 ,\u2_Display/n734 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u21  (
    .a(\u2_Display/n710 ),
    .b(1'b0),
    .c(\u2_Display/add27/c21 ),
    .o({\u2_Display/add27/c22 ,\u2_Display/n734 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u22  (
    .a(\u2_Display/n709 ),
    .b(1'b0),
    .c(\u2_Display/add27/c22 ),
    .o({\u2_Display/add27/c23 ,\u2_Display/n734 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u23  (
    .a(\u2_Display/n708 ),
    .b(1'b1),
    .c(\u2_Display/add27/c23 ),
    .o({\u2_Display/add27/c24 ,\u2_Display/n734 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u24  (
    .a(\u2_Display/n707 ),
    .b(1'b1),
    .c(\u2_Display/add27/c24 ),
    .o({\u2_Display/add27/c25 ,\u2_Display/n734 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u25  (
    .a(\u2_Display/n706 ),
    .b(1'b1),
    .c(\u2_Display/add27/c25 ),
    .o({\u2_Display/add27/c26 ,\u2_Display/n734 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u26  (
    .a(\u2_Display/n705 ),
    .b(1'b1),
    .c(\u2_Display/add27/c26 ),
    .o({\u2_Display/add27/c27 ,\u2_Display/n734 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u27  (
    .a(\u2_Display/n704 ),
    .b(1'b1),
    .c(\u2_Display/add27/c27 ),
    .o({\u2_Display/add27/c28 ,\u2_Display/n734 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u28  (
    .a(\u2_Display/n703 ),
    .b(1'b1),
    .c(\u2_Display/add27/c28 ),
    .o({\u2_Display/add27/c29 ,\u2_Display/n734 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u29  (
    .a(\u2_Display/n702 ),
    .b(1'b1),
    .c(\u2_Display/add27/c29 ),
    .o({\u2_Display/add27/c30 ,\u2_Display/n734 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u3  (
    .a(\u2_Display/n728 ),
    .b(1'b1),
    .c(\u2_Display/add27/c3 ),
    .o({\u2_Display/add27/c4 ,\u2_Display/n734 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u30  (
    .a(\u2_Display/n701 ),
    .b(1'b1),
    .c(\u2_Display/add27/c30 ),
    .o({\u2_Display/add27/c31 ,\u2_Display/n734 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u31  (
    .a(\u2_Display/n700 ),
    .b(1'b1),
    .c(\u2_Display/add27/c31 ),
    .o({open_n1127,\u2_Display/n734 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u4  (
    .a(\u2_Display/n727 ),
    .b(1'b1),
    .c(\u2_Display/add27/c4 ),
    .o({\u2_Display/add27/c5 ,\u2_Display/n734 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u5  (
    .a(\u2_Display/n726 ),
    .b(1'b1),
    .c(\u2_Display/add27/c5 ),
    .o({\u2_Display/add27/c6 ,\u2_Display/n734 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u6  (
    .a(\u2_Display/n725 ),
    .b(1'b1),
    .c(\u2_Display/add27/c6 ),
    .o({\u2_Display/add27/c7 ,\u2_Display/n734 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u7  (
    .a(\u2_Display/n724 ),
    .b(1'b1),
    .c(\u2_Display/add27/c7 ),
    .o({\u2_Display/add27/c8 ,\u2_Display/n734 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u8  (
    .a(\u2_Display/n723 ),
    .b(1'b1),
    .c(\u2_Display/add27/c8 ),
    .o({\u2_Display/add27/c9 ,\u2_Display/n734 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add27/u9  (
    .a(\u2_Display/n722 ),
    .b(1'b1),
    .c(\u2_Display/add27/c9 ),
    .o({\u2_Display/add27/c10 ,\u2_Display/n734 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add27/ucin  (
    .a(1'b1),
    .o({\u2_Display/add27/c0 ,open_n1130}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u0  (
    .a(\u2_Display/n766 ),
    .b(1'b1),
    .c(\u2_Display/add28/c0 ),
    .o({\u2_Display/add28/c1 ,\u2_Display/n769 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u1  (
    .a(\u2_Display/n765 ),
    .b(1'b1),
    .c(\u2_Display/add28/c1 ),
    .o({\u2_Display/add28/c2 ,\u2_Display/n769 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u10  (
    .a(\u2_Display/n756 ),
    .b(1'b1),
    .c(\u2_Display/add28/c10 ),
    .o({\u2_Display/add28/c11 ,\u2_Display/n769 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u11  (
    .a(\u2_Display/n755 ),
    .b(1'b1),
    .c(\u2_Display/add28/c11 ),
    .o({\u2_Display/add28/c12 ,\u2_Display/n769 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u12  (
    .a(\u2_Display/n754 ),
    .b(1'b1),
    .c(\u2_Display/add28/c12 ),
    .o({\u2_Display/add28/c13 ,\u2_Display/n769 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u13  (
    .a(\u2_Display/n753 ),
    .b(1'b1),
    .c(\u2_Display/add28/c13 ),
    .o({\u2_Display/add28/c14 ,\u2_Display/n769 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u14  (
    .a(\u2_Display/n752 ),
    .b(1'b1),
    .c(\u2_Display/add28/c14 ),
    .o({\u2_Display/add28/c15 ,\u2_Display/n769 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u15  (
    .a(\u2_Display/n751 ),
    .b(1'b0),
    .c(\u2_Display/add28/c15 ),
    .o({\u2_Display/add28/c16 ,\u2_Display/n769 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u16  (
    .a(\u2_Display/n750 ),
    .b(1'b1),
    .c(\u2_Display/add28/c16 ),
    .o({\u2_Display/add28/c17 ,\u2_Display/n769 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u17  (
    .a(\u2_Display/n749 ),
    .b(1'b0),
    .c(\u2_Display/add28/c17 ),
    .o({\u2_Display/add28/c18 ,\u2_Display/n769 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u18  (
    .a(\u2_Display/n748 ),
    .b(1'b0),
    .c(\u2_Display/add28/c18 ),
    .o({\u2_Display/add28/c19 ,\u2_Display/n769 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u19  (
    .a(\u2_Display/n747 ),
    .b(1'b0),
    .c(\u2_Display/add28/c19 ),
    .o({\u2_Display/add28/c20 ,\u2_Display/n769 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u2  (
    .a(\u2_Display/n764 ),
    .b(1'b1),
    .c(\u2_Display/add28/c2 ),
    .o({\u2_Display/add28/c3 ,\u2_Display/n769 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u20  (
    .a(\u2_Display/n746 ),
    .b(1'b0),
    .c(\u2_Display/add28/c20 ),
    .o({\u2_Display/add28/c21 ,\u2_Display/n769 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u21  (
    .a(\u2_Display/n745 ),
    .b(1'b0),
    .c(\u2_Display/add28/c21 ),
    .o({\u2_Display/add28/c22 ,\u2_Display/n769 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u22  (
    .a(\u2_Display/n744 ),
    .b(1'b1),
    .c(\u2_Display/add28/c22 ),
    .o({\u2_Display/add28/c23 ,\u2_Display/n769 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u23  (
    .a(\u2_Display/n743 ),
    .b(1'b1),
    .c(\u2_Display/add28/c23 ),
    .o({\u2_Display/add28/c24 ,\u2_Display/n769 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u24  (
    .a(\u2_Display/n742 ),
    .b(1'b1),
    .c(\u2_Display/add28/c24 ),
    .o({\u2_Display/add28/c25 ,\u2_Display/n769 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u25  (
    .a(\u2_Display/n741 ),
    .b(1'b1),
    .c(\u2_Display/add28/c25 ),
    .o({\u2_Display/add28/c26 ,\u2_Display/n769 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u26  (
    .a(\u2_Display/n740 ),
    .b(1'b1),
    .c(\u2_Display/add28/c26 ),
    .o({\u2_Display/add28/c27 ,\u2_Display/n769 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u27  (
    .a(\u2_Display/n739 ),
    .b(1'b1),
    .c(\u2_Display/add28/c27 ),
    .o({\u2_Display/add28/c28 ,\u2_Display/n769 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u28  (
    .a(\u2_Display/n738 ),
    .b(1'b1),
    .c(\u2_Display/add28/c28 ),
    .o({\u2_Display/add28/c29 ,\u2_Display/n769 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u29  (
    .a(\u2_Display/n737 ),
    .b(1'b1),
    .c(\u2_Display/add28/c29 ),
    .o({\u2_Display/add28/c30 ,\u2_Display/n769 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u3  (
    .a(\u2_Display/n763 ),
    .b(1'b1),
    .c(\u2_Display/add28/c3 ),
    .o({\u2_Display/add28/c4 ,\u2_Display/n769 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u30  (
    .a(\u2_Display/n736 ),
    .b(1'b1),
    .c(\u2_Display/add28/c30 ),
    .o({\u2_Display/add28/c31 ,\u2_Display/n769 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u31  (
    .a(\u2_Display/n735 ),
    .b(1'b1),
    .c(\u2_Display/add28/c31 ),
    .o({open_n1131,\u2_Display/n769 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u4  (
    .a(\u2_Display/n762 ),
    .b(1'b1),
    .c(\u2_Display/add28/c4 ),
    .o({\u2_Display/add28/c5 ,\u2_Display/n769 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u5  (
    .a(\u2_Display/n761 ),
    .b(1'b1),
    .c(\u2_Display/add28/c5 ),
    .o({\u2_Display/add28/c6 ,\u2_Display/n769 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u6  (
    .a(\u2_Display/n760 ),
    .b(1'b1),
    .c(\u2_Display/add28/c6 ),
    .o({\u2_Display/add28/c7 ,\u2_Display/n769 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u7  (
    .a(\u2_Display/n759 ),
    .b(1'b1),
    .c(\u2_Display/add28/c7 ),
    .o({\u2_Display/add28/c8 ,\u2_Display/n769 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u8  (
    .a(\u2_Display/n758 ),
    .b(1'b1),
    .c(\u2_Display/add28/c8 ),
    .o({\u2_Display/add28/c9 ,\u2_Display/n769 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add28/u9  (
    .a(\u2_Display/n757 ),
    .b(1'b1),
    .c(\u2_Display/add28/c9 ),
    .o({\u2_Display/add28/c10 ,\u2_Display/n769 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add28/ucin  (
    .a(1'b1),
    .o({\u2_Display/add28/c0 ,open_n1134}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u0  (
    .a(\u2_Display/n801 ),
    .b(1'b1),
    .c(\u2_Display/add29/c0 ),
    .o({\u2_Display/add29/c1 ,\u2_Display/n804 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u1  (
    .a(\u2_Display/n800 ),
    .b(1'b1),
    .c(\u2_Display/add29/c1 ),
    .o({\u2_Display/add29/c2 ,\u2_Display/n804 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u10  (
    .a(\u2_Display/n791 ),
    .b(1'b1),
    .c(\u2_Display/add29/c10 ),
    .o({\u2_Display/add29/c11 ,\u2_Display/n804 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u11  (
    .a(\u2_Display/n790 ),
    .b(1'b1),
    .c(\u2_Display/add29/c11 ),
    .o({\u2_Display/add29/c12 ,\u2_Display/n804 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u12  (
    .a(\u2_Display/n789 ),
    .b(1'b1),
    .c(\u2_Display/add29/c12 ),
    .o({\u2_Display/add29/c13 ,\u2_Display/n804 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u13  (
    .a(\u2_Display/n788 ),
    .b(1'b1),
    .c(\u2_Display/add29/c13 ),
    .o({\u2_Display/add29/c14 ,\u2_Display/n804 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u14  (
    .a(\u2_Display/n787 ),
    .b(1'b0),
    .c(\u2_Display/add29/c14 ),
    .o({\u2_Display/add29/c15 ,\u2_Display/n804 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u15  (
    .a(\u2_Display/n786 ),
    .b(1'b1),
    .c(\u2_Display/add29/c15 ),
    .o({\u2_Display/add29/c16 ,\u2_Display/n804 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u16  (
    .a(\u2_Display/n785 ),
    .b(1'b0),
    .c(\u2_Display/add29/c16 ),
    .o({\u2_Display/add29/c17 ,\u2_Display/n804 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u17  (
    .a(\u2_Display/n784 ),
    .b(1'b0),
    .c(\u2_Display/add29/c17 ),
    .o({\u2_Display/add29/c18 ,\u2_Display/n804 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u18  (
    .a(\u2_Display/n783 ),
    .b(1'b0),
    .c(\u2_Display/add29/c18 ),
    .o({\u2_Display/add29/c19 ,\u2_Display/n804 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u19  (
    .a(\u2_Display/n782 ),
    .b(1'b0),
    .c(\u2_Display/add29/c19 ),
    .o({\u2_Display/add29/c20 ,\u2_Display/n804 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u2  (
    .a(\u2_Display/n799 ),
    .b(1'b1),
    .c(\u2_Display/add29/c2 ),
    .o({\u2_Display/add29/c3 ,\u2_Display/n804 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u20  (
    .a(\u2_Display/n781 ),
    .b(1'b0),
    .c(\u2_Display/add29/c20 ),
    .o({\u2_Display/add29/c21 ,\u2_Display/n804 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u21  (
    .a(\u2_Display/n780 ),
    .b(1'b1),
    .c(\u2_Display/add29/c21 ),
    .o({\u2_Display/add29/c22 ,\u2_Display/n804 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u22  (
    .a(\u2_Display/n779 ),
    .b(1'b1),
    .c(\u2_Display/add29/c22 ),
    .o({\u2_Display/add29/c23 ,\u2_Display/n804 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u23  (
    .a(\u2_Display/n778 ),
    .b(1'b1),
    .c(\u2_Display/add29/c23 ),
    .o({\u2_Display/add29/c24 ,\u2_Display/n804 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u24  (
    .a(\u2_Display/n777 ),
    .b(1'b1),
    .c(\u2_Display/add29/c24 ),
    .o({\u2_Display/add29/c25 ,\u2_Display/n804 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u25  (
    .a(\u2_Display/n776 ),
    .b(1'b1),
    .c(\u2_Display/add29/c25 ),
    .o({\u2_Display/add29/c26 ,\u2_Display/n804 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u26  (
    .a(\u2_Display/n775 ),
    .b(1'b1),
    .c(\u2_Display/add29/c26 ),
    .o({\u2_Display/add29/c27 ,\u2_Display/n804 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u27  (
    .a(\u2_Display/n774 ),
    .b(1'b1),
    .c(\u2_Display/add29/c27 ),
    .o({\u2_Display/add29/c28 ,\u2_Display/n804 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u28  (
    .a(\u2_Display/n773 ),
    .b(1'b1),
    .c(\u2_Display/add29/c28 ),
    .o({\u2_Display/add29/c29 ,\u2_Display/n804 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u29  (
    .a(\u2_Display/n772 ),
    .b(1'b1),
    .c(\u2_Display/add29/c29 ),
    .o({\u2_Display/add29/c30 ,\u2_Display/n804 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u3  (
    .a(\u2_Display/n798 ),
    .b(1'b1),
    .c(\u2_Display/add29/c3 ),
    .o({\u2_Display/add29/c4 ,\u2_Display/n804 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u30  (
    .a(\u2_Display/n771 ),
    .b(1'b1),
    .c(\u2_Display/add29/c30 ),
    .o({\u2_Display/add29/c31 ,\u2_Display/n804 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u31  (
    .a(\u2_Display/n770 ),
    .b(1'b1),
    .c(\u2_Display/add29/c31 ),
    .o({open_n1135,\u2_Display/n804 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u4  (
    .a(\u2_Display/n797 ),
    .b(1'b1),
    .c(\u2_Display/add29/c4 ),
    .o({\u2_Display/add29/c5 ,\u2_Display/n804 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u5  (
    .a(\u2_Display/n796 ),
    .b(1'b1),
    .c(\u2_Display/add29/c5 ),
    .o({\u2_Display/add29/c6 ,\u2_Display/n804 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u6  (
    .a(\u2_Display/n795 ),
    .b(1'b1),
    .c(\u2_Display/add29/c6 ),
    .o({\u2_Display/add29/c7 ,\u2_Display/n804 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u7  (
    .a(\u2_Display/n794 ),
    .b(1'b1),
    .c(\u2_Display/add29/c7 ),
    .o({\u2_Display/add29/c8 ,\u2_Display/n804 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u8  (
    .a(\u2_Display/n793 ),
    .b(1'b1),
    .c(\u2_Display/add29/c8 ),
    .o({\u2_Display/add29/c9 ,\u2_Display/n804 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add29/u9  (
    .a(\u2_Display/n792 ),
    .b(1'b1),
    .c(\u2_Display/add29/c9 ),
    .o({\u2_Display/add29/c10 ,\u2_Display/n804 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add29/ucin  (
    .a(1'b1),
    .o({\u2_Display/add29/c0 ,open_n1138}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add2_2/u0  (
    .a(1'b1),
    .b(\u2_Display/i [8]),
    .c(\u2_Display/add2_2/c0 ),
    .o({\u2_Display/add2_2/c1 ,\u2_Display/n43 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add2_2/u1  (
    .a(1'b0),
    .b(\u2_Display/i [9]),
    .c(\u2_Display/add2_2/c1 ),
    .o({\u2_Display/add2_2/c2 ,\u2_Display/n43 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add2_2/u2  (
    .a(1'b1),
    .b(\u2_Display/i [10]),
    .c(\u2_Display/add2_2/c2 ),
    .o({\u2_Display/add2_2/c3 ,\u2_Display/n43 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add2_2/ucin  (
    .a(1'b0),
    .o({\u2_Display/add2_2/c0 ,open_n1141}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add2_2/ucout  (
    .c(\u2_Display/add2_2/c3 ),
    .o({open_n1144,\u2_Display/add2_2_co }));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u0  (
    .a(\u2_Display/n836 ),
    .b(1'b1),
    .c(\u2_Display/add30/c0 ),
    .o({\u2_Display/add30/c1 ,\u2_Display/n839 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u1  (
    .a(\u2_Display/n835 ),
    .b(1'b1),
    .c(\u2_Display/add30/c1 ),
    .o({\u2_Display/add30/c2 ,\u2_Display/n839 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u10  (
    .a(\u2_Display/n826 ),
    .b(1'b1),
    .c(\u2_Display/add30/c10 ),
    .o({\u2_Display/add30/c11 ,\u2_Display/n839 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u11  (
    .a(\u2_Display/n825 ),
    .b(1'b1),
    .c(\u2_Display/add30/c11 ),
    .o({\u2_Display/add30/c12 ,\u2_Display/n839 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u12  (
    .a(\u2_Display/n824 ),
    .b(1'b1),
    .c(\u2_Display/add30/c12 ),
    .o({\u2_Display/add30/c13 ,\u2_Display/n839 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u13  (
    .a(\u2_Display/n823 ),
    .b(1'b0),
    .c(\u2_Display/add30/c13 ),
    .o({\u2_Display/add30/c14 ,\u2_Display/n839 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u14  (
    .a(\u2_Display/n822 ),
    .b(1'b1),
    .c(\u2_Display/add30/c14 ),
    .o({\u2_Display/add30/c15 ,\u2_Display/n839 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u15  (
    .a(\u2_Display/n821 ),
    .b(1'b0),
    .c(\u2_Display/add30/c15 ),
    .o({\u2_Display/add30/c16 ,\u2_Display/n839 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u16  (
    .a(\u2_Display/n820 ),
    .b(1'b0),
    .c(\u2_Display/add30/c16 ),
    .o({\u2_Display/add30/c17 ,\u2_Display/n839 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u17  (
    .a(\u2_Display/n819 ),
    .b(1'b0),
    .c(\u2_Display/add30/c17 ),
    .o({\u2_Display/add30/c18 ,\u2_Display/n839 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u18  (
    .a(\u2_Display/n818 ),
    .b(1'b0),
    .c(\u2_Display/add30/c18 ),
    .o({\u2_Display/add30/c19 ,\u2_Display/n839 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u19  (
    .a(\u2_Display/n817 ),
    .b(1'b0),
    .c(\u2_Display/add30/c19 ),
    .o({\u2_Display/add30/c20 ,\u2_Display/n839 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u2  (
    .a(\u2_Display/n834 ),
    .b(1'b1),
    .c(\u2_Display/add30/c2 ),
    .o({\u2_Display/add30/c3 ,\u2_Display/n839 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u20  (
    .a(\u2_Display/n816 ),
    .b(1'b1),
    .c(\u2_Display/add30/c20 ),
    .o({\u2_Display/add30/c21 ,\u2_Display/n839 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u21  (
    .a(\u2_Display/n815 ),
    .b(1'b1),
    .c(\u2_Display/add30/c21 ),
    .o({\u2_Display/add30/c22 ,\u2_Display/n839 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u22  (
    .a(\u2_Display/n814 ),
    .b(1'b1),
    .c(\u2_Display/add30/c22 ),
    .o({\u2_Display/add30/c23 ,\u2_Display/n839 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u23  (
    .a(\u2_Display/n813 ),
    .b(1'b1),
    .c(\u2_Display/add30/c23 ),
    .o({\u2_Display/add30/c24 ,\u2_Display/n839 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u24  (
    .a(\u2_Display/n812 ),
    .b(1'b1),
    .c(\u2_Display/add30/c24 ),
    .o({\u2_Display/add30/c25 ,\u2_Display/n839 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u25  (
    .a(\u2_Display/n811 ),
    .b(1'b1),
    .c(\u2_Display/add30/c25 ),
    .o({\u2_Display/add30/c26 ,\u2_Display/n839 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u26  (
    .a(\u2_Display/n810 ),
    .b(1'b1),
    .c(\u2_Display/add30/c26 ),
    .o({\u2_Display/add30/c27 ,\u2_Display/n839 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u27  (
    .a(\u2_Display/n809 ),
    .b(1'b1),
    .c(\u2_Display/add30/c27 ),
    .o({\u2_Display/add30/c28 ,\u2_Display/n839 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u28  (
    .a(\u2_Display/n808 ),
    .b(1'b1),
    .c(\u2_Display/add30/c28 ),
    .o({\u2_Display/add30/c29 ,\u2_Display/n839 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u29  (
    .a(\u2_Display/n807 ),
    .b(1'b1),
    .c(\u2_Display/add30/c29 ),
    .o({\u2_Display/add30/c30 ,\u2_Display/n839 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u3  (
    .a(\u2_Display/n833 ),
    .b(1'b1),
    .c(\u2_Display/add30/c3 ),
    .o({\u2_Display/add30/c4 ,\u2_Display/n839 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u30  (
    .a(\u2_Display/n806 ),
    .b(1'b1),
    .c(\u2_Display/add30/c30 ),
    .o({\u2_Display/add30/c31 ,\u2_Display/n839 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u31  (
    .a(\u2_Display/n805 ),
    .b(1'b1),
    .c(\u2_Display/add30/c31 ),
    .o({open_n1145,\u2_Display/n839 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u4  (
    .a(\u2_Display/n832 ),
    .b(1'b1),
    .c(\u2_Display/add30/c4 ),
    .o({\u2_Display/add30/c5 ,\u2_Display/n839 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u5  (
    .a(\u2_Display/n831 ),
    .b(1'b1),
    .c(\u2_Display/add30/c5 ),
    .o({\u2_Display/add30/c6 ,\u2_Display/n839 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u6  (
    .a(\u2_Display/n830 ),
    .b(1'b1),
    .c(\u2_Display/add30/c6 ),
    .o({\u2_Display/add30/c7 ,\u2_Display/n839 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u7  (
    .a(\u2_Display/n829 ),
    .b(1'b1),
    .c(\u2_Display/add30/c7 ),
    .o({\u2_Display/add30/c8 ,\u2_Display/n839 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u8  (
    .a(\u2_Display/n828 ),
    .b(1'b1),
    .c(\u2_Display/add30/c8 ),
    .o({\u2_Display/add30/c9 ,\u2_Display/n839 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add30/u9  (
    .a(\u2_Display/n827 ),
    .b(1'b1),
    .c(\u2_Display/add30/c9 ),
    .o({\u2_Display/add30/c10 ,\u2_Display/n839 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add30/ucin  (
    .a(1'b1),
    .o({\u2_Display/add30/c0 ,open_n1148}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u0  (
    .a(\u2_Display/n871 ),
    .b(1'b1),
    .c(\u2_Display/add31/c0 ),
    .o({\u2_Display/add31/c1 ,\u2_Display/n874 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u1  (
    .a(\u2_Display/n870 ),
    .b(1'b1),
    .c(\u2_Display/add31/c1 ),
    .o({\u2_Display/add31/c2 ,\u2_Display/n874 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u10  (
    .a(\u2_Display/n861 ),
    .b(1'b1),
    .c(\u2_Display/add31/c10 ),
    .o({\u2_Display/add31/c11 ,\u2_Display/n874 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u11  (
    .a(\u2_Display/n860 ),
    .b(1'b1),
    .c(\u2_Display/add31/c11 ),
    .o({\u2_Display/add31/c12 ,\u2_Display/n874 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u12  (
    .a(\u2_Display/n859 ),
    .b(1'b0),
    .c(\u2_Display/add31/c12 ),
    .o({\u2_Display/add31/c13 ,\u2_Display/n874 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u13  (
    .a(\u2_Display/n858 ),
    .b(1'b1),
    .c(\u2_Display/add31/c13 ),
    .o({\u2_Display/add31/c14 ,\u2_Display/n874 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u14  (
    .a(\u2_Display/n857 ),
    .b(1'b0),
    .c(\u2_Display/add31/c14 ),
    .o({\u2_Display/add31/c15 ,\u2_Display/n874 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u15  (
    .a(\u2_Display/n856 ),
    .b(1'b0),
    .c(\u2_Display/add31/c15 ),
    .o({\u2_Display/add31/c16 ,\u2_Display/n874 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u16  (
    .a(\u2_Display/n855 ),
    .b(1'b0),
    .c(\u2_Display/add31/c16 ),
    .o({\u2_Display/add31/c17 ,\u2_Display/n874 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u17  (
    .a(\u2_Display/n854 ),
    .b(1'b0),
    .c(\u2_Display/add31/c17 ),
    .o({\u2_Display/add31/c18 ,\u2_Display/n874 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u18  (
    .a(\u2_Display/n853 ),
    .b(1'b0),
    .c(\u2_Display/add31/c18 ),
    .o({\u2_Display/add31/c19 ,\u2_Display/n874 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u19  (
    .a(\u2_Display/n852 ),
    .b(1'b1),
    .c(\u2_Display/add31/c19 ),
    .o({\u2_Display/add31/c20 ,\u2_Display/n874 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u2  (
    .a(\u2_Display/n869 ),
    .b(1'b1),
    .c(\u2_Display/add31/c2 ),
    .o({\u2_Display/add31/c3 ,\u2_Display/n874 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u20  (
    .a(\u2_Display/n851 ),
    .b(1'b1),
    .c(\u2_Display/add31/c20 ),
    .o({\u2_Display/add31/c21 ,\u2_Display/n874 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u21  (
    .a(\u2_Display/n850 ),
    .b(1'b1),
    .c(\u2_Display/add31/c21 ),
    .o({\u2_Display/add31/c22 ,\u2_Display/n874 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u22  (
    .a(\u2_Display/n849 ),
    .b(1'b1),
    .c(\u2_Display/add31/c22 ),
    .o({\u2_Display/add31/c23 ,\u2_Display/n874 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u23  (
    .a(\u2_Display/n848 ),
    .b(1'b1),
    .c(\u2_Display/add31/c23 ),
    .o({\u2_Display/add31/c24 ,\u2_Display/n874 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u24  (
    .a(\u2_Display/n847 ),
    .b(1'b1),
    .c(\u2_Display/add31/c24 ),
    .o({\u2_Display/add31/c25 ,\u2_Display/n874 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u25  (
    .a(\u2_Display/n846 ),
    .b(1'b1),
    .c(\u2_Display/add31/c25 ),
    .o({\u2_Display/add31/c26 ,\u2_Display/n874 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u26  (
    .a(\u2_Display/n845 ),
    .b(1'b1),
    .c(\u2_Display/add31/c26 ),
    .o({\u2_Display/add31/c27 ,\u2_Display/n874 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u27  (
    .a(\u2_Display/n844 ),
    .b(1'b1),
    .c(\u2_Display/add31/c27 ),
    .o({\u2_Display/add31/c28 ,\u2_Display/n874 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u28  (
    .a(\u2_Display/n843 ),
    .b(1'b1),
    .c(\u2_Display/add31/c28 ),
    .o({\u2_Display/add31/c29 ,\u2_Display/n874 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u29  (
    .a(\u2_Display/n842 ),
    .b(1'b1),
    .c(\u2_Display/add31/c29 ),
    .o({\u2_Display/add31/c30 ,\u2_Display/n874 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u3  (
    .a(\u2_Display/n868 ),
    .b(1'b1),
    .c(\u2_Display/add31/c3 ),
    .o({\u2_Display/add31/c4 ,\u2_Display/n874 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u30  (
    .a(\u2_Display/n841 ),
    .b(1'b1),
    .c(\u2_Display/add31/c30 ),
    .o({\u2_Display/add31/c31 ,\u2_Display/n874 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u31  (
    .a(\u2_Display/n840 ),
    .b(1'b1),
    .c(\u2_Display/add31/c31 ),
    .o({open_n1149,\u2_Display/n874 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u4  (
    .a(\u2_Display/n867 ),
    .b(1'b1),
    .c(\u2_Display/add31/c4 ),
    .o({\u2_Display/add31/c5 ,\u2_Display/n874 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u5  (
    .a(\u2_Display/n866 ),
    .b(1'b1),
    .c(\u2_Display/add31/c5 ),
    .o({\u2_Display/add31/c6 ,\u2_Display/n874 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u6  (
    .a(\u2_Display/n865 ),
    .b(1'b1),
    .c(\u2_Display/add31/c6 ),
    .o({\u2_Display/add31/c7 ,\u2_Display/n874 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u7  (
    .a(\u2_Display/n864 ),
    .b(1'b1),
    .c(\u2_Display/add31/c7 ),
    .o({\u2_Display/add31/c8 ,\u2_Display/n874 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u8  (
    .a(\u2_Display/n863 ),
    .b(1'b1),
    .c(\u2_Display/add31/c8 ),
    .o({\u2_Display/add31/c9 ,\u2_Display/n874 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add31/u9  (
    .a(\u2_Display/n862 ),
    .b(1'b1),
    .c(\u2_Display/add31/c9 ),
    .o({\u2_Display/add31/c10 ,\u2_Display/n874 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add31/ucin  (
    .a(1'b1),
    .o({\u2_Display/add31/c0 ,open_n1152}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u0  (
    .a(\u2_Display/n906 ),
    .b(1'b1),
    .c(\u2_Display/add32/c0 ),
    .o({\u2_Display/add32/c1 ,\u2_Display/n909 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u1  (
    .a(\u2_Display/n905 ),
    .b(1'b1),
    .c(\u2_Display/add32/c1 ),
    .o({\u2_Display/add32/c2 ,\u2_Display/n909 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u10  (
    .a(\u2_Display/n896 ),
    .b(1'b1),
    .c(\u2_Display/add32/c10 ),
    .o({\u2_Display/add32/c11 ,\u2_Display/n909 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u11  (
    .a(\u2_Display/n895 ),
    .b(1'b0),
    .c(\u2_Display/add32/c11 ),
    .o({\u2_Display/add32/c12 ,\u2_Display/n909 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u12  (
    .a(\u2_Display/n894 ),
    .b(1'b1),
    .c(\u2_Display/add32/c12 ),
    .o({\u2_Display/add32/c13 ,\u2_Display/n909 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u13  (
    .a(\u2_Display/n893 ),
    .b(1'b0),
    .c(\u2_Display/add32/c13 ),
    .o({\u2_Display/add32/c14 ,\u2_Display/n909 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u14  (
    .a(\u2_Display/n892 ),
    .b(1'b0),
    .c(\u2_Display/add32/c14 ),
    .o({\u2_Display/add32/c15 ,\u2_Display/n909 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u15  (
    .a(\u2_Display/n891 ),
    .b(1'b0),
    .c(\u2_Display/add32/c15 ),
    .o({\u2_Display/add32/c16 ,\u2_Display/n909 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u16  (
    .a(\u2_Display/n890 ),
    .b(1'b0),
    .c(\u2_Display/add32/c16 ),
    .o({\u2_Display/add32/c17 ,\u2_Display/n909 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u17  (
    .a(\u2_Display/n889 ),
    .b(1'b0),
    .c(\u2_Display/add32/c17 ),
    .o({\u2_Display/add32/c18 ,\u2_Display/n909 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u18  (
    .a(\u2_Display/n888 ),
    .b(1'b1),
    .c(\u2_Display/add32/c18 ),
    .o({\u2_Display/add32/c19 ,\u2_Display/n909 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u19  (
    .a(\u2_Display/n887 ),
    .b(1'b1),
    .c(\u2_Display/add32/c19 ),
    .o({\u2_Display/add32/c20 ,\u2_Display/n909 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u2  (
    .a(\u2_Display/n904 ),
    .b(1'b1),
    .c(\u2_Display/add32/c2 ),
    .o({\u2_Display/add32/c3 ,\u2_Display/n909 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u20  (
    .a(\u2_Display/n886 ),
    .b(1'b1),
    .c(\u2_Display/add32/c20 ),
    .o({\u2_Display/add32/c21 ,\u2_Display/n909 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u21  (
    .a(\u2_Display/n885 ),
    .b(1'b1),
    .c(\u2_Display/add32/c21 ),
    .o({\u2_Display/add32/c22 ,\u2_Display/n909 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u22  (
    .a(\u2_Display/n884 ),
    .b(1'b1),
    .c(\u2_Display/add32/c22 ),
    .o({\u2_Display/add32/c23 ,\u2_Display/n909 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u23  (
    .a(\u2_Display/n883 ),
    .b(1'b1),
    .c(\u2_Display/add32/c23 ),
    .o({\u2_Display/add32/c24 ,\u2_Display/n909 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u24  (
    .a(\u2_Display/n882 ),
    .b(1'b1),
    .c(\u2_Display/add32/c24 ),
    .o({\u2_Display/add32/c25 ,\u2_Display/n909 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u25  (
    .a(\u2_Display/n881 ),
    .b(1'b1),
    .c(\u2_Display/add32/c25 ),
    .o({\u2_Display/add32/c26 ,\u2_Display/n909 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u26  (
    .a(\u2_Display/n880 ),
    .b(1'b1),
    .c(\u2_Display/add32/c26 ),
    .o({\u2_Display/add32/c27 ,\u2_Display/n909 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u27  (
    .a(\u2_Display/n879 ),
    .b(1'b1),
    .c(\u2_Display/add32/c27 ),
    .o({\u2_Display/add32/c28 ,\u2_Display/n909 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u28  (
    .a(\u2_Display/n878 ),
    .b(1'b1),
    .c(\u2_Display/add32/c28 ),
    .o({\u2_Display/add32/c29 ,\u2_Display/n909 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u29  (
    .a(\u2_Display/n877 ),
    .b(1'b1),
    .c(\u2_Display/add32/c29 ),
    .o({\u2_Display/add32/c30 ,\u2_Display/n909 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u3  (
    .a(\u2_Display/n903 ),
    .b(1'b1),
    .c(\u2_Display/add32/c3 ),
    .o({\u2_Display/add32/c4 ,\u2_Display/n909 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u30  (
    .a(\u2_Display/n876 ),
    .b(1'b1),
    .c(\u2_Display/add32/c30 ),
    .o({\u2_Display/add32/c31 ,\u2_Display/n909 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u31  (
    .a(\u2_Display/n875 ),
    .b(1'b1),
    .c(\u2_Display/add32/c31 ),
    .o({open_n1153,\u2_Display/n909 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u4  (
    .a(\u2_Display/n902 ),
    .b(1'b1),
    .c(\u2_Display/add32/c4 ),
    .o({\u2_Display/add32/c5 ,\u2_Display/n909 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u5  (
    .a(\u2_Display/n901 ),
    .b(1'b1),
    .c(\u2_Display/add32/c5 ),
    .o({\u2_Display/add32/c6 ,\u2_Display/n909 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u6  (
    .a(\u2_Display/n900 ),
    .b(1'b1),
    .c(\u2_Display/add32/c6 ),
    .o({\u2_Display/add32/c7 ,\u2_Display/n909 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u7  (
    .a(\u2_Display/n899 ),
    .b(1'b1),
    .c(\u2_Display/add32/c7 ),
    .o({\u2_Display/add32/c8 ,\u2_Display/n909 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u8  (
    .a(\u2_Display/n898 ),
    .b(1'b1),
    .c(\u2_Display/add32/c8 ),
    .o({\u2_Display/add32/c9 ,\u2_Display/n909 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add32/u9  (
    .a(\u2_Display/n897 ),
    .b(1'b1),
    .c(\u2_Display/add32/c9 ),
    .o({\u2_Display/add32/c10 ,\u2_Display/n909 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add32/ucin  (
    .a(1'b1),
    .o({\u2_Display/add32/c0 ,open_n1156}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u0  (
    .a(\u2_Display/n941 ),
    .b(1'b1),
    .c(\u2_Display/add33/c0 ),
    .o({\u2_Display/add33/c1 ,\u2_Display/n944 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u1  (
    .a(\u2_Display/n940 ),
    .b(1'b1),
    .c(\u2_Display/add33/c1 ),
    .o({\u2_Display/add33/c2 ,\u2_Display/n944 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u10  (
    .a(\u2_Display/n931 ),
    .b(1'b0),
    .c(\u2_Display/add33/c10 ),
    .o({\u2_Display/add33/c11 ,\u2_Display/n944 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u11  (
    .a(\u2_Display/n930 ),
    .b(1'b1),
    .c(\u2_Display/add33/c11 ),
    .o({\u2_Display/add33/c12 ,\u2_Display/n944 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u12  (
    .a(\u2_Display/n929 ),
    .b(1'b0),
    .c(\u2_Display/add33/c12 ),
    .o({\u2_Display/add33/c13 ,\u2_Display/n944 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u13  (
    .a(\u2_Display/n928 ),
    .b(1'b0),
    .c(\u2_Display/add33/c13 ),
    .o({\u2_Display/add33/c14 ,\u2_Display/n944 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u14  (
    .a(\u2_Display/n927 ),
    .b(1'b0),
    .c(\u2_Display/add33/c14 ),
    .o({\u2_Display/add33/c15 ,\u2_Display/n944 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u15  (
    .a(\u2_Display/n926 ),
    .b(1'b0),
    .c(\u2_Display/add33/c15 ),
    .o({\u2_Display/add33/c16 ,\u2_Display/n944 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u16  (
    .a(\u2_Display/n925 ),
    .b(1'b0),
    .c(\u2_Display/add33/c16 ),
    .o({\u2_Display/add33/c17 ,\u2_Display/n944 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u17  (
    .a(\u2_Display/n924 ),
    .b(1'b1),
    .c(\u2_Display/add33/c17 ),
    .o({\u2_Display/add33/c18 ,\u2_Display/n944 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u18  (
    .a(\u2_Display/n923 ),
    .b(1'b1),
    .c(\u2_Display/add33/c18 ),
    .o({\u2_Display/add33/c19 ,\u2_Display/n944 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u19  (
    .a(\u2_Display/n922 ),
    .b(1'b1),
    .c(\u2_Display/add33/c19 ),
    .o({\u2_Display/add33/c20 ,\u2_Display/n944 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u2  (
    .a(\u2_Display/n939 ),
    .b(1'b1),
    .c(\u2_Display/add33/c2 ),
    .o({\u2_Display/add33/c3 ,\u2_Display/n944 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u20  (
    .a(\u2_Display/n921 ),
    .b(1'b1),
    .c(\u2_Display/add33/c20 ),
    .o({\u2_Display/add33/c21 ,\u2_Display/n944 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u21  (
    .a(\u2_Display/n920 ),
    .b(1'b1),
    .c(\u2_Display/add33/c21 ),
    .o({\u2_Display/add33/c22 ,\u2_Display/n944 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u22  (
    .a(\u2_Display/n919 ),
    .b(1'b1),
    .c(\u2_Display/add33/c22 ),
    .o({\u2_Display/add33/c23 ,\u2_Display/n944 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u23  (
    .a(\u2_Display/n918 ),
    .b(1'b1),
    .c(\u2_Display/add33/c23 ),
    .o({\u2_Display/add33/c24 ,\u2_Display/n944 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u24  (
    .a(\u2_Display/n917 ),
    .b(1'b1),
    .c(\u2_Display/add33/c24 ),
    .o({\u2_Display/add33/c25 ,\u2_Display/n944 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u25  (
    .a(\u2_Display/n916 ),
    .b(1'b1),
    .c(\u2_Display/add33/c25 ),
    .o({\u2_Display/add33/c26 ,\u2_Display/n944 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u26  (
    .a(\u2_Display/n915 ),
    .b(1'b1),
    .c(\u2_Display/add33/c26 ),
    .o({\u2_Display/add33/c27 ,\u2_Display/n944 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u27  (
    .a(\u2_Display/n914 ),
    .b(1'b1),
    .c(\u2_Display/add33/c27 ),
    .o({\u2_Display/add33/c28 ,\u2_Display/n944 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u28  (
    .a(\u2_Display/n913 ),
    .b(1'b1),
    .c(\u2_Display/add33/c28 ),
    .o({\u2_Display/add33/c29 ,\u2_Display/n944 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u29  (
    .a(\u2_Display/n912 ),
    .b(1'b1),
    .c(\u2_Display/add33/c29 ),
    .o({\u2_Display/add33/c30 ,\u2_Display/n944 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u3  (
    .a(\u2_Display/n938 ),
    .b(1'b1),
    .c(\u2_Display/add33/c3 ),
    .o({\u2_Display/add33/c4 ,\u2_Display/n944 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u30  (
    .a(\u2_Display/n911 ),
    .b(1'b1),
    .c(\u2_Display/add33/c30 ),
    .o({\u2_Display/add33/c31 ,\u2_Display/n944 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u31  (
    .a(\u2_Display/n910 ),
    .b(1'b1),
    .c(\u2_Display/add33/c31 ),
    .o({open_n1157,\u2_Display/n944 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u4  (
    .a(\u2_Display/n937 ),
    .b(1'b1),
    .c(\u2_Display/add33/c4 ),
    .o({\u2_Display/add33/c5 ,\u2_Display/n944 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u5  (
    .a(\u2_Display/n936 ),
    .b(1'b1),
    .c(\u2_Display/add33/c5 ),
    .o({\u2_Display/add33/c6 ,\u2_Display/n944 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u6  (
    .a(\u2_Display/n935 ),
    .b(1'b1),
    .c(\u2_Display/add33/c6 ),
    .o({\u2_Display/add33/c7 ,\u2_Display/n944 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u7  (
    .a(\u2_Display/n934 ),
    .b(1'b1),
    .c(\u2_Display/add33/c7 ),
    .o({\u2_Display/add33/c8 ,\u2_Display/n944 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u8  (
    .a(\u2_Display/n933 ),
    .b(1'b1),
    .c(\u2_Display/add33/c8 ),
    .o({\u2_Display/add33/c9 ,\u2_Display/n944 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add33/u9  (
    .a(\u2_Display/n932 ),
    .b(1'b1),
    .c(\u2_Display/add33/c9 ),
    .o({\u2_Display/add33/c10 ,\u2_Display/n944 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add33/ucin  (
    .a(1'b1),
    .o({\u2_Display/add33/c0 ,open_n1160}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u0  (
    .a(\u2_Display/n976 ),
    .b(1'b1),
    .c(\u2_Display/add34/c0 ),
    .o({\u2_Display/add34/c1 ,\u2_Display/n979 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u1  (
    .a(\u2_Display/n975 ),
    .b(1'b1),
    .c(\u2_Display/add34/c1 ),
    .o({\u2_Display/add34/c2 ,\u2_Display/n979 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u10  (
    .a(\u2_Display/n966 ),
    .b(1'b1),
    .c(\u2_Display/add34/c10 ),
    .o({\u2_Display/add34/c11 ,\u2_Display/n979 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u11  (
    .a(\u2_Display/n965 ),
    .b(1'b0),
    .c(\u2_Display/add34/c11 ),
    .o({\u2_Display/add34/c12 ,\u2_Display/n979 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u12  (
    .a(\u2_Display/n964 ),
    .b(1'b0),
    .c(\u2_Display/add34/c12 ),
    .o({\u2_Display/add34/c13 ,\u2_Display/n979 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u13  (
    .a(\u2_Display/n963 ),
    .b(1'b0),
    .c(\u2_Display/add34/c13 ),
    .o({\u2_Display/add34/c14 ,\u2_Display/n979 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u14  (
    .a(\u2_Display/n962 ),
    .b(1'b0),
    .c(\u2_Display/add34/c14 ),
    .o({\u2_Display/add34/c15 ,\u2_Display/n979 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u15  (
    .a(\u2_Display/n961 ),
    .b(1'b0),
    .c(\u2_Display/add34/c15 ),
    .o({\u2_Display/add34/c16 ,\u2_Display/n979 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u16  (
    .a(\u2_Display/n960 ),
    .b(1'b1),
    .c(\u2_Display/add34/c16 ),
    .o({\u2_Display/add34/c17 ,\u2_Display/n979 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u17  (
    .a(\u2_Display/n959 ),
    .b(1'b1),
    .c(\u2_Display/add34/c17 ),
    .o({\u2_Display/add34/c18 ,\u2_Display/n979 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u18  (
    .a(\u2_Display/n958 ),
    .b(1'b1),
    .c(\u2_Display/add34/c18 ),
    .o({\u2_Display/add34/c19 ,\u2_Display/n979 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u19  (
    .a(\u2_Display/n957 ),
    .b(1'b1),
    .c(\u2_Display/add34/c19 ),
    .o({\u2_Display/add34/c20 ,\u2_Display/n979 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u2  (
    .a(\u2_Display/n974 ),
    .b(1'b1),
    .c(\u2_Display/add34/c2 ),
    .o({\u2_Display/add34/c3 ,\u2_Display/n979 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u20  (
    .a(\u2_Display/n956 ),
    .b(1'b1),
    .c(\u2_Display/add34/c20 ),
    .o({\u2_Display/add34/c21 ,\u2_Display/n979 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u21  (
    .a(\u2_Display/n955 ),
    .b(1'b1),
    .c(\u2_Display/add34/c21 ),
    .o({\u2_Display/add34/c22 ,\u2_Display/n979 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u22  (
    .a(\u2_Display/n954 ),
    .b(1'b1),
    .c(\u2_Display/add34/c22 ),
    .o({\u2_Display/add34/c23 ,\u2_Display/n979 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u23  (
    .a(\u2_Display/n953 ),
    .b(1'b1),
    .c(\u2_Display/add34/c23 ),
    .o({\u2_Display/add34/c24 ,\u2_Display/n979 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u24  (
    .a(\u2_Display/n952 ),
    .b(1'b1),
    .c(\u2_Display/add34/c24 ),
    .o({\u2_Display/add34/c25 ,\u2_Display/n979 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u25  (
    .a(\u2_Display/n951 ),
    .b(1'b1),
    .c(\u2_Display/add34/c25 ),
    .o({\u2_Display/add34/c26 ,\u2_Display/n979 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u26  (
    .a(\u2_Display/n950 ),
    .b(1'b1),
    .c(\u2_Display/add34/c26 ),
    .o({\u2_Display/add34/c27 ,\u2_Display/n979 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u27  (
    .a(\u2_Display/n949 ),
    .b(1'b1),
    .c(\u2_Display/add34/c27 ),
    .o({\u2_Display/add34/c28 ,\u2_Display/n979 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u28  (
    .a(\u2_Display/n948 ),
    .b(1'b1),
    .c(\u2_Display/add34/c28 ),
    .o({\u2_Display/add34/c29 ,\u2_Display/n979 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u29  (
    .a(\u2_Display/n947 ),
    .b(1'b1),
    .c(\u2_Display/add34/c29 ),
    .o({\u2_Display/add34/c30 ,\u2_Display/n979 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u3  (
    .a(\u2_Display/n973 ),
    .b(1'b1),
    .c(\u2_Display/add34/c3 ),
    .o({\u2_Display/add34/c4 ,\u2_Display/n979 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u30  (
    .a(\u2_Display/n946 ),
    .b(1'b1),
    .c(\u2_Display/add34/c30 ),
    .o({\u2_Display/add34/c31 ,\u2_Display/n979 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u31  (
    .a(\u2_Display/n945 ),
    .b(1'b1),
    .c(\u2_Display/add34/c31 ),
    .o({open_n1161,\u2_Display/n979 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u4  (
    .a(\u2_Display/n972 ),
    .b(1'b1),
    .c(\u2_Display/add34/c4 ),
    .o({\u2_Display/add34/c5 ,\u2_Display/n979 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u5  (
    .a(\u2_Display/n971 ),
    .b(1'b1),
    .c(\u2_Display/add34/c5 ),
    .o({\u2_Display/add34/c6 ,\u2_Display/n979 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u6  (
    .a(\u2_Display/n970 ),
    .b(1'b1),
    .c(\u2_Display/add34/c6 ),
    .o({\u2_Display/add34/c7 ,\u2_Display/n979 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u7  (
    .a(\u2_Display/n969 ),
    .b(1'b1),
    .c(\u2_Display/add34/c7 ),
    .o({\u2_Display/add34/c8 ,\u2_Display/n979 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u8  (
    .a(\u2_Display/n968 ),
    .b(1'b1),
    .c(\u2_Display/add34/c8 ),
    .o({\u2_Display/add34/c9 ,\u2_Display/n979 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add34/u9  (
    .a(\u2_Display/n967 ),
    .b(1'b0),
    .c(\u2_Display/add34/c9 ),
    .o({\u2_Display/add34/c10 ,\u2_Display/n979 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add34/ucin  (
    .a(1'b1),
    .o({\u2_Display/add34/c0 ,open_n1164}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u0  (
    .a(\u2_Display/n1011 ),
    .b(1'b1),
    .c(\u2_Display/add35/c0 ),
    .o({\u2_Display/add35/c1 ,\u2_Display/n1014 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u1  (
    .a(\u2_Display/n1010 ),
    .b(1'b1),
    .c(\u2_Display/add35/c1 ),
    .o({\u2_Display/add35/c2 ,\u2_Display/n1014 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u10  (
    .a(\u2_Display/n1001 ),
    .b(1'b0),
    .c(\u2_Display/add35/c10 ),
    .o({\u2_Display/add35/c11 ,\u2_Display/n1014 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u11  (
    .a(\u2_Display/n1000 ),
    .b(1'b0),
    .c(\u2_Display/add35/c11 ),
    .o({\u2_Display/add35/c12 ,\u2_Display/n1014 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u12  (
    .a(\u2_Display/n999 ),
    .b(1'b0),
    .c(\u2_Display/add35/c12 ),
    .o({\u2_Display/add35/c13 ,\u2_Display/n1014 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u13  (
    .a(\u2_Display/n998 ),
    .b(1'b0),
    .c(\u2_Display/add35/c13 ),
    .o({\u2_Display/add35/c14 ,\u2_Display/n1014 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u14  (
    .a(\u2_Display/n997 ),
    .b(1'b0),
    .c(\u2_Display/add35/c14 ),
    .o({\u2_Display/add35/c15 ,\u2_Display/n1014 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u15  (
    .a(\u2_Display/n996 ),
    .b(1'b1),
    .c(\u2_Display/add35/c15 ),
    .o({\u2_Display/add35/c16 ,\u2_Display/n1014 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u16  (
    .a(\u2_Display/n995 ),
    .b(1'b1),
    .c(\u2_Display/add35/c16 ),
    .o({\u2_Display/add35/c17 ,\u2_Display/n1014 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u17  (
    .a(\u2_Display/n994 ),
    .b(1'b1),
    .c(\u2_Display/add35/c17 ),
    .o({\u2_Display/add35/c18 ,\u2_Display/n1014 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u18  (
    .a(\u2_Display/n993 ),
    .b(1'b1),
    .c(\u2_Display/add35/c18 ),
    .o({\u2_Display/add35/c19 ,\u2_Display/n1014 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u19  (
    .a(\u2_Display/n992 ),
    .b(1'b1),
    .c(\u2_Display/add35/c19 ),
    .o({\u2_Display/add35/c20 ,\u2_Display/n1014 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u2  (
    .a(\u2_Display/n1009 ),
    .b(1'b1),
    .c(\u2_Display/add35/c2 ),
    .o({\u2_Display/add35/c3 ,\u2_Display/n1014 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u20  (
    .a(\u2_Display/n991 ),
    .b(1'b1),
    .c(\u2_Display/add35/c20 ),
    .o({\u2_Display/add35/c21 ,\u2_Display/n1014 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u21  (
    .a(\u2_Display/n990 ),
    .b(1'b1),
    .c(\u2_Display/add35/c21 ),
    .o({\u2_Display/add35/c22 ,\u2_Display/n1014 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u22  (
    .a(\u2_Display/n989 ),
    .b(1'b1),
    .c(\u2_Display/add35/c22 ),
    .o({\u2_Display/add35/c23 ,\u2_Display/n1014 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u23  (
    .a(\u2_Display/n988 ),
    .b(1'b1),
    .c(\u2_Display/add35/c23 ),
    .o({\u2_Display/add35/c24 ,\u2_Display/n1014 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u24  (
    .a(\u2_Display/n987 ),
    .b(1'b1),
    .c(\u2_Display/add35/c24 ),
    .o({\u2_Display/add35/c25 ,\u2_Display/n1014 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u25  (
    .a(\u2_Display/n986 ),
    .b(1'b1),
    .c(\u2_Display/add35/c25 ),
    .o({\u2_Display/add35/c26 ,\u2_Display/n1014 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u26  (
    .a(\u2_Display/n985 ),
    .b(1'b1),
    .c(\u2_Display/add35/c26 ),
    .o({\u2_Display/add35/c27 ,\u2_Display/n1014 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u27  (
    .a(\u2_Display/n984 ),
    .b(1'b1),
    .c(\u2_Display/add35/c27 ),
    .o({\u2_Display/add35/c28 ,\u2_Display/n1014 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u28  (
    .a(\u2_Display/n983 ),
    .b(1'b1),
    .c(\u2_Display/add35/c28 ),
    .o({\u2_Display/add35/c29 ,\u2_Display/n1014 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u29  (
    .a(\u2_Display/n982 ),
    .b(1'b1),
    .c(\u2_Display/add35/c29 ),
    .o({\u2_Display/add35/c30 ,\u2_Display/n1014 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u3  (
    .a(\u2_Display/n1008 ),
    .b(1'b1),
    .c(\u2_Display/add35/c3 ),
    .o({\u2_Display/add35/c4 ,\u2_Display/n1014 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u30  (
    .a(\u2_Display/n981 ),
    .b(1'b1),
    .c(\u2_Display/add35/c30 ),
    .o({\u2_Display/add35/c31 ,\u2_Display/n1014 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u31  (
    .a(\u2_Display/n980 ),
    .b(1'b1),
    .c(\u2_Display/add35/c31 ),
    .o({open_n1165,\u2_Display/n1014 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u4  (
    .a(\u2_Display/n1007 ),
    .b(1'b1),
    .c(\u2_Display/add35/c4 ),
    .o({\u2_Display/add35/c5 ,\u2_Display/n1014 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u5  (
    .a(\u2_Display/n1006 ),
    .b(1'b1),
    .c(\u2_Display/add35/c5 ),
    .o({\u2_Display/add35/c6 ,\u2_Display/n1014 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u6  (
    .a(\u2_Display/n1005 ),
    .b(1'b1),
    .c(\u2_Display/add35/c6 ),
    .o({\u2_Display/add35/c7 ,\u2_Display/n1014 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u7  (
    .a(\u2_Display/n1004 ),
    .b(1'b1),
    .c(\u2_Display/add35/c7 ),
    .o({\u2_Display/add35/c8 ,\u2_Display/n1014 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u8  (
    .a(\u2_Display/n1003 ),
    .b(1'b0),
    .c(\u2_Display/add35/c8 ),
    .o({\u2_Display/add35/c9 ,\u2_Display/n1014 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add35/u9  (
    .a(\u2_Display/n1002 ),
    .b(1'b1),
    .c(\u2_Display/add35/c9 ),
    .o({\u2_Display/add35/c10 ,\u2_Display/n1014 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add35/ucin  (
    .a(1'b1),
    .o({\u2_Display/add35/c0 ,open_n1168}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u0  (
    .a(\u2_Display/n1046 ),
    .b(1'b1),
    .c(\u2_Display/add36/c0 ),
    .o({\u2_Display/add36/c1 ,\u2_Display/n1049 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u1  (
    .a(\u2_Display/n1045 ),
    .b(1'b1),
    .c(\u2_Display/add36/c1 ),
    .o({\u2_Display/add36/c2 ,\u2_Display/n1049 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u10  (
    .a(\u2_Display/n1036 ),
    .b(1'b0),
    .c(\u2_Display/add36/c10 ),
    .o({\u2_Display/add36/c11 ,\u2_Display/n1049 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u11  (
    .a(\u2_Display/n1035 ),
    .b(1'b0),
    .c(\u2_Display/add36/c11 ),
    .o({\u2_Display/add36/c12 ,\u2_Display/n1049 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u12  (
    .a(\u2_Display/n1034 ),
    .b(1'b0),
    .c(\u2_Display/add36/c12 ),
    .o({\u2_Display/add36/c13 ,\u2_Display/n1049 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u13  (
    .a(\u2_Display/n1033 ),
    .b(1'b0),
    .c(\u2_Display/add36/c13 ),
    .o({\u2_Display/add36/c14 ,\u2_Display/n1049 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u14  (
    .a(\u2_Display/n1032 ),
    .b(1'b1),
    .c(\u2_Display/add36/c14 ),
    .o({\u2_Display/add36/c15 ,\u2_Display/n1049 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u15  (
    .a(\u2_Display/n1031 ),
    .b(1'b1),
    .c(\u2_Display/add36/c15 ),
    .o({\u2_Display/add36/c16 ,\u2_Display/n1049 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u16  (
    .a(\u2_Display/n1030 ),
    .b(1'b1),
    .c(\u2_Display/add36/c16 ),
    .o({\u2_Display/add36/c17 ,\u2_Display/n1049 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u17  (
    .a(\u2_Display/n1029 ),
    .b(1'b1),
    .c(\u2_Display/add36/c17 ),
    .o({\u2_Display/add36/c18 ,\u2_Display/n1049 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u18  (
    .a(\u2_Display/n1028 ),
    .b(1'b1),
    .c(\u2_Display/add36/c18 ),
    .o({\u2_Display/add36/c19 ,\u2_Display/n1049 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u19  (
    .a(\u2_Display/n1027 ),
    .b(1'b1),
    .c(\u2_Display/add36/c19 ),
    .o({\u2_Display/add36/c20 ,\u2_Display/n1049 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u2  (
    .a(\u2_Display/n1044 ),
    .b(1'b1),
    .c(\u2_Display/add36/c2 ),
    .o({\u2_Display/add36/c3 ,\u2_Display/n1049 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u20  (
    .a(\u2_Display/n1026 ),
    .b(1'b1),
    .c(\u2_Display/add36/c20 ),
    .o({\u2_Display/add36/c21 ,\u2_Display/n1049 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u21  (
    .a(\u2_Display/n1025 ),
    .b(1'b1),
    .c(\u2_Display/add36/c21 ),
    .o({\u2_Display/add36/c22 ,\u2_Display/n1049 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u22  (
    .a(\u2_Display/n1024 ),
    .b(1'b1),
    .c(\u2_Display/add36/c22 ),
    .o({\u2_Display/add36/c23 ,\u2_Display/n1049 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u23  (
    .a(\u2_Display/n1023 ),
    .b(1'b1),
    .c(\u2_Display/add36/c23 ),
    .o({\u2_Display/add36/c24 ,\u2_Display/n1049 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u24  (
    .a(\u2_Display/n1022 ),
    .b(1'b1),
    .c(\u2_Display/add36/c24 ),
    .o({\u2_Display/add36/c25 ,\u2_Display/n1049 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u25  (
    .a(\u2_Display/n1021 ),
    .b(1'b1),
    .c(\u2_Display/add36/c25 ),
    .o({\u2_Display/add36/c26 ,\u2_Display/n1049 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u26  (
    .a(\u2_Display/n1020 ),
    .b(1'b1),
    .c(\u2_Display/add36/c26 ),
    .o({\u2_Display/add36/c27 ,\u2_Display/n1049 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u27  (
    .a(\u2_Display/n1019 ),
    .b(1'b1),
    .c(\u2_Display/add36/c27 ),
    .o({\u2_Display/add36/c28 ,\u2_Display/n1049 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u28  (
    .a(\u2_Display/n1018 ),
    .b(1'b1),
    .c(\u2_Display/add36/c28 ),
    .o({\u2_Display/add36/c29 ,\u2_Display/n1049 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u29  (
    .a(\u2_Display/n1017 ),
    .b(1'b1),
    .c(\u2_Display/add36/c29 ),
    .o({\u2_Display/add36/c30 ,\u2_Display/n1049 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u3  (
    .a(\u2_Display/n1043 ),
    .b(1'b1),
    .c(\u2_Display/add36/c3 ),
    .o({\u2_Display/add36/c4 ,\u2_Display/n1049 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u30  (
    .a(\u2_Display/n1016 ),
    .b(1'b1),
    .c(\u2_Display/add36/c30 ),
    .o({\u2_Display/add36/c31 ,\u2_Display/n1049 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u31  (
    .a(\u2_Display/n1015 ),
    .b(1'b1),
    .c(\u2_Display/add36/c31 ),
    .o({open_n1169,\u2_Display/n1049 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u4  (
    .a(\u2_Display/n1042 ),
    .b(1'b1),
    .c(\u2_Display/add36/c4 ),
    .o({\u2_Display/add36/c5 ,\u2_Display/n1049 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u5  (
    .a(\u2_Display/n1041 ),
    .b(1'b1),
    .c(\u2_Display/add36/c5 ),
    .o({\u2_Display/add36/c6 ,\u2_Display/n1049 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u6  (
    .a(\u2_Display/n1040 ),
    .b(1'b1),
    .c(\u2_Display/add36/c6 ),
    .o({\u2_Display/add36/c7 ,\u2_Display/n1049 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u7  (
    .a(\u2_Display/n1039 ),
    .b(1'b0),
    .c(\u2_Display/add36/c7 ),
    .o({\u2_Display/add36/c8 ,\u2_Display/n1049 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u8  (
    .a(\u2_Display/n1038 ),
    .b(1'b1),
    .c(\u2_Display/add36/c8 ),
    .o({\u2_Display/add36/c9 ,\u2_Display/n1049 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add36/u9  (
    .a(\u2_Display/n1037 ),
    .b(1'b0),
    .c(\u2_Display/add36/c9 ),
    .o({\u2_Display/add36/c10 ,\u2_Display/n1049 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add36/ucin  (
    .a(1'b1),
    .o({\u2_Display/add36/c0 ,open_n1172}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u0  (
    .a(\u2_Display/n1081 ),
    .b(1'b1),
    .c(\u2_Display/add37/c0 ),
    .o({\u2_Display/add37/c1 ,\u2_Display/n1084 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u1  (
    .a(\u2_Display/n1080 ),
    .b(1'b1),
    .c(\u2_Display/add37/c1 ),
    .o({\u2_Display/add37/c2 ,\u2_Display/n1084 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u10  (
    .a(\u2_Display/n1071 ),
    .b(1'b0),
    .c(\u2_Display/add37/c10 ),
    .o({\u2_Display/add37/c11 ,\u2_Display/n1084 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u11  (
    .a(\u2_Display/n1070 ),
    .b(1'b0),
    .c(\u2_Display/add37/c11 ),
    .o({\u2_Display/add37/c12 ,\u2_Display/n1084 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u12  (
    .a(\u2_Display/n1069 ),
    .b(1'b0),
    .c(\u2_Display/add37/c12 ),
    .o({\u2_Display/add37/c13 ,\u2_Display/n1084 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u13  (
    .a(\u2_Display/n1068 ),
    .b(1'b1),
    .c(\u2_Display/add37/c13 ),
    .o({\u2_Display/add37/c14 ,\u2_Display/n1084 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u14  (
    .a(\u2_Display/n1067 ),
    .b(1'b1),
    .c(\u2_Display/add37/c14 ),
    .o({\u2_Display/add37/c15 ,\u2_Display/n1084 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u15  (
    .a(\u2_Display/n1066 ),
    .b(1'b1),
    .c(\u2_Display/add37/c15 ),
    .o({\u2_Display/add37/c16 ,\u2_Display/n1084 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u16  (
    .a(\u2_Display/n1065 ),
    .b(1'b1),
    .c(\u2_Display/add37/c16 ),
    .o({\u2_Display/add37/c17 ,\u2_Display/n1084 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u17  (
    .a(\u2_Display/n1064 ),
    .b(1'b1),
    .c(\u2_Display/add37/c17 ),
    .o({\u2_Display/add37/c18 ,\u2_Display/n1084 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u18  (
    .a(\u2_Display/n1063 ),
    .b(1'b1),
    .c(\u2_Display/add37/c18 ),
    .o({\u2_Display/add37/c19 ,\u2_Display/n1084 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u19  (
    .a(\u2_Display/n1062 ),
    .b(1'b1),
    .c(\u2_Display/add37/c19 ),
    .o({\u2_Display/add37/c20 ,\u2_Display/n1084 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u2  (
    .a(\u2_Display/n1079 ),
    .b(1'b1),
    .c(\u2_Display/add37/c2 ),
    .o({\u2_Display/add37/c3 ,\u2_Display/n1084 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u20  (
    .a(\u2_Display/n1061 ),
    .b(1'b1),
    .c(\u2_Display/add37/c20 ),
    .o({\u2_Display/add37/c21 ,\u2_Display/n1084 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u21  (
    .a(\u2_Display/n1060 ),
    .b(1'b1),
    .c(\u2_Display/add37/c21 ),
    .o({\u2_Display/add37/c22 ,\u2_Display/n1084 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u22  (
    .a(\u2_Display/n1059 ),
    .b(1'b1),
    .c(\u2_Display/add37/c22 ),
    .o({\u2_Display/add37/c23 ,\u2_Display/n1084 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u23  (
    .a(\u2_Display/n1058 ),
    .b(1'b1),
    .c(\u2_Display/add37/c23 ),
    .o({\u2_Display/add37/c24 ,\u2_Display/n1084 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u24  (
    .a(\u2_Display/n1057 ),
    .b(1'b1),
    .c(\u2_Display/add37/c24 ),
    .o({\u2_Display/add37/c25 ,\u2_Display/n1084 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u25  (
    .a(\u2_Display/n1056 ),
    .b(1'b1),
    .c(\u2_Display/add37/c25 ),
    .o({\u2_Display/add37/c26 ,\u2_Display/n1084 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u26  (
    .a(\u2_Display/n1055 ),
    .b(1'b1),
    .c(\u2_Display/add37/c26 ),
    .o({\u2_Display/add37/c27 ,\u2_Display/n1084 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u27  (
    .a(\u2_Display/n1054 ),
    .b(1'b1),
    .c(\u2_Display/add37/c27 ),
    .o({\u2_Display/add37/c28 ,\u2_Display/n1084 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u28  (
    .a(\u2_Display/n1053 ),
    .b(1'b1),
    .c(\u2_Display/add37/c28 ),
    .o({\u2_Display/add37/c29 ,\u2_Display/n1084 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u29  (
    .a(\u2_Display/n1052 ),
    .b(1'b1),
    .c(\u2_Display/add37/c29 ),
    .o({\u2_Display/add37/c30 ,\u2_Display/n1084 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u3  (
    .a(\u2_Display/n1078 ),
    .b(1'b1),
    .c(\u2_Display/add37/c3 ),
    .o({\u2_Display/add37/c4 ,\u2_Display/n1084 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u30  (
    .a(\u2_Display/n1051 ),
    .b(1'b1),
    .c(\u2_Display/add37/c30 ),
    .o({\u2_Display/add37/c31 ,\u2_Display/n1084 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u31  (
    .a(\u2_Display/n1050 ),
    .b(1'b1),
    .c(\u2_Display/add37/c31 ),
    .o({open_n1173,\u2_Display/n1084 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u4  (
    .a(\u2_Display/n1077 ),
    .b(1'b1),
    .c(\u2_Display/add37/c4 ),
    .o({\u2_Display/add37/c5 ,\u2_Display/n1084 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u5  (
    .a(\u2_Display/n1076 ),
    .b(1'b1),
    .c(\u2_Display/add37/c5 ),
    .o({\u2_Display/add37/c6 ,\u2_Display/n1084 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u6  (
    .a(\u2_Display/n1075 ),
    .b(1'b0),
    .c(\u2_Display/add37/c6 ),
    .o({\u2_Display/add37/c7 ,\u2_Display/n1084 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u7  (
    .a(\u2_Display/n1074 ),
    .b(1'b1),
    .c(\u2_Display/add37/c7 ),
    .o({\u2_Display/add37/c8 ,\u2_Display/n1084 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u8  (
    .a(\u2_Display/n1073 ),
    .b(1'b0),
    .c(\u2_Display/add37/c8 ),
    .o({\u2_Display/add37/c9 ,\u2_Display/n1084 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add37/u9  (
    .a(\u2_Display/n1072 ),
    .b(1'b0),
    .c(\u2_Display/add37/c9 ),
    .o({\u2_Display/add37/c10 ,\u2_Display/n1084 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add37/ucin  (
    .a(1'b1),
    .o({\u2_Display/add37/c0 ,open_n1176}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u0  (
    .a(\u2_Display/n1116 ),
    .b(1'b1),
    .c(\u2_Display/add38/c0 ),
    .o({\u2_Display/add38/c1 ,\u2_Display/n1119 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u1  (
    .a(\u2_Display/n1115 ),
    .b(1'b1),
    .c(\u2_Display/add38/c1 ),
    .o({\u2_Display/add38/c2 ,\u2_Display/n1119 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u10  (
    .a(\u2_Display/n1106 ),
    .b(1'b0),
    .c(\u2_Display/add38/c10 ),
    .o({\u2_Display/add38/c11 ,\u2_Display/n1119 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u11  (
    .a(\u2_Display/n1105 ),
    .b(1'b0),
    .c(\u2_Display/add38/c11 ),
    .o({\u2_Display/add38/c12 ,\u2_Display/n1119 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u12  (
    .a(\u2_Display/n1104 ),
    .b(1'b1),
    .c(\u2_Display/add38/c12 ),
    .o({\u2_Display/add38/c13 ,\u2_Display/n1119 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u13  (
    .a(\u2_Display/n1103 ),
    .b(1'b1),
    .c(\u2_Display/add38/c13 ),
    .o({\u2_Display/add38/c14 ,\u2_Display/n1119 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u14  (
    .a(\u2_Display/n1102 ),
    .b(1'b1),
    .c(\u2_Display/add38/c14 ),
    .o({\u2_Display/add38/c15 ,\u2_Display/n1119 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u15  (
    .a(\u2_Display/n1101 ),
    .b(1'b1),
    .c(\u2_Display/add38/c15 ),
    .o({\u2_Display/add38/c16 ,\u2_Display/n1119 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u16  (
    .a(\u2_Display/n1100 ),
    .b(1'b1),
    .c(\u2_Display/add38/c16 ),
    .o({\u2_Display/add38/c17 ,\u2_Display/n1119 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u17  (
    .a(\u2_Display/n1099 ),
    .b(1'b1),
    .c(\u2_Display/add38/c17 ),
    .o({\u2_Display/add38/c18 ,\u2_Display/n1119 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u18  (
    .a(\u2_Display/n1098 ),
    .b(1'b1),
    .c(\u2_Display/add38/c18 ),
    .o({\u2_Display/add38/c19 ,\u2_Display/n1119 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u19  (
    .a(\u2_Display/n1097 ),
    .b(1'b1),
    .c(\u2_Display/add38/c19 ),
    .o({\u2_Display/add38/c20 ,\u2_Display/n1119 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u2  (
    .a(\u2_Display/n1114 ),
    .b(1'b1),
    .c(\u2_Display/add38/c2 ),
    .o({\u2_Display/add38/c3 ,\u2_Display/n1119 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u20  (
    .a(\u2_Display/n1096 ),
    .b(1'b1),
    .c(\u2_Display/add38/c20 ),
    .o({\u2_Display/add38/c21 ,\u2_Display/n1119 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u21  (
    .a(\u2_Display/n1095 ),
    .b(1'b1),
    .c(\u2_Display/add38/c21 ),
    .o({\u2_Display/add38/c22 ,\u2_Display/n1119 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u22  (
    .a(\u2_Display/n1094 ),
    .b(1'b1),
    .c(\u2_Display/add38/c22 ),
    .o({\u2_Display/add38/c23 ,\u2_Display/n1119 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u23  (
    .a(\u2_Display/n1093 ),
    .b(1'b1),
    .c(\u2_Display/add38/c23 ),
    .o({\u2_Display/add38/c24 ,\u2_Display/n1119 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u24  (
    .a(\u2_Display/n1092 ),
    .b(1'b1),
    .c(\u2_Display/add38/c24 ),
    .o({\u2_Display/add38/c25 ,\u2_Display/n1119 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u25  (
    .a(\u2_Display/n1091 ),
    .b(1'b1),
    .c(\u2_Display/add38/c25 ),
    .o({\u2_Display/add38/c26 ,\u2_Display/n1119 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u26  (
    .a(\u2_Display/n1090 ),
    .b(1'b1),
    .c(\u2_Display/add38/c26 ),
    .o({\u2_Display/add38/c27 ,\u2_Display/n1119 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u27  (
    .a(\u2_Display/n1089 ),
    .b(1'b1),
    .c(\u2_Display/add38/c27 ),
    .o({\u2_Display/add38/c28 ,\u2_Display/n1119 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u28  (
    .a(\u2_Display/n1088 ),
    .b(1'b1),
    .c(\u2_Display/add38/c28 ),
    .o({\u2_Display/add38/c29 ,\u2_Display/n1119 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u29  (
    .a(\u2_Display/n1087 ),
    .b(1'b1),
    .c(\u2_Display/add38/c29 ),
    .o({\u2_Display/add38/c30 ,\u2_Display/n1119 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u3  (
    .a(\u2_Display/n1113 ),
    .b(1'b1),
    .c(\u2_Display/add38/c3 ),
    .o({\u2_Display/add38/c4 ,\u2_Display/n1119 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u30  (
    .a(\u2_Display/n1086 ),
    .b(1'b1),
    .c(\u2_Display/add38/c30 ),
    .o({\u2_Display/add38/c31 ,\u2_Display/n1119 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u31  (
    .a(\u2_Display/n1085 ),
    .b(1'b1),
    .c(\u2_Display/add38/c31 ),
    .o({open_n1177,\u2_Display/n1119 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u4  (
    .a(\u2_Display/n1112 ),
    .b(1'b1),
    .c(\u2_Display/add38/c4 ),
    .o({\u2_Display/add38/c5 ,\u2_Display/n1119 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u5  (
    .a(\u2_Display/n1111 ),
    .b(1'b0),
    .c(\u2_Display/add38/c5 ),
    .o({\u2_Display/add38/c6 ,\u2_Display/n1119 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u6  (
    .a(\u2_Display/n1110 ),
    .b(1'b1),
    .c(\u2_Display/add38/c6 ),
    .o({\u2_Display/add38/c7 ,\u2_Display/n1119 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u7  (
    .a(\u2_Display/n1109 ),
    .b(1'b0),
    .c(\u2_Display/add38/c7 ),
    .o({\u2_Display/add38/c8 ,\u2_Display/n1119 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u8  (
    .a(\u2_Display/n1108 ),
    .b(1'b0),
    .c(\u2_Display/add38/c8 ),
    .o({\u2_Display/add38/c9 ,\u2_Display/n1119 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add38/u9  (
    .a(\u2_Display/n1107 ),
    .b(1'b0),
    .c(\u2_Display/add38/c9 ),
    .o({\u2_Display/add38/c10 ,\u2_Display/n1119 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add38/ucin  (
    .a(1'b1),
    .o({\u2_Display/add38/c0 ,open_n1180}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u0  (
    .a(\u2_Display/n1151 ),
    .b(1'b1),
    .c(\u2_Display/add39/c0 ),
    .o({\u2_Display/add39/c1 ,\u2_Display/n1154 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u1  (
    .a(\u2_Display/n1150 ),
    .b(1'b1),
    .c(\u2_Display/add39/c1 ),
    .o({\u2_Display/add39/c2 ,\u2_Display/n1154 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u10  (
    .a(\u2_Display/n1141 ),
    .b(1'b0),
    .c(\u2_Display/add39/c10 ),
    .o({\u2_Display/add39/c11 ,\u2_Display/n1154 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u11  (
    .a(\u2_Display/n1140 ),
    .b(1'b1),
    .c(\u2_Display/add39/c11 ),
    .o({\u2_Display/add39/c12 ,\u2_Display/n1154 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u12  (
    .a(\u2_Display/n1139 ),
    .b(1'b1),
    .c(\u2_Display/add39/c12 ),
    .o({\u2_Display/add39/c13 ,\u2_Display/n1154 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u13  (
    .a(\u2_Display/n1138 ),
    .b(1'b1),
    .c(\u2_Display/add39/c13 ),
    .o({\u2_Display/add39/c14 ,\u2_Display/n1154 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u14  (
    .a(\u2_Display/n1137 ),
    .b(1'b1),
    .c(\u2_Display/add39/c14 ),
    .o({\u2_Display/add39/c15 ,\u2_Display/n1154 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u15  (
    .a(\u2_Display/n1136 ),
    .b(1'b1),
    .c(\u2_Display/add39/c15 ),
    .o({\u2_Display/add39/c16 ,\u2_Display/n1154 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u16  (
    .a(\u2_Display/n1135 ),
    .b(1'b1),
    .c(\u2_Display/add39/c16 ),
    .o({\u2_Display/add39/c17 ,\u2_Display/n1154 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u17  (
    .a(\u2_Display/n1134 ),
    .b(1'b1),
    .c(\u2_Display/add39/c17 ),
    .o({\u2_Display/add39/c18 ,\u2_Display/n1154 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u18  (
    .a(\u2_Display/n1133 ),
    .b(1'b1),
    .c(\u2_Display/add39/c18 ),
    .o({\u2_Display/add39/c19 ,\u2_Display/n1154 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u19  (
    .a(\u2_Display/n1132 ),
    .b(1'b1),
    .c(\u2_Display/add39/c19 ),
    .o({\u2_Display/add39/c20 ,\u2_Display/n1154 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u2  (
    .a(\u2_Display/n1149 ),
    .b(1'b1),
    .c(\u2_Display/add39/c2 ),
    .o({\u2_Display/add39/c3 ,\u2_Display/n1154 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u20  (
    .a(\u2_Display/n1131 ),
    .b(1'b1),
    .c(\u2_Display/add39/c20 ),
    .o({\u2_Display/add39/c21 ,\u2_Display/n1154 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u21  (
    .a(\u2_Display/n1130 ),
    .b(1'b1),
    .c(\u2_Display/add39/c21 ),
    .o({\u2_Display/add39/c22 ,\u2_Display/n1154 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u22  (
    .a(\u2_Display/n1129 ),
    .b(1'b1),
    .c(\u2_Display/add39/c22 ),
    .o({\u2_Display/add39/c23 ,\u2_Display/n1154 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u23  (
    .a(\u2_Display/n1128 ),
    .b(1'b1),
    .c(\u2_Display/add39/c23 ),
    .o({\u2_Display/add39/c24 ,\u2_Display/n1154 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u24  (
    .a(\u2_Display/n1127 ),
    .b(1'b1),
    .c(\u2_Display/add39/c24 ),
    .o({\u2_Display/add39/c25 ,\u2_Display/n1154 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u25  (
    .a(\u2_Display/n1126 ),
    .b(1'b1),
    .c(\u2_Display/add39/c25 ),
    .o({\u2_Display/add39/c26 ,\u2_Display/n1154 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u26  (
    .a(\u2_Display/n1125 ),
    .b(1'b1),
    .c(\u2_Display/add39/c26 ),
    .o({\u2_Display/add39/c27 ,\u2_Display/n1154 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u27  (
    .a(\u2_Display/n1124 ),
    .b(1'b1),
    .c(\u2_Display/add39/c27 ),
    .o({\u2_Display/add39/c28 ,\u2_Display/n1154 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u28  (
    .a(\u2_Display/n1123 ),
    .b(1'b1),
    .c(\u2_Display/add39/c28 ),
    .o({\u2_Display/add39/c29 ,\u2_Display/n1154 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u29  (
    .a(\u2_Display/n1122 ),
    .b(1'b1),
    .c(\u2_Display/add39/c29 ),
    .o({\u2_Display/add39/c30 ,\u2_Display/n1154 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u3  (
    .a(\u2_Display/n1148 ),
    .b(1'b1),
    .c(\u2_Display/add39/c3 ),
    .o({\u2_Display/add39/c4 ,\u2_Display/n1154 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u30  (
    .a(\u2_Display/n1121 ),
    .b(1'b1),
    .c(\u2_Display/add39/c30 ),
    .o({\u2_Display/add39/c31 ,\u2_Display/n1154 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u31  (
    .a(\u2_Display/n1120 ),
    .b(1'b1),
    .c(\u2_Display/add39/c31 ),
    .o({open_n1181,\u2_Display/n1154 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u4  (
    .a(\u2_Display/n1147 ),
    .b(1'b0),
    .c(\u2_Display/add39/c4 ),
    .o({\u2_Display/add39/c5 ,\u2_Display/n1154 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u5  (
    .a(\u2_Display/n1146 ),
    .b(1'b1),
    .c(\u2_Display/add39/c5 ),
    .o({\u2_Display/add39/c6 ,\u2_Display/n1154 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u6  (
    .a(\u2_Display/n1145 ),
    .b(1'b0),
    .c(\u2_Display/add39/c6 ),
    .o({\u2_Display/add39/c7 ,\u2_Display/n1154 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u7  (
    .a(\u2_Display/n1144 ),
    .b(1'b0),
    .c(\u2_Display/add39/c7 ),
    .o({\u2_Display/add39/c8 ,\u2_Display/n1154 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u8  (
    .a(\u2_Display/n1143 ),
    .b(1'b0),
    .c(\u2_Display/add39/c8 ),
    .o({\u2_Display/add39/c9 ,\u2_Display/n1154 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add39/u9  (
    .a(\u2_Display/n1142 ),
    .b(1'b0),
    .c(\u2_Display/add39/c9 ),
    .o({\u2_Display/add39/c10 ,\u2_Display/n1154 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add39/ucin  (
    .a(1'b1),
    .o({\u2_Display/add39/c0 ,open_n1184}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add40/u0  (
    .a(\u2_Display/n1186 ),
    .b(1'b1),
    .c(\u2_Display/add40/c0 ),
    .o({\u2_Display/add40/c1 ,\u2_Display/n1189 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add40/u1  (
    .a(\u2_Display/n1185 ),
    .b(1'b1),
    .c(\u2_Display/add40/c1 ),
    .o({\u2_Display/add40/c2 ,\u2_Display/n1189 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add40/u2  (
    .a(\u2_Display/n1184 ),
    .b(1'b1),
    .c(\u2_Display/add40/c2 ),
    .o({\u2_Display/add40/c3 ,\u2_Display/n1189 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add40/u3  (
    .a(\u2_Display/n1183 ),
    .b(1'b0),
    .c(\u2_Display/add40/c3 ),
    .o({\u2_Display/add40/c4 ,\u2_Display/n1189 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add40/u4  (
    .a(\u2_Display/n1182 ),
    .b(1'b1),
    .c(\u2_Display/add40/c4 ),
    .o({\u2_Display/add40/c5 ,\u2_Display/n1189 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add40/u5  (
    .a(\u2_Display/n1181 ),
    .b(1'b0),
    .c(\u2_Display/add40/c5 ),
    .o({\u2_Display/add40/c6 ,\u2_Display/n1189 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add40/u6  (
    .a(\u2_Display/n1180 ),
    .b(1'b0),
    .c(\u2_Display/add40/c6 ),
    .o({\u2_Display/add40/c7 ,\u2_Display/n1189 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add40/u7  (
    .a(\u2_Display/n1179 ),
    .b(1'b0),
    .c(\u2_Display/add40/c7 ),
    .o({\u2_Display/add40/c8 ,\u2_Display/n1189 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add40/u8  (
    .a(\u2_Display/n1178 ),
    .b(1'b0),
    .c(\u2_Display/add40/c8 ),
    .o({\u2_Display/add40/c9 ,\u2_Display/n1189 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add40/u9  (
    .a(\u2_Display/n1177 ),
    .b(1'b0),
    .c(\u2_Display/add40/c9 ),
    .o({open_n1185,\u2_Display/n1189 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add40/ucin  (
    .a(1'b1),
    .o({\u2_Display/add40/c0 ,open_n1188}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add4_2/u0  (
    .a(1'b1),
    .b(\u2_Display/i [7]),
    .c(\u2_Display/add4_2/c0 ),
    .o({\u2_Display/add4_2/c1 ,\u2_Display/n94 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add4_2/u1  (
    .a(1'b0),
    .b(\u2_Display/i [8]),
    .c(\u2_Display/add4_2/c1 ),
    .o({\u2_Display/add4_2/c2 ,\u2_Display/n94 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add4_2/u2  (
    .a(1'b1),
    .b(\u2_Display/i [9]),
    .c(\u2_Display/add4_2/c2 ),
    .o({\u2_Display/add4_2/c3 ,\u2_Display/n94 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add4_2/u3  (
    .a(1'b0),
    .b(\u2_Display/i [10]),
    .c(\u2_Display/add4_2/c3 ),
    .o({\u2_Display/add4_2/c4 ,\u2_Display/n94 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add4_2/ucin  (
    .a(1'b0),
    .o({\u2_Display/add4_2/c0 ,open_n1191}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add4_2/ucout  (
    .c(\u2_Display/add4_2/c4 ),
    .o({open_n1194,\u2_Display/add4_2_co }));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u0  (
    .a(\u2_Display/counta [0]),
    .b(1'b1),
    .c(\u2_Display/add51/c0 ),
    .o({\u2_Display/add51/c1 ,\u2_Display/n1542 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u1  (
    .a(\u2_Display/counta [1]),
    .b(1'b1),
    .c(\u2_Display/add51/c1 ),
    .o({\u2_Display/add51/c2 ,\u2_Display/n1542 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u10  (
    .a(\u2_Display/counta [10]),
    .b(1'b1),
    .c(\u2_Display/add51/c10 ),
    .o({\u2_Display/add51/c11 ,\u2_Display/n1542 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u11  (
    .a(\u2_Display/counta [11]),
    .b(1'b1),
    .c(\u2_Display/add51/c11 ),
    .o({\u2_Display/add51/c12 ,\u2_Display/n1542 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u12  (
    .a(\u2_Display/counta [12]),
    .b(1'b1),
    .c(\u2_Display/add51/c12 ),
    .o({\u2_Display/add51/c13 ,\u2_Display/n1542 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u13  (
    .a(\u2_Display/counta [13]),
    .b(1'b1),
    .c(\u2_Display/add51/c13 ),
    .o({\u2_Display/add51/c14 ,\u2_Display/n1542 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u14  (
    .a(\u2_Display/counta [14]),
    .b(1'b1),
    .c(\u2_Display/add51/c14 ),
    .o({\u2_Display/add51/c15 ,\u2_Display/n1542 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u15  (
    .a(\u2_Display/counta [15]),
    .b(1'b1),
    .c(\u2_Display/add51/c15 ),
    .o({\u2_Display/add51/c16 ,\u2_Display/n1542 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u16  (
    .a(\u2_Display/counta [16]),
    .b(1'b1),
    .c(\u2_Display/add51/c16 ),
    .o({\u2_Display/add51/c17 ,\u2_Display/n1542 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u17  (
    .a(\u2_Display/counta [17]),
    .b(1'b1),
    .c(\u2_Display/add51/c17 ),
    .o({\u2_Display/add51/c18 ,\u2_Display/n1542 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u18  (
    .a(\u2_Display/counta [18]),
    .b(1'b1),
    .c(\u2_Display/add51/c18 ),
    .o({\u2_Display/add51/c19 ,\u2_Display/n1542 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u19  (
    .a(\u2_Display/counta [19]),
    .b(1'b1),
    .c(\u2_Display/add51/c19 ),
    .o({\u2_Display/add51/c20 ,\u2_Display/n1542 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u2  (
    .a(\u2_Display/counta [2]),
    .b(1'b1),
    .c(\u2_Display/add51/c2 ),
    .o({\u2_Display/add51/c3 ,\u2_Display/n1542 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u20  (
    .a(\u2_Display/counta [20]),
    .b(1'b1),
    .c(\u2_Display/add51/c20 ),
    .o({\u2_Display/add51/c21 ,\u2_Display/n1542 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u21  (
    .a(\u2_Display/counta [21]),
    .b(1'b1),
    .c(\u2_Display/add51/c21 ),
    .o({\u2_Display/add51/c22 ,\u2_Display/n1542 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u22  (
    .a(\u2_Display/counta [22]),
    .b(1'b1),
    .c(\u2_Display/add51/c22 ),
    .o({\u2_Display/add51/c23 ,\u2_Display/n1542 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u23  (
    .a(\u2_Display/counta [23]),
    .b(1'b1),
    .c(\u2_Display/add51/c23 ),
    .o({\u2_Display/add51/c24 ,\u2_Display/n1542 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u24  (
    .a(\u2_Display/counta [24]),
    .b(1'b0),
    .c(\u2_Display/add51/c24 ),
    .o({\u2_Display/add51/c25 ,\u2_Display/n1542 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u25  (
    .a(\u2_Display/counta [25]),
    .b(1'b1),
    .c(\u2_Display/add51/c25 ),
    .o({\u2_Display/add51/c26 ,\u2_Display/n1542 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u26  (
    .a(\u2_Display/counta [26]),
    .b(1'b1),
    .c(\u2_Display/add51/c26 ),
    .o({\u2_Display/add51/c27 ,\u2_Display/n1542 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u27  (
    .a(\u2_Display/counta [27]),
    .b(1'b1),
    .c(\u2_Display/add51/c27 ),
    .o({\u2_Display/add51/c28 ,\u2_Display/n1542 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u28  (
    .a(\u2_Display/counta [28]),
    .b(1'b1),
    .c(\u2_Display/add51/c28 ),
    .o({\u2_Display/add51/c29 ,\u2_Display/n1542 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u29  (
    .a(\u2_Display/counta [29]),
    .b(1'b0),
    .c(\u2_Display/add51/c29 ),
    .o({\u2_Display/add51/c30 ,\u2_Display/n1542 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u3  (
    .a(\u2_Display/counta [3]),
    .b(1'b1),
    .c(\u2_Display/add51/c3 ),
    .o({\u2_Display/add51/c4 ,\u2_Display/n1542 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u30  (
    .a(\u2_Display/counta [30]),
    .b(1'b0),
    .c(\u2_Display/add51/c30 ),
    .o({\u2_Display/add51/c31 ,\u2_Display/n1542 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u31  (
    .a(\u2_Display/counta [31]),
    .b(1'b0),
    .c(\u2_Display/add51/c31 ),
    .o({open_n1195,\u2_Display/n1542 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u4  (
    .a(\u2_Display/counta [4]),
    .b(1'b1),
    .c(\u2_Display/add51/c4 ),
    .o({\u2_Display/add51/c5 ,\u2_Display/n1542 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u5  (
    .a(\u2_Display/counta [5]),
    .b(1'b1),
    .c(\u2_Display/add51/c5 ),
    .o({\u2_Display/add51/c6 ,\u2_Display/n1542 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u6  (
    .a(\u2_Display/counta [6]),
    .b(1'b1),
    .c(\u2_Display/add51/c6 ),
    .o({\u2_Display/add51/c7 ,\u2_Display/n1542 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u7  (
    .a(\u2_Display/counta [7]),
    .b(1'b1),
    .c(\u2_Display/add51/c7 ),
    .o({\u2_Display/add51/c8 ,\u2_Display/n1542 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u8  (
    .a(\u2_Display/counta [8]),
    .b(1'b1),
    .c(\u2_Display/add51/c8 ),
    .o({\u2_Display/add51/c9 ,\u2_Display/n1542 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add51/u9  (
    .a(\u2_Display/counta [9]),
    .b(1'b1),
    .c(\u2_Display/add51/c9 ),
    .o({\u2_Display/add51/c10 ,\u2_Display/n1542 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add51/ucin  (
    .a(1'b1),
    .o({\u2_Display/add51/c0 ,open_n1198}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u0  (
    .a(\u2_Display/n1574 ),
    .b(1'b1),
    .c(\u2_Display/add52/c0 ),
    .o({\u2_Display/add52/c1 ,\u2_Display/n1577 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u1  (
    .a(\u2_Display/n1573 ),
    .b(1'b1),
    .c(\u2_Display/add52/c1 ),
    .o({\u2_Display/add52/c2 ,\u2_Display/n1577 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u10  (
    .a(\u2_Display/n1564 ),
    .b(1'b1),
    .c(\u2_Display/add52/c10 ),
    .o({\u2_Display/add52/c11 ,\u2_Display/n1577 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u11  (
    .a(\u2_Display/n1563 ),
    .b(1'b1),
    .c(\u2_Display/add52/c11 ),
    .o({\u2_Display/add52/c12 ,\u2_Display/n1577 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u12  (
    .a(\u2_Display/n1562 ),
    .b(1'b1),
    .c(\u2_Display/add52/c12 ),
    .o({\u2_Display/add52/c13 ,\u2_Display/n1577 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u13  (
    .a(\u2_Display/n1561 ),
    .b(1'b1),
    .c(\u2_Display/add52/c13 ),
    .o({\u2_Display/add52/c14 ,\u2_Display/n1577 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u14  (
    .a(\u2_Display/n1560 ),
    .b(1'b1),
    .c(\u2_Display/add52/c14 ),
    .o({\u2_Display/add52/c15 ,\u2_Display/n1577 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u15  (
    .a(\u2_Display/n1559 ),
    .b(1'b1),
    .c(\u2_Display/add52/c15 ),
    .o({\u2_Display/add52/c16 ,\u2_Display/n1577 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u16  (
    .a(\u2_Display/n1558 ),
    .b(1'b1),
    .c(\u2_Display/add52/c16 ),
    .o({\u2_Display/add52/c17 ,\u2_Display/n1577 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u17  (
    .a(\u2_Display/n1557 ),
    .b(1'b1),
    .c(\u2_Display/add52/c17 ),
    .o({\u2_Display/add52/c18 ,\u2_Display/n1577 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u18  (
    .a(\u2_Display/n1556 ),
    .b(1'b1),
    .c(\u2_Display/add52/c18 ),
    .o({\u2_Display/add52/c19 ,\u2_Display/n1577 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u19  (
    .a(\u2_Display/n1555 ),
    .b(1'b1),
    .c(\u2_Display/add52/c19 ),
    .o({\u2_Display/add52/c20 ,\u2_Display/n1577 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u2  (
    .a(\u2_Display/n1572 ),
    .b(1'b1),
    .c(\u2_Display/add52/c2 ),
    .o({\u2_Display/add52/c3 ,\u2_Display/n1577 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u20  (
    .a(\u2_Display/n1554 ),
    .b(1'b1),
    .c(\u2_Display/add52/c20 ),
    .o({\u2_Display/add52/c21 ,\u2_Display/n1577 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u21  (
    .a(\u2_Display/n1553 ),
    .b(1'b1),
    .c(\u2_Display/add52/c21 ),
    .o({\u2_Display/add52/c22 ,\u2_Display/n1577 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u22  (
    .a(\u2_Display/n1552 ),
    .b(1'b1),
    .c(\u2_Display/add52/c22 ),
    .o({\u2_Display/add52/c23 ,\u2_Display/n1577 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u23  (
    .a(\u2_Display/n1551 ),
    .b(1'b0),
    .c(\u2_Display/add52/c23 ),
    .o({\u2_Display/add52/c24 ,\u2_Display/n1577 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u24  (
    .a(\u2_Display/n1550 ),
    .b(1'b1),
    .c(\u2_Display/add52/c24 ),
    .o({\u2_Display/add52/c25 ,\u2_Display/n1577 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u25  (
    .a(\u2_Display/n1549 ),
    .b(1'b1),
    .c(\u2_Display/add52/c25 ),
    .o({\u2_Display/add52/c26 ,\u2_Display/n1577 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u26  (
    .a(\u2_Display/n1548 ),
    .b(1'b1),
    .c(\u2_Display/add52/c26 ),
    .o({\u2_Display/add52/c27 ,\u2_Display/n1577 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u27  (
    .a(\u2_Display/n1547 ),
    .b(1'b1),
    .c(\u2_Display/add52/c27 ),
    .o({\u2_Display/add52/c28 ,\u2_Display/n1577 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u28  (
    .a(\u2_Display/n1546 ),
    .b(1'b0),
    .c(\u2_Display/add52/c28 ),
    .o({\u2_Display/add52/c29 ,\u2_Display/n1577 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u29  (
    .a(\u2_Display/n1545 ),
    .b(1'b0),
    .c(\u2_Display/add52/c29 ),
    .o({\u2_Display/add52/c30 ,\u2_Display/n1577 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u3  (
    .a(\u2_Display/n1571 ),
    .b(1'b1),
    .c(\u2_Display/add52/c3 ),
    .o({\u2_Display/add52/c4 ,\u2_Display/n1577 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u30  (
    .a(\u2_Display/n1544 ),
    .b(1'b0),
    .c(\u2_Display/add52/c30 ),
    .o({\u2_Display/add52/c31 ,\u2_Display/n1577 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u31  (
    .a(\u2_Display/n1543 ),
    .b(1'b1),
    .c(\u2_Display/add52/c31 ),
    .o({open_n1199,\u2_Display/n1577 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u4  (
    .a(\u2_Display/n1570 ),
    .b(1'b1),
    .c(\u2_Display/add52/c4 ),
    .o({\u2_Display/add52/c5 ,\u2_Display/n1577 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u5  (
    .a(\u2_Display/n1569 ),
    .b(1'b1),
    .c(\u2_Display/add52/c5 ),
    .o({\u2_Display/add52/c6 ,\u2_Display/n1577 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u6  (
    .a(\u2_Display/n1568 ),
    .b(1'b1),
    .c(\u2_Display/add52/c6 ),
    .o({\u2_Display/add52/c7 ,\u2_Display/n1577 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u7  (
    .a(\u2_Display/n1567 ),
    .b(1'b1),
    .c(\u2_Display/add52/c7 ),
    .o({\u2_Display/add52/c8 ,\u2_Display/n1577 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u8  (
    .a(\u2_Display/n1566 ),
    .b(1'b1),
    .c(\u2_Display/add52/c8 ),
    .o({\u2_Display/add52/c9 ,\u2_Display/n1577 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add52/u9  (
    .a(\u2_Display/n1565 ),
    .b(1'b1),
    .c(\u2_Display/add52/c9 ),
    .o({\u2_Display/add52/c10 ,\u2_Display/n1577 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add52/ucin  (
    .a(1'b1),
    .o({\u2_Display/add52/c0 ,open_n1202}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u0  (
    .a(\u2_Display/n1609 ),
    .b(1'b1),
    .c(\u2_Display/add53/c0 ),
    .o({\u2_Display/add53/c1 ,\u2_Display/n1612 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u1  (
    .a(\u2_Display/n1608 ),
    .b(1'b1),
    .c(\u2_Display/add53/c1 ),
    .o({\u2_Display/add53/c2 ,\u2_Display/n1612 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u10  (
    .a(\u2_Display/n1599 ),
    .b(1'b1),
    .c(\u2_Display/add53/c10 ),
    .o({\u2_Display/add53/c11 ,\u2_Display/n1612 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u11  (
    .a(\u2_Display/n1598 ),
    .b(1'b1),
    .c(\u2_Display/add53/c11 ),
    .o({\u2_Display/add53/c12 ,\u2_Display/n1612 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u12  (
    .a(\u2_Display/n1597 ),
    .b(1'b1),
    .c(\u2_Display/add53/c12 ),
    .o({\u2_Display/add53/c13 ,\u2_Display/n1612 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u13  (
    .a(\u2_Display/n1596 ),
    .b(1'b1),
    .c(\u2_Display/add53/c13 ),
    .o({\u2_Display/add53/c14 ,\u2_Display/n1612 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u14  (
    .a(\u2_Display/n1595 ),
    .b(1'b1),
    .c(\u2_Display/add53/c14 ),
    .o({\u2_Display/add53/c15 ,\u2_Display/n1612 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u15  (
    .a(\u2_Display/n1594 ),
    .b(1'b1),
    .c(\u2_Display/add53/c15 ),
    .o({\u2_Display/add53/c16 ,\u2_Display/n1612 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u16  (
    .a(\u2_Display/n1593 ),
    .b(1'b1),
    .c(\u2_Display/add53/c16 ),
    .o({\u2_Display/add53/c17 ,\u2_Display/n1612 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u17  (
    .a(\u2_Display/n1592 ),
    .b(1'b1),
    .c(\u2_Display/add53/c17 ),
    .o({\u2_Display/add53/c18 ,\u2_Display/n1612 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u18  (
    .a(\u2_Display/n1591 ),
    .b(1'b1),
    .c(\u2_Display/add53/c18 ),
    .o({\u2_Display/add53/c19 ,\u2_Display/n1612 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u19  (
    .a(\u2_Display/n1590 ),
    .b(1'b1),
    .c(\u2_Display/add53/c19 ),
    .o({\u2_Display/add53/c20 ,\u2_Display/n1612 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u2  (
    .a(\u2_Display/n1607 ),
    .b(1'b1),
    .c(\u2_Display/add53/c2 ),
    .o({\u2_Display/add53/c3 ,\u2_Display/n1612 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u20  (
    .a(\u2_Display/n1589 ),
    .b(1'b1),
    .c(\u2_Display/add53/c20 ),
    .o({\u2_Display/add53/c21 ,\u2_Display/n1612 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u21  (
    .a(\u2_Display/n1588 ),
    .b(1'b1),
    .c(\u2_Display/add53/c21 ),
    .o({\u2_Display/add53/c22 ,\u2_Display/n1612 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u22  (
    .a(\u2_Display/n1587 ),
    .b(1'b0),
    .c(\u2_Display/add53/c22 ),
    .o({\u2_Display/add53/c23 ,\u2_Display/n1612 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u23  (
    .a(\u2_Display/n1586 ),
    .b(1'b1),
    .c(\u2_Display/add53/c23 ),
    .o({\u2_Display/add53/c24 ,\u2_Display/n1612 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u24  (
    .a(\u2_Display/n1585 ),
    .b(1'b1),
    .c(\u2_Display/add53/c24 ),
    .o({\u2_Display/add53/c25 ,\u2_Display/n1612 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u25  (
    .a(\u2_Display/n1584 ),
    .b(1'b1),
    .c(\u2_Display/add53/c25 ),
    .o({\u2_Display/add53/c26 ,\u2_Display/n1612 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u26  (
    .a(\u2_Display/n1583 ),
    .b(1'b1),
    .c(\u2_Display/add53/c26 ),
    .o({\u2_Display/add53/c27 ,\u2_Display/n1612 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u27  (
    .a(\u2_Display/n1582 ),
    .b(1'b0),
    .c(\u2_Display/add53/c27 ),
    .o({\u2_Display/add53/c28 ,\u2_Display/n1612 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u28  (
    .a(\u2_Display/n1581 ),
    .b(1'b0),
    .c(\u2_Display/add53/c28 ),
    .o({\u2_Display/add53/c29 ,\u2_Display/n1612 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u29  (
    .a(\u2_Display/n1580 ),
    .b(1'b0),
    .c(\u2_Display/add53/c29 ),
    .o({\u2_Display/add53/c30 ,\u2_Display/n1612 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u3  (
    .a(\u2_Display/n1606 ),
    .b(1'b1),
    .c(\u2_Display/add53/c3 ),
    .o({\u2_Display/add53/c4 ,\u2_Display/n1612 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u30  (
    .a(\u2_Display/n1579 ),
    .b(1'b1),
    .c(\u2_Display/add53/c30 ),
    .o({\u2_Display/add53/c31 ,\u2_Display/n1612 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u31  (
    .a(\u2_Display/n1578 ),
    .b(1'b1),
    .c(\u2_Display/add53/c31 ),
    .o({open_n1203,\u2_Display/n1612 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u4  (
    .a(\u2_Display/n1605 ),
    .b(1'b1),
    .c(\u2_Display/add53/c4 ),
    .o({\u2_Display/add53/c5 ,\u2_Display/n1612 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u5  (
    .a(\u2_Display/n1604 ),
    .b(1'b1),
    .c(\u2_Display/add53/c5 ),
    .o({\u2_Display/add53/c6 ,\u2_Display/n1612 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u6  (
    .a(\u2_Display/n1603 ),
    .b(1'b1),
    .c(\u2_Display/add53/c6 ),
    .o({\u2_Display/add53/c7 ,\u2_Display/n1612 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u7  (
    .a(\u2_Display/n1602 ),
    .b(1'b1),
    .c(\u2_Display/add53/c7 ),
    .o({\u2_Display/add53/c8 ,\u2_Display/n1612 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u8  (
    .a(\u2_Display/n1601 ),
    .b(1'b1),
    .c(\u2_Display/add53/c8 ),
    .o({\u2_Display/add53/c9 ,\u2_Display/n1612 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add53/u9  (
    .a(\u2_Display/n1600 ),
    .b(1'b1),
    .c(\u2_Display/add53/c9 ),
    .o({\u2_Display/add53/c10 ,\u2_Display/n1612 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add53/ucin  (
    .a(1'b1),
    .o({\u2_Display/add53/c0 ,open_n1206}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u0  (
    .a(\u2_Display/n1644 ),
    .b(1'b1),
    .c(\u2_Display/add54/c0 ),
    .o({\u2_Display/add54/c1 ,\u2_Display/n1647 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u1  (
    .a(\u2_Display/n1643 ),
    .b(1'b1),
    .c(\u2_Display/add54/c1 ),
    .o({\u2_Display/add54/c2 ,\u2_Display/n1647 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u10  (
    .a(\u2_Display/n1634 ),
    .b(1'b1),
    .c(\u2_Display/add54/c10 ),
    .o({\u2_Display/add54/c11 ,\u2_Display/n1647 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u11  (
    .a(\u2_Display/n1633 ),
    .b(1'b1),
    .c(\u2_Display/add54/c11 ),
    .o({\u2_Display/add54/c12 ,\u2_Display/n1647 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u12  (
    .a(\u2_Display/n1632 ),
    .b(1'b1),
    .c(\u2_Display/add54/c12 ),
    .o({\u2_Display/add54/c13 ,\u2_Display/n1647 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u13  (
    .a(\u2_Display/n1631 ),
    .b(1'b1),
    .c(\u2_Display/add54/c13 ),
    .o({\u2_Display/add54/c14 ,\u2_Display/n1647 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u14  (
    .a(\u2_Display/n1630 ),
    .b(1'b1),
    .c(\u2_Display/add54/c14 ),
    .o({\u2_Display/add54/c15 ,\u2_Display/n1647 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u15  (
    .a(\u2_Display/n1629 ),
    .b(1'b1),
    .c(\u2_Display/add54/c15 ),
    .o({\u2_Display/add54/c16 ,\u2_Display/n1647 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u16  (
    .a(\u2_Display/n1628 ),
    .b(1'b1),
    .c(\u2_Display/add54/c16 ),
    .o({\u2_Display/add54/c17 ,\u2_Display/n1647 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u17  (
    .a(\u2_Display/n1627 ),
    .b(1'b1),
    .c(\u2_Display/add54/c17 ),
    .o({\u2_Display/add54/c18 ,\u2_Display/n1647 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u18  (
    .a(\u2_Display/n1626 ),
    .b(1'b1),
    .c(\u2_Display/add54/c18 ),
    .o({\u2_Display/add54/c19 ,\u2_Display/n1647 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u19  (
    .a(\u2_Display/n1625 ),
    .b(1'b1),
    .c(\u2_Display/add54/c19 ),
    .o({\u2_Display/add54/c20 ,\u2_Display/n1647 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u2  (
    .a(\u2_Display/n1642 ),
    .b(1'b1),
    .c(\u2_Display/add54/c2 ),
    .o({\u2_Display/add54/c3 ,\u2_Display/n1647 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u20  (
    .a(\u2_Display/n1624 ),
    .b(1'b1),
    .c(\u2_Display/add54/c20 ),
    .o({\u2_Display/add54/c21 ,\u2_Display/n1647 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u21  (
    .a(\u2_Display/n1623 ),
    .b(1'b0),
    .c(\u2_Display/add54/c21 ),
    .o({\u2_Display/add54/c22 ,\u2_Display/n1647 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u22  (
    .a(\u2_Display/n1622 ),
    .b(1'b1),
    .c(\u2_Display/add54/c22 ),
    .o({\u2_Display/add54/c23 ,\u2_Display/n1647 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u23  (
    .a(\u2_Display/n1621 ),
    .b(1'b1),
    .c(\u2_Display/add54/c23 ),
    .o({\u2_Display/add54/c24 ,\u2_Display/n1647 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u24  (
    .a(\u2_Display/n1620 ),
    .b(1'b1),
    .c(\u2_Display/add54/c24 ),
    .o({\u2_Display/add54/c25 ,\u2_Display/n1647 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u25  (
    .a(\u2_Display/n1619 ),
    .b(1'b1),
    .c(\u2_Display/add54/c25 ),
    .o({\u2_Display/add54/c26 ,\u2_Display/n1647 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u26  (
    .a(\u2_Display/n1618 ),
    .b(1'b0),
    .c(\u2_Display/add54/c26 ),
    .o({\u2_Display/add54/c27 ,\u2_Display/n1647 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u27  (
    .a(\u2_Display/n1617 ),
    .b(1'b0),
    .c(\u2_Display/add54/c27 ),
    .o({\u2_Display/add54/c28 ,\u2_Display/n1647 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u28  (
    .a(\u2_Display/n1616 ),
    .b(1'b0),
    .c(\u2_Display/add54/c28 ),
    .o({\u2_Display/add54/c29 ,\u2_Display/n1647 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u29  (
    .a(\u2_Display/n1615 ),
    .b(1'b1),
    .c(\u2_Display/add54/c29 ),
    .o({\u2_Display/add54/c30 ,\u2_Display/n1647 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u3  (
    .a(\u2_Display/n1641 ),
    .b(1'b1),
    .c(\u2_Display/add54/c3 ),
    .o({\u2_Display/add54/c4 ,\u2_Display/n1647 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u30  (
    .a(\u2_Display/n1614 ),
    .b(1'b1),
    .c(\u2_Display/add54/c30 ),
    .o({\u2_Display/add54/c31 ,\u2_Display/n1647 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u31  (
    .a(\u2_Display/n1613 ),
    .b(1'b1),
    .c(\u2_Display/add54/c31 ),
    .o({open_n1207,\u2_Display/n1647 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u4  (
    .a(\u2_Display/n1640 ),
    .b(1'b1),
    .c(\u2_Display/add54/c4 ),
    .o({\u2_Display/add54/c5 ,\u2_Display/n1647 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u5  (
    .a(\u2_Display/n1639 ),
    .b(1'b1),
    .c(\u2_Display/add54/c5 ),
    .o({\u2_Display/add54/c6 ,\u2_Display/n1647 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u6  (
    .a(\u2_Display/n1638 ),
    .b(1'b1),
    .c(\u2_Display/add54/c6 ),
    .o({\u2_Display/add54/c7 ,\u2_Display/n1647 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u7  (
    .a(\u2_Display/n1637 ),
    .b(1'b1),
    .c(\u2_Display/add54/c7 ),
    .o({\u2_Display/add54/c8 ,\u2_Display/n1647 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u8  (
    .a(\u2_Display/n1636 ),
    .b(1'b1),
    .c(\u2_Display/add54/c8 ),
    .o({\u2_Display/add54/c9 ,\u2_Display/n1647 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add54/u9  (
    .a(\u2_Display/n1635 ),
    .b(1'b1),
    .c(\u2_Display/add54/c9 ),
    .o({\u2_Display/add54/c10 ,\u2_Display/n1647 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add54/ucin  (
    .a(1'b1),
    .o({\u2_Display/add54/c0 ,open_n1210}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u0  (
    .a(\u2_Display/n1679 ),
    .b(1'b1),
    .c(\u2_Display/add55/c0 ),
    .o({\u2_Display/add55/c1 ,\u2_Display/n1682 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u1  (
    .a(\u2_Display/n1678 ),
    .b(1'b1),
    .c(\u2_Display/add55/c1 ),
    .o({\u2_Display/add55/c2 ,\u2_Display/n1682 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u10  (
    .a(\u2_Display/n1669 ),
    .b(1'b1),
    .c(\u2_Display/add55/c10 ),
    .o({\u2_Display/add55/c11 ,\u2_Display/n1682 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u11  (
    .a(\u2_Display/n1668 ),
    .b(1'b1),
    .c(\u2_Display/add55/c11 ),
    .o({\u2_Display/add55/c12 ,\u2_Display/n1682 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u12  (
    .a(\u2_Display/n1667 ),
    .b(1'b1),
    .c(\u2_Display/add55/c12 ),
    .o({\u2_Display/add55/c13 ,\u2_Display/n1682 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u13  (
    .a(\u2_Display/n1666 ),
    .b(1'b1),
    .c(\u2_Display/add55/c13 ),
    .o({\u2_Display/add55/c14 ,\u2_Display/n1682 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u14  (
    .a(\u2_Display/n1665 ),
    .b(1'b1),
    .c(\u2_Display/add55/c14 ),
    .o({\u2_Display/add55/c15 ,\u2_Display/n1682 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u15  (
    .a(\u2_Display/n1664 ),
    .b(1'b1),
    .c(\u2_Display/add55/c15 ),
    .o({\u2_Display/add55/c16 ,\u2_Display/n1682 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u16  (
    .a(\u2_Display/n1663 ),
    .b(1'b1),
    .c(\u2_Display/add55/c16 ),
    .o({\u2_Display/add55/c17 ,\u2_Display/n1682 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u17  (
    .a(\u2_Display/n1662 ),
    .b(1'b1),
    .c(\u2_Display/add55/c17 ),
    .o({\u2_Display/add55/c18 ,\u2_Display/n1682 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u18  (
    .a(\u2_Display/n1661 ),
    .b(1'b1),
    .c(\u2_Display/add55/c18 ),
    .o({\u2_Display/add55/c19 ,\u2_Display/n1682 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u19  (
    .a(\u2_Display/n1660 ),
    .b(1'b1),
    .c(\u2_Display/add55/c19 ),
    .o({\u2_Display/add55/c20 ,\u2_Display/n1682 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u2  (
    .a(\u2_Display/n1677 ),
    .b(1'b1),
    .c(\u2_Display/add55/c2 ),
    .o({\u2_Display/add55/c3 ,\u2_Display/n1682 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u20  (
    .a(\u2_Display/n1659 ),
    .b(1'b0),
    .c(\u2_Display/add55/c20 ),
    .o({\u2_Display/add55/c21 ,\u2_Display/n1682 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u21  (
    .a(\u2_Display/n1658 ),
    .b(1'b1),
    .c(\u2_Display/add55/c21 ),
    .o({\u2_Display/add55/c22 ,\u2_Display/n1682 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u22  (
    .a(\u2_Display/n1657 ),
    .b(1'b1),
    .c(\u2_Display/add55/c22 ),
    .o({\u2_Display/add55/c23 ,\u2_Display/n1682 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u23  (
    .a(\u2_Display/n1656 ),
    .b(1'b1),
    .c(\u2_Display/add55/c23 ),
    .o({\u2_Display/add55/c24 ,\u2_Display/n1682 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u24  (
    .a(\u2_Display/n1655 ),
    .b(1'b1),
    .c(\u2_Display/add55/c24 ),
    .o({\u2_Display/add55/c25 ,\u2_Display/n1682 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u25  (
    .a(\u2_Display/n1654 ),
    .b(1'b0),
    .c(\u2_Display/add55/c25 ),
    .o({\u2_Display/add55/c26 ,\u2_Display/n1682 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u26  (
    .a(\u2_Display/n1653 ),
    .b(1'b0),
    .c(\u2_Display/add55/c26 ),
    .o({\u2_Display/add55/c27 ,\u2_Display/n1682 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u27  (
    .a(\u2_Display/n1652 ),
    .b(1'b0),
    .c(\u2_Display/add55/c27 ),
    .o({\u2_Display/add55/c28 ,\u2_Display/n1682 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u28  (
    .a(\u2_Display/n1651 ),
    .b(1'b1),
    .c(\u2_Display/add55/c28 ),
    .o({\u2_Display/add55/c29 ,\u2_Display/n1682 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u29  (
    .a(\u2_Display/n1650 ),
    .b(1'b1),
    .c(\u2_Display/add55/c29 ),
    .o({\u2_Display/add55/c30 ,\u2_Display/n1682 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u3  (
    .a(\u2_Display/n1676 ),
    .b(1'b1),
    .c(\u2_Display/add55/c3 ),
    .o({\u2_Display/add55/c4 ,\u2_Display/n1682 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u30  (
    .a(\u2_Display/n1649 ),
    .b(1'b1),
    .c(\u2_Display/add55/c30 ),
    .o({\u2_Display/add55/c31 ,\u2_Display/n1682 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u31  (
    .a(\u2_Display/n1648 ),
    .b(1'b1),
    .c(\u2_Display/add55/c31 ),
    .o({open_n1211,\u2_Display/n1682 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u4  (
    .a(\u2_Display/n1675 ),
    .b(1'b1),
    .c(\u2_Display/add55/c4 ),
    .o({\u2_Display/add55/c5 ,\u2_Display/n1682 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u5  (
    .a(\u2_Display/n1674 ),
    .b(1'b1),
    .c(\u2_Display/add55/c5 ),
    .o({\u2_Display/add55/c6 ,\u2_Display/n1682 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u6  (
    .a(\u2_Display/n1673 ),
    .b(1'b1),
    .c(\u2_Display/add55/c6 ),
    .o({\u2_Display/add55/c7 ,\u2_Display/n1682 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u7  (
    .a(\u2_Display/n1672 ),
    .b(1'b1),
    .c(\u2_Display/add55/c7 ),
    .o({\u2_Display/add55/c8 ,\u2_Display/n1682 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u8  (
    .a(\u2_Display/n1671 ),
    .b(1'b1),
    .c(\u2_Display/add55/c8 ),
    .o({\u2_Display/add55/c9 ,\u2_Display/n1682 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add55/u9  (
    .a(\u2_Display/n1670 ),
    .b(1'b1),
    .c(\u2_Display/add55/c9 ),
    .o({\u2_Display/add55/c10 ,\u2_Display/n1682 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add55/ucin  (
    .a(1'b1),
    .o({\u2_Display/add55/c0 ,open_n1214}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u0  (
    .a(\u2_Display/n1714 ),
    .b(1'b1),
    .c(\u2_Display/add56/c0 ),
    .o({\u2_Display/add56/c1 ,\u2_Display/n1717 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u1  (
    .a(\u2_Display/n1713 ),
    .b(1'b1),
    .c(\u2_Display/add56/c1 ),
    .o({\u2_Display/add56/c2 ,\u2_Display/n1717 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u10  (
    .a(\u2_Display/n1704 ),
    .b(1'b1),
    .c(\u2_Display/add56/c10 ),
    .o({\u2_Display/add56/c11 ,\u2_Display/n1717 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u11  (
    .a(\u2_Display/n1703 ),
    .b(1'b1),
    .c(\u2_Display/add56/c11 ),
    .o({\u2_Display/add56/c12 ,\u2_Display/n1717 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u12  (
    .a(\u2_Display/n1702 ),
    .b(1'b1),
    .c(\u2_Display/add56/c12 ),
    .o({\u2_Display/add56/c13 ,\u2_Display/n1717 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u13  (
    .a(\u2_Display/n1701 ),
    .b(1'b1),
    .c(\u2_Display/add56/c13 ),
    .o({\u2_Display/add56/c14 ,\u2_Display/n1717 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u14  (
    .a(\u2_Display/n1700 ),
    .b(1'b1),
    .c(\u2_Display/add56/c14 ),
    .o({\u2_Display/add56/c15 ,\u2_Display/n1717 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u15  (
    .a(\u2_Display/n1699 ),
    .b(1'b1),
    .c(\u2_Display/add56/c15 ),
    .o({\u2_Display/add56/c16 ,\u2_Display/n1717 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u16  (
    .a(\u2_Display/n1698 ),
    .b(1'b1),
    .c(\u2_Display/add56/c16 ),
    .o({\u2_Display/add56/c17 ,\u2_Display/n1717 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u17  (
    .a(\u2_Display/n1697 ),
    .b(1'b1),
    .c(\u2_Display/add56/c17 ),
    .o({\u2_Display/add56/c18 ,\u2_Display/n1717 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u18  (
    .a(\u2_Display/n1696 ),
    .b(1'b1),
    .c(\u2_Display/add56/c18 ),
    .o({\u2_Display/add56/c19 ,\u2_Display/n1717 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u19  (
    .a(\u2_Display/n1695 ),
    .b(1'b0),
    .c(\u2_Display/add56/c19 ),
    .o({\u2_Display/add56/c20 ,\u2_Display/n1717 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u2  (
    .a(\u2_Display/n1712 ),
    .b(1'b1),
    .c(\u2_Display/add56/c2 ),
    .o({\u2_Display/add56/c3 ,\u2_Display/n1717 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u20  (
    .a(\u2_Display/n1694 ),
    .b(1'b1),
    .c(\u2_Display/add56/c20 ),
    .o({\u2_Display/add56/c21 ,\u2_Display/n1717 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u21  (
    .a(\u2_Display/n1693 ),
    .b(1'b1),
    .c(\u2_Display/add56/c21 ),
    .o({\u2_Display/add56/c22 ,\u2_Display/n1717 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u22  (
    .a(\u2_Display/n1692 ),
    .b(1'b1),
    .c(\u2_Display/add56/c22 ),
    .o({\u2_Display/add56/c23 ,\u2_Display/n1717 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u23  (
    .a(\u2_Display/n1691 ),
    .b(1'b1),
    .c(\u2_Display/add56/c23 ),
    .o({\u2_Display/add56/c24 ,\u2_Display/n1717 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u24  (
    .a(\u2_Display/n1690 ),
    .b(1'b0),
    .c(\u2_Display/add56/c24 ),
    .o({\u2_Display/add56/c25 ,\u2_Display/n1717 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u25  (
    .a(\u2_Display/n1689 ),
    .b(1'b0),
    .c(\u2_Display/add56/c25 ),
    .o({\u2_Display/add56/c26 ,\u2_Display/n1717 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u26  (
    .a(\u2_Display/n1688 ),
    .b(1'b0),
    .c(\u2_Display/add56/c26 ),
    .o({\u2_Display/add56/c27 ,\u2_Display/n1717 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u27  (
    .a(\u2_Display/n1687 ),
    .b(1'b1),
    .c(\u2_Display/add56/c27 ),
    .o({\u2_Display/add56/c28 ,\u2_Display/n1717 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u28  (
    .a(\u2_Display/n1686 ),
    .b(1'b1),
    .c(\u2_Display/add56/c28 ),
    .o({\u2_Display/add56/c29 ,\u2_Display/n1717 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u29  (
    .a(\u2_Display/n1685 ),
    .b(1'b1),
    .c(\u2_Display/add56/c29 ),
    .o({\u2_Display/add56/c30 ,\u2_Display/n1717 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u3  (
    .a(\u2_Display/n1711 ),
    .b(1'b1),
    .c(\u2_Display/add56/c3 ),
    .o({\u2_Display/add56/c4 ,\u2_Display/n1717 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u30  (
    .a(\u2_Display/n1684 ),
    .b(1'b1),
    .c(\u2_Display/add56/c30 ),
    .o({\u2_Display/add56/c31 ,\u2_Display/n1717 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u31  (
    .a(\u2_Display/n1683 ),
    .b(1'b1),
    .c(\u2_Display/add56/c31 ),
    .o({open_n1215,\u2_Display/n1717 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u4  (
    .a(\u2_Display/n1710 ),
    .b(1'b1),
    .c(\u2_Display/add56/c4 ),
    .o({\u2_Display/add56/c5 ,\u2_Display/n1717 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u5  (
    .a(\u2_Display/n1709 ),
    .b(1'b1),
    .c(\u2_Display/add56/c5 ),
    .o({\u2_Display/add56/c6 ,\u2_Display/n1717 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u6  (
    .a(\u2_Display/n1708 ),
    .b(1'b1),
    .c(\u2_Display/add56/c6 ),
    .o({\u2_Display/add56/c7 ,\u2_Display/n1717 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u7  (
    .a(\u2_Display/n1707 ),
    .b(1'b1),
    .c(\u2_Display/add56/c7 ),
    .o({\u2_Display/add56/c8 ,\u2_Display/n1717 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u8  (
    .a(\u2_Display/n1706 ),
    .b(1'b1),
    .c(\u2_Display/add56/c8 ),
    .o({\u2_Display/add56/c9 ,\u2_Display/n1717 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add56/u9  (
    .a(\u2_Display/n1705 ),
    .b(1'b1),
    .c(\u2_Display/add56/c9 ),
    .o({\u2_Display/add56/c10 ,\u2_Display/n1717 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add56/ucin  (
    .a(1'b1),
    .o({\u2_Display/add56/c0 ,open_n1218}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u0  (
    .a(\u2_Display/n1749 ),
    .b(1'b1),
    .c(\u2_Display/add57/c0 ),
    .o({\u2_Display/add57/c1 ,\u2_Display/n1752 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u1  (
    .a(\u2_Display/n1748 ),
    .b(1'b1),
    .c(\u2_Display/add57/c1 ),
    .o({\u2_Display/add57/c2 ,\u2_Display/n1752 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u10  (
    .a(\u2_Display/n1739 ),
    .b(1'b1),
    .c(\u2_Display/add57/c10 ),
    .o({\u2_Display/add57/c11 ,\u2_Display/n1752 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u11  (
    .a(\u2_Display/n1738 ),
    .b(1'b1),
    .c(\u2_Display/add57/c11 ),
    .o({\u2_Display/add57/c12 ,\u2_Display/n1752 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u12  (
    .a(\u2_Display/n1737 ),
    .b(1'b1),
    .c(\u2_Display/add57/c12 ),
    .o({\u2_Display/add57/c13 ,\u2_Display/n1752 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u13  (
    .a(\u2_Display/n1736 ),
    .b(1'b1),
    .c(\u2_Display/add57/c13 ),
    .o({\u2_Display/add57/c14 ,\u2_Display/n1752 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u14  (
    .a(\u2_Display/n1735 ),
    .b(1'b1),
    .c(\u2_Display/add57/c14 ),
    .o({\u2_Display/add57/c15 ,\u2_Display/n1752 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u15  (
    .a(\u2_Display/n1734 ),
    .b(1'b1),
    .c(\u2_Display/add57/c15 ),
    .o({\u2_Display/add57/c16 ,\u2_Display/n1752 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u16  (
    .a(\u2_Display/n1733 ),
    .b(1'b1),
    .c(\u2_Display/add57/c16 ),
    .o({\u2_Display/add57/c17 ,\u2_Display/n1752 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u17  (
    .a(\u2_Display/n1732 ),
    .b(1'b1),
    .c(\u2_Display/add57/c17 ),
    .o({\u2_Display/add57/c18 ,\u2_Display/n1752 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u18  (
    .a(\u2_Display/n1731 ),
    .b(1'b0),
    .c(\u2_Display/add57/c18 ),
    .o({\u2_Display/add57/c19 ,\u2_Display/n1752 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u19  (
    .a(\u2_Display/n1730 ),
    .b(1'b1),
    .c(\u2_Display/add57/c19 ),
    .o({\u2_Display/add57/c20 ,\u2_Display/n1752 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u2  (
    .a(\u2_Display/n1747 ),
    .b(1'b1),
    .c(\u2_Display/add57/c2 ),
    .o({\u2_Display/add57/c3 ,\u2_Display/n1752 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u20  (
    .a(\u2_Display/n1729 ),
    .b(1'b1),
    .c(\u2_Display/add57/c20 ),
    .o({\u2_Display/add57/c21 ,\u2_Display/n1752 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u21  (
    .a(\u2_Display/n1728 ),
    .b(1'b1),
    .c(\u2_Display/add57/c21 ),
    .o({\u2_Display/add57/c22 ,\u2_Display/n1752 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u22  (
    .a(\u2_Display/n1727 ),
    .b(1'b1),
    .c(\u2_Display/add57/c22 ),
    .o({\u2_Display/add57/c23 ,\u2_Display/n1752 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u23  (
    .a(\u2_Display/n1726 ),
    .b(1'b0),
    .c(\u2_Display/add57/c23 ),
    .o({\u2_Display/add57/c24 ,\u2_Display/n1752 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u24  (
    .a(\u2_Display/n1725 ),
    .b(1'b0),
    .c(\u2_Display/add57/c24 ),
    .o({\u2_Display/add57/c25 ,\u2_Display/n1752 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u25  (
    .a(\u2_Display/n1724 ),
    .b(1'b0),
    .c(\u2_Display/add57/c25 ),
    .o({\u2_Display/add57/c26 ,\u2_Display/n1752 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u26  (
    .a(\u2_Display/n1723 ),
    .b(1'b1),
    .c(\u2_Display/add57/c26 ),
    .o({\u2_Display/add57/c27 ,\u2_Display/n1752 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u27  (
    .a(\u2_Display/n1722 ),
    .b(1'b1),
    .c(\u2_Display/add57/c27 ),
    .o({\u2_Display/add57/c28 ,\u2_Display/n1752 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u28  (
    .a(\u2_Display/n1721 ),
    .b(1'b1),
    .c(\u2_Display/add57/c28 ),
    .o({\u2_Display/add57/c29 ,\u2_Display/n1752 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u29  (
    .a(\u2_Display/n1720 ),
    .b(1'b1),
    .c(\u2_Display/add57/c29 ),
    .o({\u2_Display/add57/c30 ,\u2_Display/n1752 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u3  (
    .a(\u2_Display/n1746 ),
    .b(1'b1),
    .c(\u2_Display/add57/c3 ),
    .o({\u2_Display/add57/c4 ,\u2_Display/n1752 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u30  (
    .a(\u2_Display/n1719 ),
    .b(1'b1),
    .c(\u2_Display/add57/c30 ),
    .o({\u2_Display/add57/c31 ,\u2_Display/n1752 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u31  (
    .a(\u2_Display/n1718 ),
    .b(1'b1),
    .c(\u2_Display/add57/c31 ),
    .o({open_n1219,\u2_Display/n1752 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u4  (
    .a(\u2_Display/n1745 ),
    .b(1'b1),
    .c(\u2_Display/add57/c4 ),
    .o({\u2_Display/add57/c5 ,\u2_Display/n1752 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u5  (
    .a(\u2_Display/n1744 ),
    .b(1'b1),
    .c(\u2_Display/add57/c5 ),
    .o({\u2_Display/add57/c6 ,\u2_Display/n1752 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u6  (
    .a(\u2_Display/n1743 ),
    .b(1'b1),
    .c(\u2_Display/add57/c6 ),
    .o({\u2_Display/add57/c7 ,\u2_Display/n1752 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u7  (
    .a(\u2_Display/n1742 ),
    .b(1'b1),
    .c(\u2_Display/add57/c7 ),
    .o({\u2_Display/add57/c8 ,\u2_Display/n1752 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u8  (
    .a(\u2_Display/n1741 ),
    .b(1'b1),
    .c(\u2_Display/add57/c8 ),
    .o({\u2_Display/add57/c9 ,\u2_Display/n1752 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add57/u9  (
    .a(\u2_Display/n1740 ),
    .b(1'b1),
    .c(\u2_Display/add57/c9 ),
    .o({\u2_Display/add57/c10 ,\u2_Display/n1752 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add57/ucin  (
    .a(1'b1),
    .o({\u2_Display/add57/c0 ,open_n1222}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u0  (
    .a(\u2_Display/n1784 ),
    .b(1'b1),
    .c(\u2_Display/add58/c0 ),
    .o({\u2_Display/add58/c1 ,\u2_Display/n1787 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u1  (
    .a(\u2_Display/n1783 ),
    .b(1'b1),
    .c(\u2_Display/add58/c1 ),
    .o({\u2_Display/add58/c2 ,\u2_Display/n1787 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u10  (
    .a(\u2_Display/n1774 ),
    .b(1'b1),
    .c(\u2_Display/add58/c10 ),
    .o({\u2_Display/add58/c11 ,\u2_Display/n1787 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u11  (
    .a(\u2_Display/n1773 ),
    .b(1'b1),
    .c(\u2_Display/add58/c11 ),
    .o({\u2_Display/add58/c12 ,\u2_Display/n1787 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u12  (
    .a(\u2_Display/n1772 ),
    .b(1'b1),
    .c(\u2_Display/add58/c12 ),
    .o({\u2_Display/add58/c13 ,\u2_Display/n1787 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u13  (
    .a(\u2_Display/n1771 ),
    .b(1'b1),
    .c(\u2_Display/add58/c13 ),
    .o({\u2_Display/add58/c14 ,\u2_Display/n1787 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u14  (
    .a(\u2_Display/n1770 ),
    .b(1'b1),
    .c(\u2_Display/add58/c14 ),
    .o({\u2_Display/add58/c15 ,\u2_Display/n1787 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u15  (
    .a(\u2_Display/n1769 ),
    .b(1'b1),
    .c(\u2_Display/add58/c15 ),
    .o({\u2_Display/add58/c16 ,\u2_Display/n1787 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u16  (
    .a(\u2_Display/n1768 ),
    .b(1'b1),
    .c(\u2_Display/add58/c16 ),
    .o({\u2_Display/add58/c17 ,\u2_Display/n1787 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u17  (
    .a(\u2_Display/n1767 ),
    .b(1'b0),
    .c(\u2_Display/add58/c17 ),
    .o({\u2_Display/add58/c18 ,\u2_Display/n1787 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u18  (
    .a(\u2_Display/n1766 ),
    .b(1'b1),
    .c(\u2_Display/add58/c18 ),
    .o({\u2_Display/add58/c19 ,\u2_Display/n1787 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u19  (
    .a(\u2_Display/n1765 ),
    .b(1'b1),
    .c(\u2_Display/add58/c19 ),
    .o({\u2_Display/add58/c20 ,\u2_Display/n1787 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u2  (
    .a(\u2_Display/n1782 ),
    .b(1'b1),
    .c(\u2_Display/add58/c2 ),
    .o({\u2_Display/add58/c3 ,\u2_Display/n1787 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u20  (
    .a(\u2_Display/n1764 ),
    .b(1'b1),
    .c(\u2_Display/add58/c20 ),
    .o({\u2_Display/add58/c21 ,\u2_Display/n1787 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u21  (
    .a(\u2_Display/n1763 ),
    .b(1'b1),
    .c(\u2_Display/add58/c21 ),
    .o({\u2_Display/add58/c22 ,\u2_Display/n1787 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u22  (
    .a(\u2_Display/n1762 ),
    .b(1'b0),
    .c(\u2_Display/add58/c22 ),
    .o({\u2_Display/add58/c23 ,\u2_Display/n1787 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u23  (
    .a(\u2_Display/n1761 ),
    .b(1'b0),
    .c(\u2_Display/add58/c23 ),
    .o({\u2_Display/add58/c24 ,\u2_Display/n1787 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u24  (
    .a(\u2_Display/n1760 ),
    .b(1'b0),
    .c(\u2_Display/add58/c24 ),
    .o({\u2_Display/add58/c25 ,\u2_Display/n1787 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u25  (
    .a(\u2_Display/n1759 ),
    .b(1'b1),
    .c(\u2_Display/add58/c25 ),
    .o({\u2_Display/add58/c26 ,\u2_Display/n1787 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u26  (
    .a(\u2_Display/n1758 ),
    .b(1'b1),
    .c(\u2_Display/add58/c26 ),
    .o({\u2_Display/add58/c27 ,\u2_Display/n1787 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u27  (
    .a(\u2_Display/n1757 ),
    .b(1'b1),
    .c(\u2_Display/add58/c27 ),
    .o({\u2_Display/add58/c28 ,\u2_Display/n1787 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u28  (
    .a(\u2_Display/n1756 ),
    .b(1'b1),
    .c(\u2_Display/add58/c28 ),
    .o({\u2_Display/add58/c29 ,\u2_Display/n1787 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u29  (
    .a(\u2_Display/n1755 ),
    .b(1'b1),
    .c(\u2_Display/add58/c29 ),
    .o({\u2_Display/add58/c30 ,\u2_Display/n1787 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u3  (
    .a(\u2_Display/n1781 ),
    .b(1'b1),
    .c(\u2_Display/add58/c3 ),
    .o({\u2_Display/add58/c4 ,\u2_Display/n1787 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u30  (
    .a(\u2_Display/n1754 ),
    .b(1'b1),
    .c(\u2_Display/add58/c30 ),
    .o({\u2_Display/add58/c31 ,\u2_Display/n1787 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u31  (
    .a(\u2_Display/n1753 ),
    .b(1'b1),
    .c(\u2_Display/add58/c31 ),
    .o({open_n1223,\u2_Display/n1787 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u4  (
    .a(\u2_Display/n1780 ),
    .b(1'b1),
    .c(\u2_Display/add58/c4 ),
    .o({\u2_Display/add58/c5 ,\u2_Display/n1787 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u5  (
    .a(\u2_Display/n1779 ),
    .b(1'b1),
    .c(\u2_Display/add58/c5 ),
    .o({\u2_Display/add58/c6 ,\u2_Display/n1787 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u6  (
    .a(\u2_Display/n1778 ),
    .b(1'b1),
    .c(\u2_Display/add58/c6 ),
    .o({\u2_Display/add58/c7 ,\u2_Display/n1787 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u7  (
    .a(\u2_Display/n1777 ),
    .b(1'b1),
    .c(\u2_Display/add58/c7 ),
    .o({\u2_Display/add58/c8 ,\u2_Display/n1787 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u8  (
    .a(\u2_Display/n1776 ),
    .b(1'b1),
    .c(\u2_Display/add58/c8 ),
    .o({\u2_Display/add58/c9 ,\u2_Display/n1787 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add58/u9  (
    .a(\u2_Display/n1775 ),
    .b(1'b1),
    .c(\u2_Display/add58/c9 ),
    .o({\u2_Display/add58/c10 ,\u2_Display/n1787 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add58/ucin  (
    .a(1'b1),
    .o({\u2_Display/add58/c0 ,open_n1226}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u0  (
    .a(\u2_Display/n1819 ),
    .b(1'b1),
    .c(\u2_Display/add59/c0 ),
    .o({\u2_Display/add59/c1 ,\u2_Display/n1822 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u1  (
    .a(\u2_Display/n1818 ),
    .b(1'b1),
    .c(\u2_Display/add59/c1 ),
    .o({\u2_Display/add59/c2 ,\u2_Display/n1822 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u10  (
    .a(\u2_Display/n1809 ),
    .b(1'b1),
    .c(\u2_Display/add59/c10 ),
    .o({\u2_Display/add59/c11 ,\u2_Display/n1822 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u11  (
    .a(\u2_Display/n1808 ),
    .b(1'b1),
    .c(\u2_Display/add59/c11 ),
    .o({\u2_Display/add59/c12 ,\u2_Display/n1822 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u12  (
    .a(\u2_Display/n1807 ),
    .b(1'b1),
    .c(\u2_Display/add59/c12 ),
    .o({\u2_Display/add59/c13 ,\u2_Display/n1822 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u13  (
    .a(\u2_Display/n1806 ),
    .b(1'b1),
    .c(\u2_Display/add59/c13 ),
    .o({\u2_Display/add59/c14 ,\u2_Display/n1822 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u14  (
    .a(\u2_Display/n1805 ),
    .b(1'b1),
    .c(\u2_Display/add59/c14 ),
    .o({\u2_Display/add59/c15 ,\u2_Display/n1822 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u15  (
    .a(\u2_Display/n1804 ),
    .b(1'b1),
    .c(\u2_Display/add59/c15 ),
    .o({\u2_Display/add59/c16 ,\u2_Display/n1822 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u16  (
    .a(\u2_Display/n1803 ),
    .b(1'b0),
    .c(\u2_Display/add59/c16 ),
    .o({\u2_Display/add59/c17 ,\u2_Display/n1822 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u17  (
    .a(\u2_Display/n1802 ),
    .b(1'b1),
    .c(\u2_Display/add59/c17 ),
    .o({\u2_Display/add59/c18 ,\u2_Display/n1822 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u18  (
    .a(\u2_Display/n1801 ),
    .b(1'b1),
    .c(\u2_Display/add59/c18 ),
    .o({\u2_Display/add59/c19 ,\u2_Display/n1822 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u19  (
    .a(\u2_Display/n1800 ),
    .b(1'b1),
    .c(\u2_Display/add59/c19 ),
    .o({\u2_Display/add59/c20 ,\u2_Display/n1822 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u2  (
    .a(\u2_Display/n1817 ),
    .b(1'b1),
    .c(\u2_Display/add59/c2 ),
    .o({\u2_Display/add59/c3 ,\u2_Display/n1822 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u20  (
    .a(\u2_Display/n1799 ),
    .b(1'b1),
    .c(\u2_Display/add59/c20 ),
    .o({\u2_Display/add59/c21 ,\u2_Display/n1822 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u21  (
    .a(\u2_Display/n1798 ),
    .b(1'b0),
    .c(\u2_Display/add59/c21 ),
    .o({\u2_Display/add59/c22 ,\u2_Display/n1822 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u22  (
    .a(\u2_Display/n1797 ),
    .b(1'b0),
    .c(\u2_Display/add59/c22 ),
    .o({\u2_Display/add59/c23 ,\u2_Display/n1822 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u23  (
    .a(\u2_Display/n1796 ),
    .b(1'b0),
    .c(\u2_Display/add59/c23 ),
    .o({\u2_Display/add59/c24 ,\u2_Display/n1822 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u24  (
    .a(\u2_Display/n1795 ),
    .b(1'b1),
    .c(\u2_Display/add59/c24 ),
    .o({\u2_Display/add59/c25 ,\u2_Display/n1822 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u25  (
    .a(\u2_Display/n1794 ),
    .b(1'b1),
    .c(\u2_Display/add59/c25 ),
    .o({\u2_Display/add59/c26 ,\u2_Display/n1822 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u26  (
    .a(\u2_Display/n1793 ),
    .b(1'b1),
    .c(\u2_Display/add59/c26 ),
    .o({\u2_Display/add59/c27 ,\u2_Display/n1822 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u27  (
    .a(\u2_Display/n1792 ),
    .b(1'b1),
    .c(\u2_Display/add59/c27 ),
    .o({\u2_Display/add59/c28 ,\u2_Display/n1822 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u28  (
    .a(\u2_Display/n1791 ),
    .b(1'b1),
    .c(\u2_Display/add59/c28 ),
    .o({\u2_Display/add59/c29 ,\u2_Display/n1822 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u29  (
    .a(\u2_Display/n1790 ),
    .b(1'b1),
    .c(\u2_Display/add59/c29 ),
    .o({\u2_Display/add59/c30 ,\u2_Display/n1822 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u3  (
    .a(\u2_Display/n1816 ),
    .b(1'b1),
    .c(\u2_Display/add59/c3 ),
    .o({\u2_Display/add59/c4 ,\u2_Display/n1822 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u30  (
    .a(\u2_Display/n1789 ),
    .b(1'b1),
    .c(\u2_Display/add59/c30 ),
    .o({\u2_Display/add59/c31 ,\u2_Display/n1822 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u31  (
    .a(\u2_Display/n1788 ),
    .b(1'b1),
    .c(\u2_Display/add59/c31 ),
    .o({open_n1227,\u2_Display/n1822 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u4  (
    .a(\u2_Display/n1815 ),
    .b(1'b1),
    .c(\u2_Display/add59/c4 ),
    .o({\u2_Display/add59/c5 ,\u2_Display/n1822 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u5  (
    .a(\u2_Display/n1814 ),
    .b(1'b1),
    .c(\u2_Display/add59/c5 ),
    .o({\u2_Display/add59/c6 ,\u2_Display/n1822 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u6  (
    .a(\u2_Display/n1813 ),
    .b(1'b1),
    .c(\u2_Display/add59/c6 ),
    .o({\u2_Display/add59/c7 ,\u2_Display/n1822 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u7  (
    .a(\u2_Display/n1812 ),
    .b(1'b1),
    .c(\u2_Display/add59/c7 ),
    .o({\u2_Display/add59/c8 ,\u2_Display/n1822 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u8  (
    .a(\u2_Display/n1811 ),
    .b(1'b1),
    .c(\u2_Display/add59/c8 ),
    .o({\u2_Display/add59/c9 ,\u2_Display/n1822 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add59/u9  (
    .a(\u2_Display/n1810 ),
    .b(1'b1),
    .c(\u2_Display/add59/c9 ),
    .o({\u2_Display/add59/c10 ,\u2_Display/n1822 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add59/ucin  (
    .a(1'b1),
    .o({\u2_Display/add59/c0 ,open_n1230}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u0  (
    .a(\u2_Display/n1854 ),
    .b(1'b1),
    .c(\u2_Display/add60/c0 ),
    .o({\u2_Display/add60/c1 ,\u2_Display/n1857 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u1  (
    .a(\u2_Display/n1853 ),
    .b(1'b1),
    .c(\u2_Display/add60/c1 ),
    .o({\u2_Display/add60/c2 ,\u2_Display/n1857 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u10  (
    .a(\u2_Display/n1844 ),
    .b(1'b1),
    .c(\u2_Display/add60/c10 ),
    .o({\u2_Display/add60/c11 ,\u2_Display/n1857 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u11  (
    .a(\u2_Display/n1843 ),
    .b(1'b1),
    .c(\u2_Display/add60/c11 ),
    .o({\u2_Display/add60/c12 ,\u2_Display/n1857 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u12  (
    .a(\u2_Display/n1842 ),
    .b(1'b1),
    .c(\u2_Display/add60/c12 ),
    .o({\u2_Display/add60/c13 ,\u2_Display/n1857 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u13  (
    .a(\u2_Display/n1841 ),
    .b(1'b1),
    .c(\u2_Display/add60/c13 ),
    .o({\u2_Display/add60/c14 ,\u2_Display/n1857 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u14  (
    .a(\u2_Display/n1840 ),
    .b(1'b1),
    .c(\u2_Display/add60/c14 ),
    .o({\u2_Display/add60/c15 ,\u2_Display/n1857 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u15  (
    .a(\u2_Display/n1839 ),
    .b(1'b0),
    .c(\u2_Display/add60/c15 ),
    .o({\u2_Display/add60/c16 ,\u2_Display/n1857 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u16  (
    .a(\u2_Display/n1838 ),
    .b(1'b1),
    .c(\u2_Display/add60/c16 ),
    .o({\u2_Display/add60/c17 ,\u2_Display/n1857 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u17  (
    .a(\u2_Display/n1837 ),
    .b(1'b1),
    .c(\u2_Display/add60/c17 ),
    .o({\u2_Display/add60/c18 ,\u2_Display/n1857 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u18  (
    .a(\u2_Display/n1836 ),
    .b(1'b1),
    .c(\u2_Display/add60/c18 ),
    .o({\u2_Display/add60/c19 ,\u2_Display/n1857 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u19  (
    .a(\u2_Display/n1835 ),
    .b(1'b1),
    .c(\u2_Display/add60/c19 ),
    .o({\u2_Display/add60/c20 ,\u2_Display/n1857 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u2  (
    .a(\u2_Display/n1852 ),
    .b(1'b1),
    .c(\u2_Display/add60/c2 ),
    .o({\u2_Display/add60/c3 ,\u2_Display/n1857 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u20  (
    .a(\u2_Display/n1834 ),
    .b(1'b0),
    .c(\u2_Display/add60/c20 ),
    .o({\u2_Display/add60/c21 ,\u2_Display/n1857 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u21  (
    .a(\u2_Display/n1833 ),
    .b(1'b0),
    .c(\u2_Display/add60/c21 ),
    .o({\u2_Display/add60/c22 ,\u2_Display/n1857 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u22  (
    .a(\u2_Display/n1832 ),
    .b(1'b0),
    .c(\u2_Display/add60/c22 ),
    .o({\u2_Display/add60/c23 ,\u2_Display/n1857 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u23  (
    .a(\u2_Display/n1831 ),
    .b(1'b1),
    .c(\u2_Display/add60/c23 ),
    .o({\u2_Display/add60/c24 ,\u2_Display/n1857 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u24  (
    .a(\u2_Display/n1830 ),
    .b(1'b1),
    .c(\u2_Display/add60/c24 ),
    .o({\u2_Display/add60/c25 ,\u2_Display/n1857 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u25  (
    .a(\u2_Display/n1829 ),
    .b(1'b1),
    .c(\u2_Display/add60/c25 ),
    .o({\u2_Display/add60/c26 ,\u2_Display/n1857 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u26  (
    .a(\u2_Display/n1828 ),
    .b(1'b1),
    .c(\u2_Display/add60/c26 ),
    .o({\u2_Display/add60/c27 ,\u2_Display/n1857 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u27  (
    .a(\u2_Display/n1827 ),
    .b(1'b1),
    .c(\u2_Display/add60/c27 ),
    .o({\u2_Display/add60/c28 ,\u2_Display/n1857 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u28  (
    .a(\u2_Display/n1826 ),
    .b(1'b1),
    .c(\u2_Display/add60/c28 ),
    .o({\u2_Display/add60/c29 ,\u2_Display/n1857 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u29  (
    .a(\u2_Display/n1825 ),
    .b(1'b1),
    .c(\u2_Display/add60/c29 ),
    .o({\u2_Display/add60/c30 ,\u2_Display/n1857 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u3  (
    .a(\u2_Display/n1851 ),
    .b(1'b1),
    .c(\u2_Display/add60/c3 ),
    .o({\u2_Display/add60/c4 ,\u2_Display/n1857 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u30  (
    .a(\u2_Display/n1824 ),
    .b(1'b1),
    .c(\u2_Display/add60/c30 ),
    .o({\u2_Display/add60/c31 ,\u2_Display/n1857 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u31  (
    .a(\u2_Display/n1823 ),
    .b(1'b1),
    .c(\u2_Display/add60/c31 ),
    .o({open_n1231,\u2_Display/n1857 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u4  (
    .a(\u2_Display/n1850 ),
    .b(1'b1),
    .c(\u2_Display/add60/c4 ),
    .o({\u2_Display/add60/c5 ,\u2_Display/n1857 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u5  (
    .a(\u2_Display/n1849 ),
    .b(1'b1),
    .c(\u2_Display/add60/c5 ),
    .o({\u2_Display/add60/c6 ,\u2_Display/n1857 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u6  (
    .a(\u2_Display/n1848 ),
    .b(1'b1),
    .c(\u2_Display/add60/c6 ),
    .o({\u2_Display/add60/c7 ,\u2_Display/n1857 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u7  (
    .a(\u2_Display/n1847 ),
    .b(1'b1),
    .c(\u2_Display/add60/c7 ),
    .o({\u2_Display/add60/c8 ,\u2_Display/n1857 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u8  (
    .a(\u2_Display/n1846 ),
    .b(1'b1),
    .c(\u2_Display/add60/c8 ),
    .o({\u2_Display/add60/c9 ,\u2_Display/n1857 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add60/u9  (
    .a(\u2_Display/n1845 ),
    .b(1'b1),
    .c(\u2_Display/add60/c9 ),
    .o({\u2_Display/add60/c10 ,\u2_Display/n1857 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add60/ucin  (
    .a(1'b1),
    .o({\u2_Display/add60/c0 ,open_n1234}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u0  (
    .a(\u2_Display/n1889 ),
    .b(1'b1),
    .c(\u2_Display/add61/c0 ),
    .o({\u2_Display/add61/c1 ,\u2_Display/n1892 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u1  (
    .a(\u2_Display/n1888 ),
    .b(1'b1),
    .c(\u2_Display/add61/c1 ),
    .o({\u2_Display/add61/c2 ,\u2_Display/n1892 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u10  (
    .a(\u2_Display/n1879 ),
    .b(1'b1),
    .c(\u2_Display/add61/c10 ),
    .o({\u2_Display/add61/c11 ,\u2_Display/n1892 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u11  (
    .a(\u2_Display/n1878 ),
    .b(1'b1),
    .c(\u2_Display/add61/c11 ),
    .o({\u2_Display/add61/c12 ,\u2_Display/n1892 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u12  (
    .a(\u2_Display/n1877 ),
    .b(1'b1),
    .c(\u2_Display/add61/c12 ),
    .o({\u2_Display/add61/c13 ,\u2_Display/n1892 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u13  (
    .a(\u2_Display/n1876 ),
    .b(1'b1),
    .c(\u2_Display/add61/c13 ),
    .o({\u2_Display/add61/c14 ,\u2_Display/n1892 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u14  (
    .a(\u2_Display/n1875 ),
    .b(1'b0),
    .c(\u2_Display/add61/c14 ),
    .o({\u2_Display/add61/c15 ,\u2_Display/n1892 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u15  (
    .a(\u2_Display/n1874 ),
    .b(1'b1),
    .c(\u2_Display/add61/c15 ),
    .o({\u2_Display/add61/c16 ,\u2_Display/n1892 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u16  (
    .a(\u2_Display/n1873 ),
    .b(1'b1),
    .c(\u2_Display/add61/c16 ),
    .o({\u2_Display/add61/c17 ,\u2_Display/n1892 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u17  (
    .a(\u2_Display/n1872 ),
    .b(1'b1),
    .c(\u2_Display/add61/c17 ),
    .o({\u2_Display/add61/c18 ,\u2_Display/n1892 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u18  (
    .a(\u2_Display/n1871 ),
    .b(1'b1),
    .c(\u2_Display/add61/c18 ),
    .o({\u2_Display/add61/c19 ,\u2_Display/n1892 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u19  (
    .a(\u2_Display/n1870 ),
    .b(1'b0),
    .c(\u2_Display/add61/c19 ),
    .o({\u2_Display/add61/c20 ,\u2_Display/n1892 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u2  (
    .a(\u2_Display/n1887 ),
    .b(1'b1),
    .c(\u2_Display/add61/c2 ),
    .o({\u2_Display/add61/c3 ,\u2_Display/n1892 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u20  (
    .a(\u2_Display/n1869 ),
    .b(1'b0),
    .c(\u2_Display/add61/c20 ),
    .o({\u2_Display/add61/c21 ,\u2_Display/n1892 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u21  (
    .a(\u2_Display/n1868 ),
    .b(1'b0),
    .c(\u2_Display/add61/c21 ),
    .o({\u2_Display/add61/c22 ,\u2_Display/n1892 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u22  (
    .a(\u2_Display/n1867 ),
    .b(1'b1),
    .c(\u2_Display/add61/c22 ),
    .o({\u2_Display/add61/c23 ,\u2_Display/n1892 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u23  (
    .a(\u2_Display/n1866 ),
    .b(1'b1),
    .c(\u2_Display/add61/c23 ),
    .o({\u2_Display/add61/c24 ,\u2_Display/n1892 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u24  (
    .a(\u2_Display/n1865 ),
    .b(1'b1),
    .c(\u2_Display/add61/c24 ),
    .o({\u2_Display/add61/c25 ,\u2_Display/n1892 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u25  (
    .a(\u2_Display/n1864 ),
    .b(1'b1),
    .c(\u2_Display/add61/c25 ),
    .o({\u2_Display/add61/c26 ,\u2_Display/n1892 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u26  (
    .a(\u2_Display/n1863 ),
    .b(1'b1),
    .c(\u2_Display/add61/c26 ),
    .o({\u2_Display/add61/c27 ,\u2_Display/n1892 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u27  (
    .a(\u2_Display/n1862 ),
    .b(1'b1),
    .c(\u2_Display/add61/c27 ),
    .o({\u2_Display/add61/c28 ,\u2_Display/n1892 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u28  (
    .a(\u2_Display/n1861 ),
    .b(1'b1),
    .c(\u2_Display/add61/c28 ),
    .o({\u2_Display/add61/c29 ,\u2_Display/n1892 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u29  (
    .a(\u2_Display/n1860 ),
    .b(1'b1),
    .c(\u2_Display/add61/c29 ),
    .o({\u2_Display/add61/c30 ,\u2_Display/n1892 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u3  (
    .a(\u2_Display/n1886 ),
    .b(1'b1),
    .c(\u2_Display/add61/c3 ),
    .o({\u2_Display/add61/c4 ,\u2_Display/n1892 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u30  (
    .a(\u2_Display/n1859 ),
    .b(1'b1),
    .c(\u2_Display/add61/c30 ),
    .o({\u2_Display/add61/c31 ,\u2_Display/n1892 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u31  (
    .a(\u2_Display/n1858 ),
    .b(1'b1),
    .c(\u2_Display/add61/c31 ),
    .o({open_n1235,\u2_Display/n1892 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u4  (
    .a(\u2_Display/n1885 ),
    .b(1'b1),
    .c(\u2_Display/add61/c4 ),
    .o({\u2_Display/add61/c5 ,\u2_Display/n1892 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u5  (
    .a(\u2_Display/n1884 ),
    .b(1'b1),
    .c(\u2_Display/add61/c5 ),
    .o({\u2_Display/add61/c6 ,\u2_Display/n1892 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u6  (
    .a(\u2_Display/n1883 ),
    .b(1'b1),
    .c(\u2_Display/add61/c6 ),
    .o({\u2_Display/add61/c7 ,\u2_Display/n1892 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u7  (
    .a(\u2_Display/n1882 ),
    .b(1'b1),
    .c(\u2_Display/add61/c7 ),
    .o({\u2_Display/add61/c8 ,\u2_Display/n1892 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u8  (
    .a(\u2_Display/n1881 ),
    .b(1'b1),
    .c(\u2_Display/add61/c8 ),
    .o({\u2_Display/add61/c9 ,\u2_Display/n1892 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add61/u9  (
    .a(\u2_Display/n1880 ),
    .b(1'b1),
    .c(\u2_Display/add61/c9 ),
    .o({\u2_Display/add61/c10 ,\u2_Display/n1892 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add61/ucin  (
    .a(1'b1),
    .o({\u2_Display/add61/c0 ,open_n1238}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u0  (
    .a(\u2_Display/n1924 ),
    .b(1'b1),
    .c(\u2_Display/add62/c0 ),
    .o({\u2_Display/add62/c1 ,\u2_Display/n1927 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u1  (
    .a(\u2_Display/n1923 ),
    .b(1'b1),
    .c(\u2_Display/add62/c1 ),
    .o({\u2_Display/add62/c2 ,\u2_Display/n1927 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u10  (
    .a(\u2_Display/n1914 ),
    .b(1'b1),
    .c(\u2_Display/add62/c10 ),
    .o({\u2_Display/add62/c11 ,\u2_Display/n1927 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u11  (
    .a(\u2_Display/n1913 ),
    .b(1'b1),
    .c(\u2_Display/add62/c11 ),
    .o({\u2_Display/add62/c12 ,\u2_Display/n1927 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u12  (
    .a(\u2_Display/n1912 ),
    .b(1'b1),
    .c(\u2_Display/add62/c12 ),
    .o({\u2_Display/add62/c13 ,\u2_Display/n1927 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u13  (
    .a(\u2_Display/n1911 ),
    .b(1'b0),
    .c(\u2_Display/add62/c13 ),
    .o({\u2_Display/add62/c14 ,\u2_Display/n1927 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u14  (
    .a(\u2_Display/n1910 ),
    .b(1'b1),
    .c(\u2_Display/add62/c14 ),
    .o({\u2_Display/add62/c15 ,\u2_Display/n1927 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u15  (
    .a(\u2_Display/n1909 ),
    .b(1'b1),
    .c(\u2_Display/add62/c15 ),
    .o({\u2_Display/add62/c16 ,\u2_Display/n1927 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u16  (
    .a(\u2_Display/n1908 ),
    .b(1'b1),
    .c(\u2_Display/add62/c16 ),
    .o({\u2_Display/add62/c17 ,\u2_Display/n1927 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u17  (
    .a(\u2_Display/n1907 ),
    .b(1'b1),
    .c(\u2_Display/add62/c17 ),
    .o({\u2_Display/add62/c18 ,\u2_Display/n1927 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u18  (
    .a(\u2_Display/n1906 ),
    .b(1'b0),
    .c(\u2_Display/add62/c18 ),
    .o({\u2_Display/add62/c19 ,\u2_Display/n1927 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u19  (
    .a(\u2_Display/n1905 ),
    .b(1'b0),
    .c(\u2_Display/add62/c19 ),
    .o({\u2_Display/add62/c20 ,\u2_Display/n1927 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u2  (
    .a(\u2_Display/n1922 ),
    .b(1'b1),
    .c(\u2_Display/add62/c2 ),
    .o({\u2_Display/add62/c3 ,\u2_Display/n1927 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u20  (
    .a(\u2_Display/n1904 ),
    .b(1'b0),
    .c(\u2_Display/add62/c20 ),
    .o({\u2_Display/add62/c21 ,\u2_Display/n1927 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u21  (
    .a(\u2_Display/n1903 ),
    .b(1'b1),
    .c(\u2_Display/add62/c21 ),
    .o({\u2_Display/add62/c22 ,\u2_Display/n1927 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u22  (
    .a(\u2_Display/n1902 ),
    .b(1'b1),
    .c(\u2_Display/add62/c22 ),
    .o({\u2_Display/add62/c23 ,\u2_Display/n1927 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u23  (
    .a(\u2_Display/n1901 ),
    .b(1'b1),
    .c(\u2_Display/add62/c23 ),
    .o({\u2_Display/add62/c24 ,\u2_Display/n1927 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u24  (
    .a(\u2_Display/n1900 ),
    .b(1'b1),
    .c(\u2_Display/add62/c24 ),
    .o({\u2_Display/add62/c25 ,\u2_Display/n1927 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u25  (
    .a(\u2_Display/n1899 ),
    .b(1'b1),
    .c(\u2_Display/add62/c25 ),
    .o({\u2_Display/add62/c26 ,\u2_Display/n1927 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u26  (
    .a(\u2_Display/n1898 ),
    .b(1'b1),
    .c(\u2_Display/add62/c26 ),
    .o({\u2_Display/add62/c27 ,\u2_Display/n1927 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u27  (
    .a(\u2_Display/n1897 ),
    .b(1'b1),
    .c(\u2_Display/add62/c27 ),
    .o({\u2_Display/add62/c28 ,\u2_Display/n1927 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u28  (
    .a(\u2_Display/n1896 ),
    .b(1'b1),
    .c(\u2_Display/add62/c28 ),
    .o({\u2_Display/add62/c29 ,\u2_Display/n1927 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u29  (
    .a(\u2_Display/n1895 ),
    .b(1'b1),
    .c(\u2_Display/add62/c29 ),
    .o({\u2_Display/add62/c30 ,\u2_Display/n1927 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u3  (
    .a(\u2_Display/n1921 ),
    .b(1'b1),
    .c(\u2_Display/add62/c3 ),
    .o({\u2_Display/add62/c4 ,\u2_Display/n1927 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u30  (
    .a(\u2_Display/n1894 ),
    .b(1'b1),
    .c(\u2_Display/add62/c30 ),
    .o({\u2_Display/add62/c31 ,\u2_Display/n1927 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u31  (
    .a(\u2_Display/n1893 ),
    .b(1'b1),
    .c(\u2_Display/add62/c31 ),
    .o({open_n1239,\u2_Display/n1927 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u4  (
    .a(\u2_Display/n1920 ),
    .b(1'b1),
    .c(\u2_Display/add62/c4 ),
    .o({\u2_Display/add62/c5 ,\u2_Display/n1927 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u5  (
    .a(\u2_Display/n1919 ),
    .b(1'b1),
    .c(\u2_Display/add62/c5 ),
    .o({\u2_Display/add62/c6 ,\u2_Display/n1927 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u6  (
    .a(\u2_Display/n1918 ),
    .b(1'b1),
    .c(\u2_Display/add62/c6 ),
    .o({\u2_Display/add62/c7 ,\u2_Display/n1927 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u7  (
    .a(\u2_Display/n1917 ),
    .b(1'b1),
    .c(\u2_Display/add62/c7 ),
    .o({\u2_Display/add62/c8 ,\u2_Display/n1927 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u8  (
    .a(\u2_Display/n1916 ),
    .b(1'b1),
    .c(\u2_Display/add62/c8 ),
    .o({\u2_Display/add62/c9 ,\u2_Display/n1927 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add62/u9  (
    .a(\u2_Display/n1915 ),
    .b(1'b1),
    .c(\u2_Display/add62/c9 ),
    .o({\u2_Display/add62/c10 ,\u2_Display/n1927 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add62/ucin  (
    .a(1'b1),
    .o({\u2_Display/add62/c0 ,open_n1242}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u0  (
    .a(\u2_Display/n1959 ),
    .b(1'b1),
    .c(\u2_Display/add63/c0 ),
    .o({\u2_Display/add63/c1 ,\u2_Display/n1962 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u1  (
    .a(\u2_Display/n1958 ),
    .b(1'b1),
    .c(\u2_Display/add63/c1 ),
    .o({\u2_Display/add63/c2 ,\u2_Display/n1962 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u10  (
    .a(\u2_Display/n1949 ),
    .b(1'b1),
    .c(\u2_Display/add63/c10 ),
    .o({\u2_Display/add63/c11 ,\u2_Display/n1962 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u11  (
    .a(\u2_Display/n1948 ),
    .b(1'b1),
    .c(\u2_Display/add63/c11 ),
    .o({\u2_Display/add63/c12 ,\u2_Display/n1962 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u12  (
    .a(\u2_Display/n1947 ),
    .b(1'b0),
    .c(\u2_Display/add63/c12 ),
    .o({\u2_Display/add63/c13 ,\u2_Display/n1962 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u13  (
    .a(\u2_Display/n1946 ),
    .b(1'b1),
    .c(\u2_Display/add63/c13 ),
    .o({\u2_Display/add63/c14 ,\u2_Display/n1962 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u14  (
    .a(\u2_Display/n1945 ),
    .b(1'b1),
    .c(\u2_Display/add63/c14 ),
    .o({\u2_Display/add63/c15 ,\u2_Display/n1962 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u15  (
    .a(\u2_Display/n1944 ),
    .b(1'b1),
    .c(\u2_Display/add63/c15 ),
    .o({\u2_Display/add63/c16 ,\u2_Display/n1962 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u16  (
    .a(\u2_Display/n1943 ),
    .b(1'b1),
    .c(\u2_Display/add63/c16 ),
    .o({\u2_Display/add63/c17 ,\u2_Display/n1962 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u17  (
    .a(\u2_Display/n1942 ),
    .b(1'b0),
    .c(\u2_Display/add63/c17 ),
    .o({\u2_Display/add63/c18 ,\u2_Display/n1962 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u18  (
    .a(\u2_Display/n1941 ),
    .b(1'b0),
    .c(\u2_Display/add63/c18 ),
    .o({\u2_Display/add63/c19 ,\u2_Display/n1962 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u19  (
    .a(\u2_Display/n1940 ),
    .b(1'b0),
    .c(\u2_Display/add63/c19 ),
    .o({\u2_Display/add63/c20 ,\u2_Display/n1962 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u2  (
    .a(\u2_Display/n1957 ),
    .b(1'b1),
    .c(\u2_Display/add63/c2 ),
    .o({\u2_Display/add63/c3 ,\u2_Display/n1962 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u20  (
    .a(\u2_Display/n1939 ),
    .b(1'b1),
    .c(\u2_Display/add63/c20 ),
    .o({\u2_Display/add63/c21 ,\u2_Display/n1962 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u21  (
    .a(\u2_Display/n1938 ),
    .b(1'b1),
    .c(\u2_Display/add63/c21 ),
    .o({\u2_Display/add63/c22 ,\u2_Display/n1962 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u22  (
    .a(\u2_Display/n1937 ),
    .b(1'b1),
    .c(\u2_Display/add63/c22 ),
    .o({\u2_Display/add63/c23 ,\u2_Display/n1962 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u23  (
    .a(\u2_Display/n1936 ),
    .b(1'b1),
    .c(\u2_Display/add63/c23 ),
    .o({\u2_Display/add63/c24 ,\u2_Display/n1962 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u24  (
    .a(\u2_Display/n1935 ),
    .b(1'b1),
    .c(\u2_Display/add63/c24 ),
    .o({\u2_Display/add63/c25 ,\u2_Display/n1962 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u25  (
    .a(\u2_Display/n1934 ),
    .b(1'b1),
    .c(\u2_Display/add63/c25 ),
    .o({\u2_Display/add63/c26 ,\u2_Display/n1962 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u26  (
    .a(\u2_Display/n1933 ),
    .b(1'b1),
    .c(\u2_Display/add63/c26 ),
    .o({\u2_Display/add63/c27 ,\u2_Display/n1962 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u27  (
    .a(\u2_Display/n1932 ),
    .b(1'b1),
    .c(\u2_Display/add63/c27 ),
    .o({\u2_Display/add63/c28 ,\u2_Display/n1962 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u28  (
    .a(\u2_Display/n1931 ),
    .b(1'b1),
    .c(\u2_Display/add63/c28 ),
    .o({\u2_Display/add63/c29 ,\u2_Display/n1962 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u29  (
    .a(\u2_Display/n1930 ),
    .b(1'b1),
    .c(\u2_Display/add63/c29 ),
    .o({\u2_Display/add63/c30 ,\u2_Display/n1962 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u3  (
    .a(\u2_Display/n1956 ),
    .b(1'b1),
    .c(\u2_Display/add63/c3 ),
    .o({\u2_Display/add63/c4 ,\u2_Display/n1962 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u30  (
    .a(\u2_Display/n1929 ),
    .b(1'b1),
    .c(\u2_Display/add63/c30 ),
    .o({\u2_Display/add63/c31 ,\u2_Display/n1962 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u31  (
    .a(\u2_Display/n1928 ),
    .b(1'b1),
    .c(\u2_Display/add63/c31 ),
    .o({open_n1243,\u2_Display/n1962 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u4  (
    .a(\u2_Display/n1955 ),
    .b(1'b1),
    .c(\u2_Display/add63/c4 ),
    .o({\u2_Display/add63/c5 ,\u2_Display/n1962 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u5  (
    .a(\u2_Display/n1954 ),
    .b(1'b1),
    .c(\u2_Display/add63/c5 ),
    .o({\u2_Display/add63/c6 ,\u2_Display/n1962 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u6  (
    .a(\u2_Display/n1953 ),
    .b(1'b1),
    .c(\u2_Display/add63/c6 ),
    .o({\u2_Display/add63/c7 ,\u2_Display/n1962 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u7  (
    .a(\u2_Display/n1952 ),
    .b(1'b1),
    .c(\u2_Display/add63/c7 ),
    .o({\u2_Display/add63/c8 ,\u2_Display/n1962 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u8  (
    .a(\u2_Display/n1951 ),
    .b(1'b1),
    .c(\u2_Display/add63/c8 ),
    .o({\u2_Display/add63/c9 ,\u2_Display/n1962 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add63/u9  (
    .a(\u2_Display/n1950 ),
    .b(1'b1),
    .c(\u2_Display/add63/c9 ),
    .o({\u2_Display/add63/c10 ,\u2_Display/n1962 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add63/ucin  (
    .a(1'b1),
    .o({\u2_Display/add63/c0 ,open_n1246}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u0  (
    .a(\u2_Display/n1994 ),
    .b(1'b1),
    .c(\u2_Display/add64/c0 ),
    .o({\u2_Display/add64/c1 ,\u2_Display/n1997 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u1  (
    .a(\u2_Display/n1993 ),
    .b(1'b1),
    .c(\u2_Display/add64/c1 ),
    .o({\u2_Display/add64/c2 ,\u2_Display/n1997 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u10  (
    .a(\u2_Display/n1984 ),
    .b(1'b1),
    .c(\u2_Display/add64/c10 ),
    .o({\u2_Display/add64/c11 ,\u2_Display/n1997 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u11  (
    .a(\u2_Display/n1983 ),
    .b(1'b0),
    .c(\u2_Display/add64/c11 ),
    .o({\u2_Display/add64/c12 ,\u2_Display/n1997 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u12  (
    .a(\u2_Display/n1982 ),
    .b(1'b1),
    .c(\u2_Display/add64/c12 ),
    .o({\u2_Display/add64/c13 ,\u2_Display/n1997 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u13  (
    .a(\u2_Display/n1981 ),
    .b(1'b1),
    .c(\u2_Display/add64/c13 ),
    .o({\u2_Display/add64/c14 ,\u2_Display/n1997 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u14  (
    .a(\u2_Display/n1980 ),
    .b(1'b1),
    .c(\u2_Display/add64/c14 ),
    .o({\u2_Display/add64/c15 ,\u2_Display/n1997 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u15  (
    .a(\u2_Display/n1979 ),
    .b(1'b1),
    .c(\u2_Display/add64/c15 ),
    .o({\u2_Display/add64/c16 ,\u2_Display/n1997 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u16  (
    .a(\u2_Display/n1978 ),
    .b(1'b0),
    .c(\u2_Display/add64/c16 ),
    .o({\u2_Display/add64/c17 ,\u2_Display/n1997 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u17  (
    .a(\u2_Display/n1977 ),
    .b(1'b0),
    .c(\u2_Display/add64/c17 ),
    .o({\u2_Display/add64/c18 ,\u2_Display/n1997 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u18  (
    .a(\u2_Display/n1976 ),
    .b(1'b0),
    .c(\u2_Display/add64/c18 ),
    .o({\u2_Display/add64/c19 ,\u2_Display/n1997 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u19  (
    .a(\u2_Display/n1975 ),
    .b(1'b1),
    .c(\u2_Display/add64/c19 ),
    .o({\u2_Display/add64/c20 ,\u2_Display/n1997 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u2  (
    .a(\u2_Display/n1992 ),
    .b(1'b1),
    .c(\u2_Display/add64/c2 ),
    .o({\u2_Display/add64/c3 ,\u2_Display/n1997 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u20  (
    .a(\u2_Display/n1974 ),
    .b(1'b1),
    .c(\u2_Display/add64/c20 ),
    .o({\u2_Display/add64/c21 ,\u2_Display/n1997 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u21  (
    .a(\u2_Display/n1973 ),
    .b(1'b1),
    .c(\u2_Display/add64/c21 ),
    .o({\u2_Display/add64/c22 ,\u2_Display/n1997 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u22  (
    .a(\u2_Display/n1972 ),
    .b(1'b1),
    .c(\u2_Display/add64/c22 ),
    .o({\u2_Display/add64/c23 ,\u2_Display/n1997 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u23  (
    .a(\u2_Display/n1971 ),
    .b(1'b1),
    .c(\u2_Display/add64/c23 ),
    .o({\u2_Display/add64/c24 ,\u2_Display/n1997 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u24  (
    .a(\u2_Display/n1970 ),
    .b(1'b1),
    .c(\u2_Display/add64/c24 ),
    .o({\u2_Display/add64/c25 ,\u2_Display/n1997 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u25  (
    .a(\u2_Display/n1969 ),
    .b(1'b1),
    .c(\u2_Display/add64/c25 ),
    .o({\u2_Display/add64/c26 ,\u2_Display/n1997 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u26  (
    .a(\u2_Display/n1968 ),
    .b(1'b1),
    .c(\u2_Display/add64/c26 ),
    .o({\u2_Display/add64/c27 ,\u2_Display/n1997 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u27  (
    .a(\u2_Display/n1967 ),
    .b(1'b1),
    .c(\u2_Display/add64/c27 ),
    .o({\u2_Display/add64/c28 ,\u2_Display/n1997 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u28  (
    .a(\u2_Display/n1966 ),
    .b(1'b1),
    .c(\u2_Display/add64/c28 ),
    .o({\u2_Display/add64/c29 ,\u2_Display/n1997 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u29  (
    .a(\u2_Display/n1965 ),
    .b(1'b1),
    .c(\u2_Display/add64/c29 ),
    .o({\u2_Display/add64/c30 ,\u2_Display/n1997 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u3  (
    .a(\u2_Display/n1991 ),
    .b(1'b1),
    .c(\u2_Display/add64/c3 ),
    .o({\u2_Display/add64/c4 ,\u2_Display/n1997 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u30  (
    .a(\u2_Display/n1964 ),
    .b(1'b1),
    .c(\u2_Display/add64/c30 ),
    .o({\u2_Display/add64/c31 ,\u2_Display/n1997 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u31  (
    .a(\u2_Display/n1963 ),
    .b(1'b1),
    .c(\u2_Display/add64/c31 ),
    .o({open_n1247,\u2_Display/n1997 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u4  (
    .a(\u2_Display/n1990 ),
    .b(1'b1),
    .c(\u2_Display/add64/c4 ),
    .o({\u2_Display/add64/c5 ,\u2_Display/n1997 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u5  (
    .a(\u2_Display/n1989 ),
    .b(1'b1),
    .c(\u2_Display/add64/c5 ),
    .o({\u2_Display/add64/c6 ,\u2_Display/n1997 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u6  (
    .a(\u2_Display/n1988 ),
    .b(1'b1),
    .c(\u2_Display/add64/c6 ),
    .o({\u2_Display/add64/c7 ,\u2_Display/n1997 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u7  (
    .a(\u2_Display/n1987 ),
    .b(1'b1),
    .c(\u2_Display/add64/c7 ),
    .o({\u2_Display/add64/c8 ,\u2_Display/n1997 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u8  (
    .a(\u2_Display/n1986 ),
    .b(1'b1),
    .c(\u2_Display/add64/c8 ),
    .o({\u2_Display/add64/c9 ,\u2_Display/n1997 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add64/u9  (
    .a(\u2_Display/n1985 ),
    .b(1'b1),
    .c(\u2_Display/add64/c9 ),
    .o({\u2_Display/add64/c10 ,\u2_Display/n1997 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add64/ucin  (
    .a(1'b1),
    .o({\u2_Display/add64/c0 ,open_n1250}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u0  (
    .a(\u2_Display/n2029 ),
    .b(1'b1),
    .c(\u2_Display/add65/c0 ),
    .o({\u2_Display/add65/c1 ,\u2_Display/n2032 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u1  (
    .a(\u2_Display/n2028 ),
    .b(1'b1),
    .c(\u2_Display/add65/c1 ),
    .o({\u2_Display/add65/c2 ,\u2_Display/n2032 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u10  (
    .a(\u2_Display/n2019 ),
    .b(1'b0),
    .c(\u2_Display/add65/c10 ),
    .o({\u2_Display/add65/c11 ,\u2_Display/n2032 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u11  (
    .a(\u2_Display/n2018 ),
    .b(1'b1),
    .c(\u2_Display/add65/c11 ),
    .o({\u2_Display/add65/c12 ,\u2_Display/n2032 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u12  (
    .a(\u2_Display/n2017 ),
    .b(1'b1),
    .c(\u2_Display/add65/c12 ),
    .o({\u2_Display/add65/c13 ,\u2_Display/n2032 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u13  (
    .a(\u2_Display/n2016 ),
    .b(1'b1),
    .c(\u2_Display/add65/c13 ),
    .o({\u2_Display/add65/c14 ,\u2_Display/n2032 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u14  (
    .a(\u2_Display/n2015 ),
    .b(1'b1),
    .c(\u2_Display/add65/c14 ),
    .o({\u2_Display/add65/c15 ,\u2_Display/n2032 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u15  (
    .a(\u2_Display/n2014 ),
    .b(1'b0),
    .c(\u2_Display/add65/c15 ),
    .o({\u2_Display/add65/c16 ,\u2_Display/n2032 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u16  (
    .a(\u2_Display/n2013 ),
    .b(1'b0),
    .c(\u2_Display/add65/c16 ),
    .o({\u2_Display/add65/c17 ,\u2_Display/n2032 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u17  (
    .a(\u2_Display/n2012 ),
    .b(1'b0),
    .c(\u2_Display/add65/c17 ),
    .o({\u2_Display/add65/c18 ,\u2_Display/n2032 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u18  (
    .a(\u2_Display/n2011 ),
    .b(1'b1),
    .c(\u2_Display/add65/c18 ),
    .o({\u2_Display/add65/c19 ,\u2_Display/n2032 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u19  (
    .a(\u2_Display/n2010 ),
    .b(1'b1),
    .c(\u2_Display/add65/c19 ),
    .o({\u2_Display/add65/c20 ,\u2_Display/n2032 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u2  (
    .a(\u2_Display/n2027 ),
    .b(1'b1),
    .c(\u2_Display/add65/c2 ),
    .o({\u2_Display/add65/c3 ,\u2_Display/n2032 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u20  (
    .a(\u2_Display/n2009 ),
    .b(1'b1),
    .c(\u2_Display/add65/c20 ),
    .o({\u2_Display/add65/c21 ,\u2_Display/n2032 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u21  (
    .a(\u2_Display/n2008 ),
    .b(1'b1),
    .c(\u2_Display/add65/c21 ),
    .o({\u2_Display/add65/c22 ,\u2_Display/n2032 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u22  (
    .a(\u2_Display/n2007 ),
    .b(1'b1),
    .c(\u2_Display/add65/c22 ),
    .o({\u2_Display/add65/c23 ,\u2_Display/n2032 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u23  (
    .a(\u2_Display/n2006 ),
    .b(1'b1),
    .c(\u2_Display/add65/c23 ),
    .o({\u2_Display/add65/c24 ,\u2_Display/n2032 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u24  (
    .a(\u2_Display/n2005 ),
    .b(1'b1),
    .c(\u2_Display/add65/c24 ),
    .o({\u2_Display/add65/c25 ,\u2_Display/n2032 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u25  (
    .a(\u2_Display/n2004 ),
    .b(1'b1),
    .c(\u2_Display/add65/c25 ),
    .o({\u2_Display/add65/c26 ,\u2_Display/n2032 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u26  (
    .a(\u2_Display/n2003 ),
    .b(1'b1),
    .c(\u2_Display/add65/c26 ),
    .o({\u2_Display/add65/c27 ,\u2_Display/n2032 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u27  (
    .a(\u2_Display/n2002 ),
    .b(1'b1),
    .c(\u2_Display/add65/c27 ),
    .o({\u2_Display/add65/c28 ,\u2_Display/n2032 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u28  (
    .a(\u2_Display/n2001 ),
    .b(1'b1),
    .c(\u2_Display/add65/c28 ),
    .o({\u2_Display/add65/c29 ,\u2_Display/n2032 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u29  (
    .a(\u2_Display/n2000 ),
    .b(1'b1),
    .c(\u2_Display/add65/c29 ),
    .o({\u2_Display/add65/c30 ,\u2_Display/n2032 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u3  (
    .a(\u2_Display/n2026 ),
    .b(1'b1),
    .c(\u2_Display/add65/c3 ),
    .o({\u2_Display/add65/c4 ,\u2_Display/n2032 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u30  (
    .a(\u2_Display/n1999 ),
    .b(1'b1),
    .c(\u2_Display/add65/c30 ),
    .o({\u2_Display/add65/c31 ,\u2_Display/n2032 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u31  (
    .a(\u2_Display/n1998 ),
    .b(1'b1),
    .c(\u2_Display/add65/c31 ),
    .o({open_n1251,\u2_Display/n2032 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u4  (
    .a(\u2_Display/n2025 ),
    .b(1'b1),
    .c(\u2_Display/add65/c4 ),
    .o({\u2_Display/add65/c5 ,\u2_Display/n2032 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u5  (
    .a(\u2_Display/n2024 ),
    .b(1'b1),
    .c(\u2_Display/add65/c5 ),
    .o({\u2_Display/add65/c6 ,\u2_Display/n2032 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u6  (
    .a(\u2_Display/n2023 ),
    .b(1'b1),
    .c(\u2_Display/add65/c6 ),
    .o({\u2_Display/add65/c7 ,\u2_Display/n2032 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u7  (
    .a(\u2_Display/n2022 ),
    .b(1'b1),
    .c(\u2_Display/add65/c7 ),
    .o({\u2_Display/add65/c8 ,\u2_Display/n2032 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u8  (
    .a(\u2_Display/n2021 ),
    .b(1'b1),
    .c(\u2_Display/add65/c8 ),
    .o({\u2_Display/add65/c9 ,\u2_Display/n2032 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add65/u9  (
    .a(\u2_Display/n2020 ),
    .b(1'b1),
    .c(\u2_Display/add65/c9 ),
    .o({\u2_Display/add65/c10 ,\u2_Display/n2032 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add65/ucin  (
    .a(1'b1),
    .o({\u2_Display/add65/c0 ,open_n1254}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u0  (
    .a(\u2_Display/n2064 ),
    .b(1'b1),
    .c(\u2_Display/add66/c0 ),
    .o({\u2_Display/add66/c1 ,\u2_Display/n2067 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u1  (
    .a(\u2_Display/n2063 ),
    .b(1'b1),
    .c(\u2_Display/add66/c1 ),
    .o({\u2_Display/add66/c2 ,\u2_Display/n2067 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u10  (
    .a(\u2_Display/n2054 ),
    .b(1'b1),
    .c(\u2_Display/add66/c10 ),
    .o({\u2_Display/add66/c11 ,\u2_Display/n2067 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u11  (
    .a(\u2_Display/n2053 ),
    .b(1'b1),
    .c(\u2_Display/add66/c11 ),
    .o({\u2_Display/add66/c12 ,\u2_Display/n2067 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u12  (
    .a(\u2_Display/n2052 ),
    .b(1'b1),
    .c(\u2_Display/add66/c12 ),
    .o({\u2_Display/add66/c13 ,\u2_Display/n2067 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u13  (
    .a(\u2_Display/n2051 ),
    .b(1'b1),
    .c(\u2_Display/add66/c13 ),
    .o({\u2_Display/add66/c14 ,\u2_Display/n2067 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u14  (
    .a(\u2_Display/n2050 ),
    .b(1'b0),
    .c(\u2_Display/add66/c14 ),
    .o({\u2_Display/add66/c15 ,\u2_Display/n2067 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u15  (
    .a(\u2_Display/n2049 ),
    .b(1'b0),
    .c(\u2_Display/add66/c15 ),
    .o({\u2_Display/add66/c16 ,\u2_Display/n2067 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u16  (
    .a(\u2_Display/n2048 ),
    .b(1'b0),
    .c(\u2_Display/add66/c16 ),
    .o({\u2_Display/add66/c17 ,\u2_Display/n2067 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u17  (
    .a(\u2_Display/n2047 ),
    .b(1'b1),
    .c(\u2_Display/add66/c17 ),
    .o({\u2_Display/add66/c18 ,\u2_Display/n2067 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u18  (
    .a(\u2_Display/n2046 ),
    .b(1'b1),
    .c(\u2_Display/add66/c18 ),
    .o({\u2_Display/add66/c19 ,\u2_Display/n2067 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u19  (
    .a(\u2_Display/n2045 ),
    .b(1'b1),
    .c(\u2_Display/add66/c19 ),
    .o({\u2_Display/add66/c20 ,\u2_Display/n2067 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u2  (
    .a(\u2_Display/n2062 ),
    .b(1'b1),
    .c(\u2_Display/add66/c2 ),
    .o({\u2_Display/add66/c3 ,\u2_Display/n2067 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u20  (
    .a(\u2_Display/n2044 ),
    .b(1'b1),
    .c(\u2_Display/add66/c20 ),
    .o({\u2_Display/add66/c21 ,\u2_Display/n2067 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u21  (
    .a(\u2_Display/n2043 ),
    .b(1'b1),
    .c(\u2_Display/add66/c21 ),
    .o({\u2_Display/add66/c22 ,\u2_Display/n2067 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u22  (
    .a(\u2_Display/n2042 ),
    .b(1'b1),
    .c(\u2_Display/add66/c22 ),
    .o({\u2_Display/add66/c23 ,\u2_Display/n2067 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u23  (
    .a(\u2_Display/n2041 ),
    .b(1'b1),
    .c(\u2_Display/add66/c23 ),
    .o({\u2_Display/add66/c24 ,\u2_Display/n2067 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u24  (
    .a(\u2_Display/n2040 ),
    .b(1'b1),
    .c(\u2_Display/add66/c24 ),
    .o({\u2_Display/add66/c25 ,\u2_Display/n2067 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u25  (
    .a(\u2_Display/n2039 ),
    .b(1'b1),
    .c(\u2_Display/add66/c25 ),
    .o({\u2_Display/add66/c26 ,\u2_Display/n2067 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u26  (
    .a(\u2_Display/n2038 ),
    .b(1'b1),
    .c(\u2_Display/add66/c26 ),
    .o({\u2_Display/add66/c27 ,\u2_Display/n2067 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u27  (
    .a(\u2_Display/n2037 ),
    .b(1'b1),
    .c(\u2_Display/add66/c27 ),
    .o({\u2_Display/add66/c28 ,\u2_Display/n2067 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u28  (
    .a(\u2_Display/n2036 ),
    .b(1'b1),
    .c(\u2_Display/add66/c28 ),
    .o({\u2_Display/add66/c29 ,\u2_Display/n2067 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u29  (
    .a(\u2_Display/n2035 ),
    .b(1'b1),
    .c(\u2_Display/add66/c29 ),
    .o({\u2_Display/add66/c30 ,\u2_Display/n2067 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u3  (
    .a(\u2_Display/n2061 ),
    .b(1'b1),
    .c(\u2_Display/add66/c3 ),
    .o({\u2_Display/add66/c4 ,\u2_Display/n2067 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u30  (
    .a(\u2_Display/n2034 ),
    .b(1'b1),
    .c(\u2_Display/add66/c30 ),
    .o({\u2_Display/add66/c31 ,\u2_Display/n2067 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u31  (
    .a(\u2_Display/n2033 ),
    .b(1'b1),
    .c(\u2_Display/add66/c31 ),
    .o({open_n1255,\u2_Display/n2067 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u4  (
    .a(\u2_Display/n2060 ),
    .b(1'b1),
    .c(\u2_Display/add66/c4 ),
    .o({\u2_Display/add66/c5 ,\u2_Display/n2067 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u5  (
    .a(\u2_Display/n2059 ),
    .b(1'b1),
    .c(\u2_Display/add66/c5 ),
    .o({\u2_Display/add66/c6 ,\u2_Display/n2067 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u6  (
    .a(\u2_Display/n2058 ),
    .b(1'b1),
    .c(\u2_Display/add66/c6 ),
    .o({\u2_Display/add66/c7 ,\u2_Display/n2067 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u7  (
    .a(\u2_Display/n2057 ),
    .b(1'b1),
    .c(\u2_Display/add66/c7 ),
    .o({\u2_Display/add66/c8 ,\u2_Display/n2067 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u8  (
    .a(\u2_Display/n2056 ),
    .b(1'b1),
    .c(\u2_Display/add66/c8 ),
    .o({\u2_Display/add66/c9 ,\u2_Display/n2067 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add66/u9  (
    .a(\u2_Display/n2055 ),
    .b(1'b0),
    .c(\u2_Display/add66/c9 ),
    .o({\u2_Display/add66/c10 ,\u2_Display/n2067 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add66/ucin  (
    .a(1'b1),
    .o({\u2_Display/add66/c0 ,open_n1258}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u0  (
    .a(\u2_Display/n2099 ),
    .b(1'b1),
    .c(\u2_Display/add67/c0 ),
    .o({\u2_Display/add67/c1 ,\u2_Display/n2102 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u1  (
    .a(\u2_Display/n2098 ),
    .b(1'b1),
    .c(\u2_Display/add67/c1 ),
    .o({\u2_Display/add67/c2 ,\u2_Display/n2102 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u10  (
    .a(\u2_Display/n2089 ),
    .b(1'b1),
    .c(\u2_Display/add67/c10 ),
    .o({\u2_Display/add67/c11 ,\u2_Display/n2102 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u11  (
    .a(\u2_Display/n2088 ),
    .b(1'b1),
    .c(\u2_Display/add67/c11 ),
    .o({\u2_Display/add67/c12 ,\u2_Display/n2102 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u12  (
    .a(\u2_Display/n2087 ),
    .b(1'b1),
    .c(\u2_Display/add67/c12 ),
    .o({\u2_Display/add67/c13 ,\u2_Display/n2102 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u13  (
    .a(\u2_Display/n2086 ),
    .b(1'b0),
    .c(\u2_Display/add67/c13 ),
    .o({\u2_Display/add67/c14 ,\u2_Display/n2102 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u14  (
    .a(\u2_Display/n2085 ),
    .b(1'b0),
    .c(\u2_Display/add67/c14 ),
    .o({\u2_Display/add67/c15 ,\u2_Display/n2102 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u15  (
    .a(\u2_Display/n2084 ),
    .b(1'b0),
    .c(\u2_Display/add67/c15 ),
    .o({\u2_Display/add67/c16 ,\u2_Display/n2102 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u16  (
    .a(\u2_Display/n2083 ),
    .b(1'b1),
    .c(\u2_Display/add67/c16 ),
    .o({\u2_Display/add67/c17 ,\u2_Display/n2102 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u17  (
    .a(\u2_Display/n2082 ),
    .b(1'b1),
    .c(\u2_Display/add67/c17 ),
    .o({\u2_Display/add67/c18 ,\u2_Display/n2102 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u18  (
    .a(\u2_Display/n2081 ),
    .b(1'b1),
    .c(\u2_Display/add67/c18 ),
    .o({\u2_Display/add67/c19 ,\u2_Display/n2102 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u19  (
    .a(\u2_Display/n2080 ),
    .b(1'b1),
    .c(\u2_Display/add67/c19 ),
    .o({\u2_Display/add67/c20 ,\u2_Display/n2102 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u2  (
    .a(\u2_Display/n2097 ),
    .b(1'b1),
    .c(\u2_Display/add67/c2 ),
    .o({\u2_Display/add67/c3 ,\u2_Display/n2102 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u20  (
    .a(\u2_Display/n2079 ),
    .b(1'b1),
    .c(\u2_Display/add67/c20 ),
    .o({\u2_Display/add67/c21 ,\u2_Display/n2102 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u21  (
    .a(\u2_Display/n2078 ),
    .b(1'b1),
    .c(\u2_Display/add67/c21 ),
    .o({\u2_Display/add67/c22 ,\u2_Display/n2102 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u22  (
    .a(\u2_Display/n2077 ),
    .b(1'b1),
    .c(\u2_Display/add67/c22 ),
    .o({\u2_Display/add67/c23 ,\u2_Display/n2102 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u23  (
    .a(\u2_Display/n2076 ),
    .b(1'b1),
    .c(\u2_Display/add67/c23 ),
    .o({\u2_Display/add67/c24 ,\u2_Display/n2102 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u24  (
    .a(\u2_Display/n2075 ),
    .b(1'b1),
    .c(\u2_Display/add67/c24 ),
    .o({\u2_Display/add67/c25 ,\u2_Display/n2102 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u25  (
    .a(\u2_Display/n2074 ),
    .b(1'b1),
    .c(\u2_Display/add67/c25 ),
    .o({\u2_Display/add67/c26 ,\u2_Display/n2102 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u26  (
    .a(\u2_Display/n2073 ),
    .b(1'b1),
    .c(\u2_Display/add67/c26 ),
    .o({\u2_Display/add67/c27 ,\u2_Display/n2102 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u27  (
    .a(\u2_Display/n2072 ),
    .b(1'b1),
    .c(\u2_Display/add67/c27 ),
    .o({\u2_Display/add67/c28 ,\u2_Display/n2102 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u28  (
    .a(\u2_Display/n2071 ),
    .b(1'b1),
    .c(\u2_Display/add67/c28 ),
    .o({\u2_Display/add67/c29 ,\u2_Display/n2102 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u29  (
    .a(\u2_Display/n2070 ),
    .b(1'b1),
    .c(\u2_Display/add67/c29 ),
    .o({\u2_Display/add67/c30 ,\u2_Display/n2102 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u3  (
    .a(\u2_Display/n2096 ),
    .b(1'b1),
    .c(\u2_Display/add67/c3 ),
    .o({\u2_Display/add67/c4 ,\u2_Display/n2102 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u30  (
    .a(\u2_Display/n2069 ),
    .b(1'b1),
    .c(\u2_Display/add67/c30 ),
    .o({\u2_Display/add67/c31 ,\u2_Display/n2102 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u31  (
    .a(\u2_Display/n2068 ),
    .b(1'b1),
    .c(\u2_Display/add67/c31 ),
    .o({open_n1259,\u2_Display/n2102 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u4  (
    .a(\u2_Display/n2095 ),
    .b(1'b1),
    .c(\u2_Display/add67/c4 ),
    .o({\u2_Display/add67/c5 ,\u2_Display/n2102 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u5  (
    .a(\u2_Display/n2094 ),
    .b(1'b1),
    .c(\u2_Display/add67/c5 ),
    .o({\u2_Display/add67/c6 ,\u2_Display/n2102 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u6  (
    .a(\u2_Display/n2093 ),
    .b(1'b1),
    .c(\u2_Display/add67/c6 ),
    .o({\u2_Display/add67/c7 ,\u2_Display/n2102 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u7  (
    .a(\u2_Display/n2092 ),
    .b(1'b1),
    .c(\u2_Display/add67/c7 ),
    .o({\u2_Display/add67/c8 ,\u2_Display/n2102 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u8  (
    .a(\u2_Display/n2091 ),
    .b(1'b0),
    .c(\u2_Display/add67/c8 ),
    .o({\u2_Display/add67/c9 ,\u2_Display/n2102 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add67/u9  (
    .a(\u2_Display/n2090 ),
    .b(1'b1),
    .c(\u2_Display/add67/c9 ),
    .o({\u2_Display/add67/c10 ,\u2_Display/n2102 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add67/ucin  (
    .a(1'b1),
    .o({\u2_Display/add67/c0 ,open_n1262}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u0  (
    .a(\u2_Display/n2134 ),
    .b(1'b1),
    .c(\u2_Display/add68/c0 ),
    .o({\u2_Display/add68/c1 ,\u2_Display/n2137 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u1  (
    .a(\u2_Display/n2133 ),
    .b(1'b1),
    .c(\u2_Display/add68/c1 ),
    .o({\u2_Display/add68/c2 ,\u2_Display/n2137 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u10  (
    .a(\u2_Display/n2124 ),
    .b(1'b1),
    .c(\u2_Display/add68/c10 ),
    .o({\u2_Display/add68/c11 ,\u2_Display/n2137 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u11  (
    .a(\u2_Display/n2123 ),
    .b(1'b1),
    .c(\u2_Display/add68/c11 ),
    .o({\u2_Display/add68/c12 ,\u2_Display/n2137 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u12  (
    .a(\u2_Display/n2122 ),
    .b(1'b0),
    .c(\u2_Display/add68/c12 ),
    .o({\u2_Display/add68/c13 ,\u2_Display/n2137 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u13  (
    .a(\u2_Display/n2121 ),
    .b(1'b0),
    .c(\u2_Display/add68/c13 ),
    .o({\u2_Display/add68/c14 ,\u2_Display/n2137 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u14  (
    .a(\u2_Display/n2120 ),
    .b(1'b0),
    .c(\u2_Display/add68/c14 ),
    .o({\u2_Display/add68/c15 ,\u2_Display/n2137 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u15  (
    .a(\u2_Display/n2119 ),
    .b(1'b1),
    .c(\u2_Display/add68/c15 ),
    .o({\u2_Display/add68/c16 ,\u2_Display/n2137 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u16  (
    .a(\u2_Display/n2118 ),
    .b(1'b1),
    .c(\u2_Display/add68/c16 ),
    .o({\u2_Display/add68/c17 ,\u2_Display/n2137 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u17  (
    .a(\u2_Display/n2117 ),
    .b(1'b1),
    .c(\u2_Display/add68/c17 ),
    .o({\u2_Display/add68/c18 ,\u2_Display/n2137 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u18  (
    .a(\u2_Display/n2116 ),
    .b(1'b1),
    .c(\u2_Display/add68/c18 ),
    .o({\u2_Display/add68/c19 ,\u2_Display/n2137 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u19  (
    .a(\u2_Display/n2115 ),
    .b(1'b1),
    .c(\u2_Display/add68/c19 ),
    .o({\u2_Display/add68/c20 ,\u2_Display/n2137 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u2  (
    .a(\u2_Display/n2132 ),
    .b(1'b1),
    .c(\u2_Display/add68/c2 ),
    .o({\u2_Display/add68/c3 ,\u2_Display/n2137 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u20  (
    .a(\u2_Display/n2114 ),
    .b(1'b1),
    .c(\u2_Display/add68/c20 ),
    .o({\u2_Display/add68/c21 ,\u2_Display/n2137 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u21  (
    .a(\u2_Display/n2113 ),
    .b(1'b1),
    .c(\u2_Display/add68/c21 ),
    .o({\u2_Display/add68/c22 ,\u2_Display/n2137 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u22  (
    .a(\u2_Display/n2112 ),
    .b(1'b1),
    .c(\u2_Display/add68/c22 ),
    .o({\u2_Display/add68/c23 ,\u2_Display/n2137 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u23  (
    .a(\u2_Display/n2111 ),
    .b(1'b1),
    .c(\u2_Display/add68/c23 ),
    .o({\u2_Display/add68/c24 ,\u2_Display/n2137 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u24  (
    .a(\u2_Display/n2110 ),
    .b(1'b1),
    .c(\u2_Display/add68/c24 ),
    .o({\u2_Display/add68/c25 ,\u2_Display/n2137 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u25  (
    .a(\u2_Display/n2109 ),
    .b(1'b1),
    .c(\u2_Display/add68/c25 ),
    .o({\u2_Display/add68/c26 ,\u2_Display/n2137 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u26  (
    .a(\u2_Display/n2108 ),
    .b(1'b1),
    .c(\u2_Display/add68/c26 ),
    .o({\u2_Display/add68/c27 ,\u2_Display/n2137 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u27  (
    .a(\u2_Display/n2107 ),
    .b(1'b1),
    .c(\u2_Display/add68/c27 ),
    .o({\u2_Display/add68/c28 ,\u2_Display/n2137 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u28  (
    .a(\u2_Display/n2106 ),
    .b(1'b1),
    .c(\u2_Display/add68/c28 ),
    .o({\u2_Display/add68/c29 ,\u2_Display/n2137 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u29  (
    .a(\u2_Display/n2105 ),
    .b(1'b1),
    .c(\u2_Display/add68/c29 ),
    .o({\u2_Display/add68/c30 ,\u2_Display/n2137 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u3  (
    .a(\u2_Display/n2131 ),
    .b(1'b1),
    .c(\u2_Display/add68/c3 ),
    .o({\u2_Display/add68/c4 ,\u2_Display/n2137 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u30  (
    .a(\u2_Display/n2104 ),
    .b(1'b1),
    .c(\u2_Display/add68/c30 ),
    .o({\u2_Display/add68/c31 ,\u2_Display/n2137 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u31  (
    .a(\u2_Display/n2103 ),
    .b(1'b1),
    .c(\u2_Display/add68/c31 ),
    .o({open_n1263,\u2_Display/n2137 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u4  (
    .a(\u2_Display/n2130 ),
    .b(1'b1),
    .c(\u2_Display/add68/c4 ),
    .o({\u2_Display/add68/c5 ,\u2_Display/n2137 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u5  (
    .a(\u2_Display/n2129 ),
    .b(1'b1),
    .c(\u2_Display/add68/c5 ),
    .o({\u2_Display/add68/c6 ,\u2_Display/n2137 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u6  (
    .a(\u2_Display/n2128 ),
    .b(1'b1),
    .c(\u2_Display/add68/c6 ),
    .o({\u2_Display/add68/c7 ,\u2_Display/n2137 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u7  (
    .a(\u2_Display/n2127 ),
    .b(1'b0),
    .c(\u2_Display/add68/c7 ),
    .o({\u2_Display/add68/c8 ,\u2_Display/n2137 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u8  (
    .a(\u2_Display/n2126 ),
    .b(1'b1),
    .c(\u2_Display/add68/c8 ),
    .o({\u2_Display/add68/c9 ,\u2_Display/n2137 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add68/u9  (
    .a(\u2_Display/n2125 ),
    .b(1'b1),
    .c(\u2_Display/add68/c9 ),
    .o({\u2_Display/add68/c10 ,\u2_Display/n2137 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add68/ucin  (
    .a(1'b1),
    .o({\u2_Display/add68/c0 ,open_n1266}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u0  (
    .a(\u2_Display/n2169 ),
    .b(1'b1),
    .c(\u2_Display/add69/c0 ),
    .o({\u2_Display/add69/c1 ,\u2_Display/n2172 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u1  (
    .a(\u2_Display/n2168 ),
    .b(1'b1),
    .c(\u2_Display/add69/c1 ),
    .o({\u2_Display/add69/c2 ,\u2_Display/n2172 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u10  (
    .a(\u2_Display/n2159 ),
    .b(1'b1),
    .c(\u2_Display/add69/c10 ),
    .o({\u2_Display/add69/c11 ,\u2_Display/n2172 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u11  (
    .a(\u2_Display/n2158 ),
    .b(1'b0),
    .c(\u2_Display/add69/c11 ),
    .o({\u2_Display/add69/c12 ,\u2_Display/n2172 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u12  (
    .a(\u2_Display/n2157 ),
    .b(1'b0),
    .c(\u2_Display/add69/c12 ),
    .o({\u2_Display/add69/c13 ,\u2_Display/n2172 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u13  (
    .a(\u2_Display/n2156 ),
    .b(1'b0),
    .c(\u2_Display/add69/c13 ),
    .o({\u2_Display/add69/c14 ,\u2_Display/n2172 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u14  (
    .a(\u2_Display/n2155 ),
    .b(1'b1),
    .c(\u2_Display/add69/c14 ),
    .o({\u2_Display/add69/c15 ,\u2_Display/n2172 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u15  (
    .a(\u2_Display/n2154 ),
    .b(1'b1),
    .c(\u2_Display/add69/c15 ),
    .o({\u2_Display/add69/c16 ,\u2_Display/n2172 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u16  (
    .a(\u2_Display/n2153 ),
    .b(1'b1),
    .c(\u2_Display/add69/c16 ),
    .o({\u2_Display/add69/c17 ,\u2_Display/n2172 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u17  (
    .a(\u2_Display/n2152 ),
    .b(1'b1),
    .c(\u2_Display/add69/c17 ),
    .o({\u2_Display/add69/c18 ,\u2_Display/n2172 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u18  (
    .a(\u2_Display/n2151 ),
    .b(1'b1),
    .c(\u2_Display/add69/c18 ),
    .o({\u2_Display/add69/c19 ,\u2_Display/n2172 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u19  (
    .a(\u2_Display/n2150 ),
    .b(1'b1),
    .c(\u2_Display/add69/c19 ),
    .o({\u2_Display/add69/c20 ,\u2_Display/n2172 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u2  (
    .a(\u2_Display/n2167 ),
    .b(1'b1),
    .c(\u2_Display/add69/c2 ),
    .o({\u2_Display/add69/c3 ,\u2_Display/n2172 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u20  (
    .a(\u2_Display/n2149 ),
    .b(1'b1),
    .c(\u2_Display/add69/c20 ),
    .o({\u2_Display/add69/c21 ,\u2_Display/n2172 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u21  (
    .a(\u2_Display/n2148 ),
    .b(1'b1),
    .c(\u2_Display/add69/c21 ),
    .o({\u2_Display/add69/c22 ,\u2_Display/n2172 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u22  (
    .a(\u2_Display/n2147 ),
    .b(1'b1),
    .c(\u2_Display/add69/c22 ),
    .o({\u2_Display/add69/c23 ,\u2_Display/n2172 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u23  (
    .a(\u2_Display/n2146 ),
    .b(1'b1),
    .c(\u2_Display/add69/c23 ),
    .o({\u2_Display/add69/c24 ,\u2_Display/n2172 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u24  (
    .a(\u2_Display/n2145 ),
    .b(1'b1),
    .c(\u2_Display/add69/c24 ),
    .o({\u2_Display/add69/c25 ,\u2_Display/n2172 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u25  (
    .a(\u2_Display/n2144 ),
    .b(1'b1),
    .c(\u2_Display/add69/c25 ),
    .o({\u2_Display/add69/c26 ,\u2_Display/n2172 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u26  (
    .a(\u2_Display/n2143 ),
    .b(1'b1),
    .c(\u2_Display/add69/c26 ),
    .o({\u2_Display/add69/c27 ,\u2_Display/n2172 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u27  (
    .a(\u2_Display/n2142 ),
    .b(1'b1),
    .c(\u2_Display/add69/c27 ),
    .o({\u2_Display/add69/c28 ,\u2_Display/n2172 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u28  (
    .a(\u2_Display/n2141 ),
    .b(1'b1),
    .c(\u2_Display/add69/c28 ),
    .o({\u2_Display/add69/c29 ,\u2_Display/n2172 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u29  (
    .a(\u2_Display/n2140 ),
    .b(1'b1),
    .c(\u2_Display/add69/c29 ),
    .o({\u2_Display/add69/c30 ,\u2_Display/n2172 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u3  (
    .a(\u2_Display/n2166 ),
    .b(1'b1),
    .c(\u2_Display/add69/c3 ),
    .o({\u2_Display/add69/c4 ,\u2_Display/n2172 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u30  (
    .a(\u2_Display/n2139 ),
    .b(1'b1),
    .c(\u2_Display/add69/c30 ),
    .o({\u2_Display/add69/c31 ,\u2_Display/n2172 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u31  (
    .a(\u2_Display/n2138 ),
    .b(1'b1),
    .c(\u2_Display/add69/c31 ),
    .o({open_n1267,\u2_Display/n2172 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u4  (
    .a(\u2_Display/n2165 ),
    .b(1'b1),
    .c(\u2_Display/add69/c4 ),
    .o({\u2_Display/add69/c5 ,\u2_Display/n2172 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u5  (
    .a(\u2_Display/n2164 ),
    .b(1'b1),
    .c(\u2_Display/add69/c5 ),
    .o({\u2_Display/add69/c6 ,\u2_Display/n2172 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u6  (
    .a(\u2_Display/n2163 ),
    .b(1'b0),
    .c(\u2_Display/add69/c6 ),
    .o({\u2_Display/add69/c7 ,\u2_Display/n2172 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u7  (
    .a(\u2_Display/n2162 ),
    .b(1'b1),
    .c(\u2_Display/add69/c7 ),
    .o({\u2_Display/add69/c8 ,\u2_Display/n2172 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u8  (
    .a(\u2_Display/n2161 ),
    .b(1'b1),
    .c(\u2_Display/add69/c8 ),
    .o({\u2_Display/add69/c9 ,\u2_Display/n2172 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add69/u9  (
    .a(\u2_Display/n2160 ),
    .b(1'b1),
    .c(\u2_Display/add69/c9 ),
    .o({\u2_Display/add69/c10 ,\u2_Display/n2172 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add69/ucin  (
    .a(1'b1),
    .o({\u2_Display/add69/c0 ,open_n1270}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add6_2/u0  (
    .a(1'b1),
    .b(\u2_Display/j [7]),
    .c(\u2_Display/add6_2/c0 ),
    .o({\u2_Display/add6_2/c1 ,\u2_Display/n135 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add6_2/u1  (
    .a(1'b0),
    .b(\u2_Display/j [8]),
    .c(\u2_Display/add6_2/c1 ),
    .o({\u2_Display/add6_2/c2 ,\u2_Display/n135 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add6_2/u2  (
    .a(1'b1),
    .b(\u2_Display/j [9]),
    .c(\u2_Display/add6_2/c2 ),
    .o({\u2_Display/add6_2/c3 ,\u2_Display/n135 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add6_2/ucin  (
    .a(1'b0),
    .o({\u2_Display/add6_2/c0 ,open_n1273}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add6_2/ucout  (
    .c(\u2_Display/add6_2/c3 ),
    .o({open_n1276,\u2_Display/add6_2_co }));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u0  (
    .a(\u2_Display/n2204 ),
    .b(1'b1),
    .c(\u2_Display/add70/c0 ),
    .o({\u2_Display/add70/c1 ,\u2_Display/n2207 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u1  (
    .a(\u2_Display/n2203 ),
    .b(1'b1),
    .c(\u2_Display/add70/c1 ),
    .o({\u2_Display/add70/c2 ,\u2_Display/n2207 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u10  (
    .a(\u2_Display/n2194 ),
    .b(1'b0),
    .c(\u2_Display/add70/c10 ),
    .o({\u2_Display/add70/c11 ,\u2_Display/n2207 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u11  (
    .a(\u2_Display/n2193 ),
    .b(1'b0),
    .c(\u2_Display/add70/c11 ),
    .o({\u2_Display/add70/c12 ,\u2_Display/n2207 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u12  (
    .a(\u2_Display/n2192 ),
    .b(1'b0),
    .c(\u2_Display/add70/c12 ),
    .o({\u2_Display/add70/c13 ,\u2_Display/n2207 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u13  (
    .a(\u2_Display/n2191 ),
    .b(1'b1),
    .c(\u2_Display/add70/c13 ),
    .o({\u2_Display/add70/c14 ,\u2_Display/n2207 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u14  (
    .a(\u2_Display/n2190 ),
    .b(1'b1),
    .c(\u2_Display/add70/c14 ),
    .o({\u2_Display/add70/c15 ,\u2_Display/n2207 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u15  (
    .a(\u2_Display/n2189 ),
    .b(1'b1),
    .c(\u2_Display/add70/c15 ),
    .o({\u2_Display/add70/c16 ,\u2_Display/n2207 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u16  (
    .a(\u2_Display/n2188 ),
    .b(1'b1),
    .c(\u2_Display/add70/c16 ),
    .o({\u2_Display/add70/c17 ,\u2_Display/n2207 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u17  (
    .a(\u2_Display/n2187 ),
    .b(1'b1),
    .c(\u2_Display/add70/c17 ),
    .o({\u2_Display/add70/c18 ,\u2_Display/n2207 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u18  (
    .a(\u2_Display/n2186 ),
    .b(1'b1),
    .c(\u2_Display/add70/c18 ),
    .o({\u2_Display/add70/c19 ,\u2_Display/n2207 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u19  (
    .a(\u2_Display/n2185 ),
    .b(1'b1),
    .c(\u2_Display/add70/c19 ),
    .o({\u2_Display/add70/c20 ,\u2_Display/n2207 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u2  (
    .a(\u2_Display/n2202 ),
    .b(1'b1),
    .c(\u2_Display/add70/c2 ),
    .o({\u2_Display/add70/c3 ,\u2_Display/n2207 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u20  (
    .a(\u2_Display/n2184 ),
    .b(1'b1),
    .c(\u2_Display/add70/c20 ),
    .o({\u2_Display/add70/c21 ,\u2_Display/n2207 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u21  (
    .a(\u2_Display/n2183 ),
    .b(1'b1),
    .c(\u2_Display/add70/c21 ),
    .o({\u2_Display/add70/c22 ,\u2_Display/n2207 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u22  (
    .a(\u2_Display/n2182 ),
    .b(1'b1),
    .c(\u2_Display/add70/c22 ),
    .o({\u2_Display/add70/c23 ,\u2_Display/n2207 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u23  (
    .a(\u2_Display/n2181 ),
    .b(1'b1),
    .c(\u2_Display/add70/c23 ),
    .o({\u2_Display/add70/c24 ,\u2_Display/n2207 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u24  (
    .a(\u2_Display/n2180 ),
    .b(1'b1),
    .c(\u2_Display/add70/c24 ),
    .o({\u2_Display/add70/c25 ,\u2_Display/n2207 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u25  (
    .a(\u2_Display/n2179 ),
    .b(1'b1),
    .c(\u2_Display/add70/c25 ),
    .o({\u2_Display/add70/c26 ,\u2_Display/n2207 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u26  (
    .a(\u2_Display/n2178 ),
    .b(1'b1),
    .c(\u2_Display/add70/c26 ),
    .o({\u2_Display/add70/c27 ,\u2_Display/n2207 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u27  (
    .a(\u2_Display/n2177 ),
    .b(1'b1),
    .c(\u2_Display/add70/c27 ),
    .o({\u2_Display/add70/c28 ,\u2_Display/n2207 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u28  (
    .a(\u2_Display/n2176 ),
    .b(1'b1),
    .c(\u2_Display/add70/c28 ),
    .o({\u2_Display/add70/c29 ,\u2_Display/n2207 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u29  (
    .a(\u2_Display/n2175 ),
    .b(1'b1),
    .c(\u2_Display/add70/c29 ),
    .o({\u2_Display/add70/c30 ,\u2_Display/n2207 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u3  (
    .a(\u2_Display/n2201 ),
    .b(1'b1),
    .c(\u2_Display/add70/c3 ),
    .o({\u2_Display/add70/c4 ,\u2_Display/n2207 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u30  (
    .a(\u2_Display/n2174 ),
    .b(1'b1),
    .c(\u2_Display/add70/c30 ),
    .o({\u2_Display/add70/c31 ,\u2_Display/n2207 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u31  (
    .a(\u2_Display/n2173 ),
    .b(1'b1),
    .c(\u2_Display/add70/c31 ),
    .o({open_n1277,\u2_Display/n2207 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u4  (
    .a(\u2_Display/n2200 ),
    .b(1'b1),
    .c(\u2_Display/add70/c4 ),
    .o({\u2_Display/add70/c5 ,\u2_Display/n2207 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u5  (
    .a(\u2_Display/n2199 ),
    .b(1'b0),
    .c(\u2_Display/add70/c5 ),
    .o({\u2_Display/add70/c6 ,\u2_Display/n2207 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u6  (
    .a(\u2_Display/n2198 ),
    .b(1'b1),
    .c(\u2_Display/add70/c6 ),
    .o({\u2_Display/add70/c7 ,\u2_Display/n2207 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u7  (
    .a(\u2_Display/n2197 ),
    .b(1'b1),
    .c(\u2_Display/add70/c7 ),
    .o({\u2_Display/add70/c8 ,\u2_Display/n2207 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u8  (
    .a(\u2_Display/n2196 ),
    .b(1'b1),
    .c(\u2_Display/add70/c8 ),
    .o({\u2_Display/add70/c9 ,\u2_Display/n2207 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add70/u9  (
    .a(\u2_Display/n2195 ),
    .b(1'b1),
    .c(\u2_Display/add70/c9 ),
    .o({\u2_Display/add70/c10 ,\u2_Display/n2207 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add70/ucin  (
    .a(1'b1),
    .o({\u2_Display/add70/c0 ,open_n1280}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u0  (
    .a(\u2_Display/n2239 ),
    .b(1'b1),
    .c(\u2_Display/add71/c0 ),
    .o({\u2_Display/add71/c1 ,\u2_Display/n2242 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u1  (
    .a(\u2_Display/n2238 ),
    .b(1'b1),
    .c(\u2_Display/add71/c1 ),
    .o({\u2_Display/add71/c2 ,\u2_Display/n2242 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u10  (
    .a(\u2_Display/n2229 ),
    .b(1'b0),
    .c(\u2_Display/add71/c10 ),
    .o({\u2_Display/add71/c11 ,\u2_Display/n2242 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u11  (
    .a(\u2_Display/n2228 ),
    .b(1'b0),
    .c(\u2_Display/add71/c11 ),
    .o({\u2_Display/add71/c12 ,\u2_Display/n2242 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u12  (
    .a(\u2_Display/n2227 ),
    .b(1'b1),
    .c(\u2_Display/add71/c12 ),
    .o({\u2_Display/add71/c13 ,\u2_Display/n2242 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u13  (
    .a(\u2_Display/n2226 ),
    .b(1'b1),
    .c(\u2_Display/add71/c13 ),
    .o({\u2_Display/add71/c14 ,\u2_Display/n2242 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u14  (
    .a(\u2_Display/n2225 ),
    .b(1'b1),
    .c(\u2_Display/add71/c14 ),
    .o({\u2_Display/add71/c15 ,\u2_Display/n2242 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u15  (
    .a(\u2_Display/n2224 ),
    .b(1'b1),
    .c(\u2_Display/add71/c15 ),
    .o({\u2_Display/add71/c16 ,\u2_Display/n2242 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u16  (
    .a(\u2_Display/n2223 ),
    .b(1'b1),
    .c(\u2_Display/add71/c16 ),
    .o({\u2_Display/add71/c17 ,\u2_Display/n2242 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u17  (
    .a(\u2_Display/n2222 ),
    .b(1'b1),
    .c(\u2_Display/add71/c17 ),
    .o({\u2_Display/add71/c18 ,\u2_Display/n2242 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u18  (
    .a(\u2_Display/n2221 ),
    .b(1'b1),
    .c(\u2_Display/add71/c18 ),
    .o({\u2_Display/add71/c19 ,\u2_Display/n2242 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u19  (
    .a(\u2_Display/n2220 ),
    .b(1'b1),
    .c(\u2_Display/add71/c19 ),
    .o({\u2_Display/add71/c20 ,\u2_Display/n2242 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u2  (
    .a(\u2_Display/n2237 ),
    .b(1'b1),
    .c(\u2_Display/add71/c2 ),
    .o({\u2_Display/add71/c3 ,\u2_Display/n2242 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u20  (
    .a(\u2_Display/n2219 ),
    .b(1'b1),
    .c(\u2_Display/add71/c20 ),
    .o({\u2_Display/add71/c21 ,\u2_Display/n2242 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u21  (
    .a(\u2_Display/n2218 ),
    .b(1'b1),
    .c(\u2_Display/add71/c21 ),
    .o({\u2_Display/add71/c22 ,\u2_Display/n2242 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u22  (
    .a(\u2_Display/n2217 ),
    .b(1'b1),
    .c(\u2_Display/add71/c22 ),
    .o({\u2_Display/add71/c23 ,\u2_Display/n2242 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u23  (
    .a(\u2_Display/n2216 ),
    .b(1'b1),
    .c(\u2_Display/add71/c23 ),
    .o({\u2_Display/add71/c24 ,\u2_Display/n2242 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u24  (
    .a(\u2_Display/n2215 ),
    .b(1'b1),
    .c(\u2_Display/add71/c24 ),
    .o({\u2_Display/add71/c25 ,\u2_Display/n2242 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u25  (
    .a(\u2_Display/n2214 ),
    .b(1'b1),
    .c(\u2_Display/add71/c25 ),
    .o({\u2_Display/add71/c26 ,\u2_Display/n2242 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u26  (
    .a(\u2_Display/n2213 ),
    .b(1'b1),
    .c(\u2_Display/add71/c26 ),
    .o({\u2_Display/add71/c27 ,\u2_Display/n2242 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u27  (
    .a(\u2_Display/n2212 ),
    .b(1'b1),
    .c(\u2_Display/add71/c27 ),
    .o({\u2_Display/add71/c28 ,\u2_Display/n2242 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u28  (
    .a(\u2_Display/n2211 ),
    .b(1'b1),
    .c(\u2_Display/add71/c28 ),
    .o({\u2_Display/add71/c29 ,\u2_Display/n2242 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u29  (
    .a(\u2_Display/n2210 ),
    .b(1'b1),
    .c(\u2_Display/add71/c29 ),
    .o({\u2_Display/add71/c30 ,\u2_Display/n2242 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u3  (
    .a(\u2_Display/n2236 ),
    .b(1'b1),
    .c(\u2_Display/add71/c3 ),
    .o({\u2_Display/add71/c4 ,\u2_Display/n2242 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u30  (
    .a(\u2_Display/n2209 ),
    .b(1'b1),
    .c(\u2_Display/add71/c30 ),
    .o({\u2_Display/add71/c31 ,\u2_Display/n2242 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u31  (
    .a(\u2_Display/n2208 ),
    .b(1'b1),
    .c(\u2_Display/add71/c31 ),
    .o({open_n1281,\u2_Display/n2242 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u4  (
    .a(\u2_Display/n2235 ),
    .b(1'b0),
    .c(\u2_Display/add71/c4 ),
    .o({\u2_Display/add71/c5 ,\u2_Display/n2242 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u5  (
    .a(\u2_Display/n2234 ),
    .b(1'b1),
    .c(\u2_Display/add71/c5 ),
    .o({\u2_Display/add71/c6 ,\u2_Display/n2242 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u6  (
    .a(\u2_Display/n2233 ),
    .b(1'b1),
    .c(\u2_Display/add71/c6 ),
    .o({\u2_Display/add71/c7 ,\u2_Display/n2242 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u7  (
    .a(\u2_Display/n2232 ),
    .b(1'b1),
    .c(\u2_Display/add71/c7 ),
    .o({\u2_Display/add71/c8 ,\u2_Display/n2242 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u8  (
    .a(\u2_Display/n2231 ),
    .b(1'b1),
    .c(\u2_Display/add71/c8 ),
    .o({\u2_Display/add71/c9 ,\u2_Display/n2242 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add71/u9  (
    .a(\u2_Display/n2230 ),
    .b(1'b0),
    .c(\u2_Display/add71/c9 ),
    .o({\u2_Display/add71/c10 ,\u2_Display/n2242 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add71/ucin  (
    .a(1'b1),
    .o({\u2_Display/add71/c0 ,open_n1284}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u0  (
    .a(\u2_Display/n2274 ),
    .b(1'b1),
    .c(\u2_Display/add72/c0 ),
    .o({\u2_Display/add72/c1 ,\u2_Display/n2277 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u1  (
    .a(\u2_Display/n2273 ),
    .b(1'b1),
    .c(\u2_Display/add72/c1 ),
    .o({\u2_Display/add72/c2 ,\u2_Display/n2277 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u10  (
    .a(\u2_Display/n2264 ),
    .b(1'b0),
    .c(\u2_Display/add72/c10 ),
    .o({\u2_Display/add72/c11 ,\u2_Display/n2277 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u11  (
    .a(\u2_Display/n2263 ),
    .b(1'b1),
    .c(\u2_Display/add72/c11 ),
    .o({\u2_Display/add72/c12 ,\u2_Display/n2277 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u12  (
    .a(\u2_Display/n2262 ),
    .b(1'b1),
    .c(\u2_Display/add72/c12 ),
    .o({\u2_Display/add72/c13 ,\u2_Display/n2277 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u13  (
    .a(\u2_Display/n2261 ),
    .b(1'b1),
    .c(\u2_Display/add72/c13 ),
    .o({\u2_Display/add72/c14 ,\u2_Display/n2277 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u14  (
    .a(\u2_Display/n2260 ),
    .b(1'b1),
    .c(\u2_Display/add72/c14 ),
    .o({\u2_Display/add72/c15 ,\u2_Display/n2277 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u15  (
    .a(\u2_Display/n2259 ),
    .b(1'b1),
    .c(\u2_Display/add72/c15 ),
    .o({\u2_Display/add72/c16 ,\u2_Display/n2277 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u16  (
    .a(\u2_Display/n2258 ),
    .b(1'b1),
    .c(\u2_Display/add72/c16 ),
    .o({\u2_Display/add72/c17 ,\u2_Display/n2277 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u17  (
    .a(\u2_Display/n2257 ),
    .b(1'b1),
    .c(\u2_Display/add72/c17 ),
    .o({\u2_Display/add72/c18 ,\u2_Display/n2277 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u18  (
    .a(\u2_Display/n2256 ),
    .b(1'b1),
    .c(\u2_Display/add72/c18 ),
    .o({\u2_Display/add72/c19 ,\u2_Display/n2277 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u19  (
    .a(\u2_Display/n2255 ),
    .b(1'b1),
    .c(\u2_Display/add72/c19 ),
    .o({\u2_Display/add72/c20 ,\u2_Display/n2277 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u2  (
    .a(\u2_Display/n2272 ),
    .b(1'b1),
    .c(\u2_Display/add72/c2 ),
    .o({\u2_Display/add72/c3 ,\u2_Display/n2277 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u20  (
    .a(\u2_Display/n2254 ),
    .b(1'b1),
    .c(\u2_Display/add72/c20 ),
    .o({\u2_Display/add72/c21 ,\u2_Display/n2277 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u21  (
    .a(\u2_Display/n2253 ),
    .b(1'b1),
    .c(\u2_Display/add72/c21 ),
    .o({\u2_Display/add72/c22 ,\u2_Display/n2277 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u22  (
    .a(\u2_Display/n2252 ),
    .b(1'b1),
    .c(\u2_Display/add72/c22 ),
    .o({\u2_Display/add72/c23 ,\u2_Display/n2277 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u23  (
    .a(\u2_Display/n2251 ),
    .b(1'b1),
    .c(\u2_Display/add72/c23 ),
    .o({\u2_Display/add72/c24 ,\u2_Display/n2277 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u24  (
    .a(\u2_Display/n2250 ),
    .b(1'b1),
    .c(\u2_Display/add72/c24 ),
    .o({\u2_Display/add72/c25 ,\u2_Display/n2277 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u25  (
    .a(\u2_Display/n2249 ),
    .b(1'b1),
    .c(\u2_Display/add72/c25 ),
    .o({\u2_Display/add72/c26 ,\u2_Display/n2277 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u26  (
    .a(\u2_Display/n2248 ),
    .b(1'b1),
    .c(\u2_Display/add72/c26 ),
    .o({\u2_Display/add72/c27 ,\u2_Display/n2277 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u27  (
    .a(\u2_Display/n2247 ),
    .b(1'b1),
    .c(\u2_Display/add72/c27 ),
    .o({\u2_Display/add72/c28 ,\u2_Display/n2277 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u28  (
    .a(\u2_Display/n2246 ),
    .b(1'b1),
    .c(\u2_Display/add72/c28 ),
    .o({\u2_Display/add72/c29 ,\u2_Display/n2277 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u29  (
    .a(\u2_Display/n2245 ),
    .b(1'b1),
    .c(\u2_Display/add72/c29 ),
    .o({\u2_Display/add72/c30 ,\u2_Display/n2277 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u3  (
    .a(\u2_Display/n2271 ),
    .b(1'b0),
    .c(\u2_Display/add72/c3 ),
    .o({\u2_Display/add72/c4 ,\u2_Display/n2277 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u30  (
    .a(\u2_Display/n2244 ),
    .b(1'b1),
    .c(\u2_Display/add72/c30 ),
    .o({\u2_Display/add72/c31 ,\u2_Display/n2277 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u31  (
    .a(\u2_Display/n2243 ),
    .b(1'b1),
    .c(\u2_Display/add72/c31 ),
    .o({open_n1285,\u2_Display/n2277 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u4  (
    .a(\u2_Display/n2270 ),
    .b(1'b1),
    .c(\u2_Display/add72/c4 ),
    .o({\u2_Display/add72/c5 ,\u2_Display/n2277 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u5  (
    .a(\u2_Display/n2269 ),
    .b(1'b1),
    .c(\u2_Display/add72/c5 ),
    .o({\u2_Display/add72/c6 ,\u2_Display/n2277 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u6  (
    .a(\u2_Display/n2268 ),
    .b(1'b1),
    .c(\u2_Display/add72/c6 ),
    .o({\u2_Display/add72/c7 ,\u2_Display/n2277 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u7  (
    .a(\u2_Display/n2267 ),
    .b(1'b1),
    .c(\u2_Display/add72/c7 ),
    .o({\u2_Display/add72/c8 ,\u2_Display/n2277 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u8  (
    .a(\u2_Display/n2266 ),
    .b(1'b0),
    .c(\u2_Display/add72/c8 ),
    .o({\u2_Display/add72/c9 ,\u2_Display/n2277 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add72/u9  (
    .a(\u2_Display/n2265 ),
    .b(1'b0),
    .c(\u2_Display/add72/c9 ),
    .o({\u2_Display/add72/c10 ,\u2_Display/n2277 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add72/ucin  (
    .a(1'b1),
    .o({\u2_Display/add72/c0 ,open_n1288}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add73/u0  (
    .a(\u2_Display/n2309 ),
    .b(1'b1),
    .c(\u2_Display/add73/c0 ),
    .o({\u2_Display/add73/c1 ,\u2_Display/n2312 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add73/u1  (
    .a(\u2_Display/n2308 ),
    .b(1'b1),
    .c(\u2_Display/add73/c1 ),
    .o({\u2_Display/add73/c2 ,\u2_Display/n2312 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add73/u2  (
    .a(\u2_Display/n2307 ),
    .b(1'b0),
    .c(\u2_Display/add73/c2 ),
    .o({\u2_Display/add73/c3 ,\u2_Display/n2312 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add73/u3  (
    .a(\u2_Display/n2306 ),
    .b(1'b1),
    .c(\u2_Display/add73/c3 ),
    .o({\u2_Display/add73/c4 ,\u2_Display/n2312 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add73/u4  (
    .a(\u2_Display/n2305 ),
    .b(1'b1),
    .c(\u2_Display/add73/c4 ),
    .o({\u2_Display/add73/c5 ,\u2_Display/n2312 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add73/u5  (
    .a(\u2_Display/n2304 ),
    .b(1'b1),
    .c(\u2_Display/add73/c5 ),
    .o({\u2_Display/add73/c6 ,\u2_Display/n2312 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add73/u6  (
    .a(\u2_Display/n2303 ),
    .b(1'b1),
    .c(\u2_Display/add73/c6 ),
    .o({\u2_Display/add73/c7 ,\u2_Display/n2312 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add73/u7  (
    .a(\u2_Display/n2302 ),
    .b(1'b0),
    .c(\u2_Display/add73/c7 ),
    .o({\u2_Display/add73/c8 ,\u2_Display/n2312 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add73/u8  (
    .a(\u2_Display/n2301 ),
    .b(1'b0),
    .c(\u2_Display/add73/c8 ),
    .o({\u2_Display/add73/c9 ,\u2_Display/n2312 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add73/u9  (
    .a(\u2_Display/n2300 ),
    .b(1'b0),
    .c(\u2_Display/add73/c9 ),
    .o({open_n1289,\u2_Display/n2312 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add73/ucin  (
    .a(1'b1),
    .o({\u2_Display/add73/c0 ,open_n1292}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u0  (
    .a(\u2_Display/counta [0]),
    .b(1'b1),
    .c(\u2_Display/add84/c0 ),
    .o({\u2_Display/add84/c1 ,\u2_Display/n2665 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u1  (
    .a(\u2_Display/counta [1]),
    .b(1'b1),
    .c(\u2_Display/add84/c1 ),
    .o({\u2_Display/add84/c2 ,\u2_Display/n2665 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u10  (
    .a(\u2_Display/counta [10]),
    .b(1'b1),
    .c(\u2_Display/add84/c10 ),
    .o({\u2_Display/add84/c11 ,\u2_Display/n2665 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u11  (
    .a(\u2_Display/counta [11]),
    .b(1'b1),
    .c(\u2_Display/add84/c11 ),
    .o({\u2_Display/add84/c12 ,\u2_Display/n2665 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u12  (
    .a(\u2_Display/counta [12]),
    .b(1'b1),
    .c(\u2_Display/add84/c12 ),
    .o({\u2_Display/add84/c13 ,\u2_Display/n2665 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u13  (
    .a(\u2_Display/counta [13]),
    .b(1'b1),
    .c(\u2_Display/add84/c13 ),
    .o({\u2_Display/add84/c14 ,\u2_Display/n2665 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u14  (
    .a(\u2_Display/counta [14]),
    .b(1'b1),
    .c(\u2_Display/add84/c14 ),
    .o({\u2_Display/add84/c15 ,\u2_Display/n2665 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u15  (
    .a(\u2_Display/counta [15]),
    .b(1'b1),
    .c(\u2_Display/add84/c15 ),
    .o({\u2_Display/add84/c16 ,\u2_Display/n2665 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u16  (
    .a(\u2_Display/counta [16]),
    .b(1'b1),
    .c(\u2_Display/add84/c16 ),
    .o({\u2_Display/add84/c17 ,\u2_Display/n2665 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u17  (
    .a(\u2_Display/counta [17]),
    .b(1'b1),
    .c(\u2_Display/add84/c17 ),
    .o({\u2_Display/add84/c18 ,\u2_Display/n2665 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u18  (
    .a(\u2_Display/counta [18]),
    .b(1'b1),
    .c(\u2_Display/add84/c18 ),
    .o({\u2_Display/add84/c19 ,\u2_Display/n2665 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u19  (
    .a(\u2_Display/counta [19]),
    .b(1'b1),
    .c(\u2_Display/add84/c19 ),
    .o({\u2_Display/add84/c20 ,\u2_Display/n2665 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u2  (
    .a(\u2_Display/counta [2]),
    .b(1'b1),
    .c(\u2_Display/add84/c2 ),
    .o({\u2_Display/add84/c3 ,\u2_Display/n2665 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u20  (
    .a(\u2_Display/counta [20]),
    .b(1'b1),
    .c(\u2_Display/add84/c20 ),
    .o({\u2_Display/add84/c21 ,\u2_Display/n2665 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u21  (
    .a(\u2_Display/counta [21]),
    .b(1'b1),
    .c(\u2_Display/add84/c21 ),
    .o({\u2_Display/add84/c22 ,\u2_Display/n2665 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u22  (
    .a(\u2_Display/counta [22]),
    .b(1'b1),
    .c(\u2_Display/add84/c22 ),
    .o({\u2_Display/add84/c23 ,\u2_Display/n2665 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u23  (
    .a(\u2_Display/counta [23]),
    .b(1'b1),
    .c(\u2_Display/add84/c23 ),
    .o({\u2_Display/add84/c24 ,\u2_Display/n2665 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u24  (
    .a(\u2_Display/counta [24]),
    .b(1'b1),
    .c(\u2_Display/add84/c24 ),
    .o({\u2_Display/add84/c25 ,\u2_Display/n2665 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u25  (
    .a(\u2_Display/counta [25]),
    .b(1'b0),
    .c(\u2_Display/add84/c25 ),
    .o({\u2_Display/add84/c26 ,\u2_Display/n2665 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u26  (
    .a(\u2_Display/counta [26]),
    .b(1'b0),
    .c(\u2_Display/add84/c26 ),
    .o({\u2_Display/add84/c27 ,\u2_Display/n2665 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u27  (
    .a(\u2_Display/counta [27]),
    .b(1'b1),
    .c(\u2_Display/add84/c27 ),
    .o({\u2_Display/add84/c28 ,\u2_Display/n2665 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u28  (
    .a(\u2_Display/counta [28]),
    .b(1'b0),
    .c(\u2_Display/add84/c28 ),
    .o({\u2_Display/add84/c29 ,\u2_Display/n2665 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u29  (
    .a(\u2_Display/counta [29]),
    .b(1'b1),
    .c(\u2_Display/add84/c29 ),
    .o({\u2_Display/add84/c30 ,\u2_Display/n2665 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u3  (
    .a(\u2_Display/counta [3]),
    .b(1'b1),
    .c(\u2_Display/add84/c3 ),
    .o({\u2_Display/add84/c4 ,\u2_Display/n2665 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u30  (
    .a(\u2_Display/counta [30]),
    .b(1'b1),
    .c(\u2_Display/add84/c30 ),
    .o({\u2_Display/add84/c31 ,\u2_Display/n2665 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u31  (
    .a(\u2_Display/counta [31]),
    .b(1'b0),
    .c(\u2_Display/add84/c31 ),
    .o({open_n1293,\u2_Display/n2665 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u4  (
    .a(\u2_Display/counta [4]),
    .b(1'b1),
    .c(\u2_Display/add84/c4 ),
    .o({\u2_Display/add84/c5 ,\u2_Display/n2665 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u5  (
    .a(\u2_Display/counta [5]),
    .b(1'b1),
    .c(\u2_Display/add84/c5 ),
    .o({\u2_Display/add84/c6 ,\u2_Display/n2665 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u6  (
    .a(\u2_Display/counta [6]),
    .b(1'b1),
    .c(\u2_Display/add84/c6 ),
    .o({\u2_Display/add84/c7 ,\u2_Display/n2665 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u7  (
    .a(\u2_Display/counta [7]),
    .b(1'b1),
    .c(\u2_Display/add84/c7 ),
    .o({\u2_Display/add84/c8 ,\u2_Display/n2665 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u8  (
    .a(\u2_Display/counta [8]),
    .b(1'b1),
    .c(\u2_Display/add84/c8 ),
    .o({\u2_Display/add84/c9 ,\u2_Display/n2665 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add84/u9  (
    .a(\u2_Display/counta [9]),
    .b(1'b1),
    .c(\u2_Display/add84/c9 ),
    .o({\u2_Display/add84/c10 ,\u2_Display/n2665 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add84/ucin  (
    .a(1'b1),
    .o({\u2_Display/add84/c0 ,open_n1296}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u0  (
    .a(\u2_Display/n2697 ),
    .b(1'b1),
    .c(\u2_Display/add85/c0 ),
    .o({\u2_Display/add85/c1 ,\u2_Display/n2700 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u1  (
    .a(\u2_Display/n2696 ),
    .b(1'b1),
    .c(\u2_Display/add85/c1 ),
    .o({\u2_Display/add85/c2 ,\u2_Display/n2700 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u10  (
    .a(\u2_Display/n2687 ),
    .b(1'b1),
    .c(\u2_Display/add85/c10 ),
    .o({\u2_Display/add85/c11 ,\u2_Display/n2700 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u11  (
    .a(\u2_Display/n2686 ),
    .b(1'b1),
    .c(\u2_Display/add85/c11 ),
    .o({\u2_Display/add85/c12 ,\u2_Display/n2700 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u12  (
    .a(\u2_Display/n2685 ),
    .b(1'b1),
    .c(\u2_Display/add85/c12 ),
    .o({\u2_Display/add85/c13 ,\u2_Display/n2700 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u13  (
    .a(\u2_Display/n2684 ),
    .b(1'b1),
    .c(\u2_Display/add85/c13 ),
    .o({\u2_Display/add85/c14 ,\u2_Display/n2700 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u14  (
    .a(\u2_Display/n2683 ),
    .b(1'b1),
    .c(\u2_Display/add85/c14 ),
    .o({\u2_Display/add85/c15 ,\u2_Display/n2700 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u15  (
    .a(\u2_Display/n2682 ),
    .b(1'b1),
    .c(\u2_Display/add85/c15 ),
    .o({\u2_Display/add85/c16 ,\u2_Display/n2700 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u16  (
    .a(\u2_Display/n2681 ),
    .b(1'b1),
    .c(\u2_Display/add85/c16 ),
    .o({\u2_Display/add85/c17 ,\u2_Display/n2700 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u17  (
    .a(\u2_Display/n2680 ),
    .b(1'b1),
    .c(\u2_Display/add85/c17 ),
    .o({\u2_Display/add85/c18 ,\u2_Display/n2700 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u18  (
    .a(\u2_Display/n2679 ),
    .b(1'b1),
    .c(\u2_Display/add85/c18 ),
    .o({\u2_Display/add85/c19 ,\u2_Display/n2700 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u19  (
    .a(\u2_Display/n2678 ),
    .b(1'b1),
    .c(\u2_Display/add85/c19 ),
    .o({\u2_Display/add85/c20 ,\u2_Display/n2700 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u2  (
    .a(\u2_Display/n2695 ),
    .b(1'b1),
    .c(\u2_Display/add85/c2 ),
    .o({\u2_Display/add85/c3 ,\u2_Display/n2700 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u20  (
    .a(\u2_Display/n2677 ),
    .b(1'b1),
    .c(\u2_Display/add85/c20 ),
    .o({\u2_Display/add85/c21 ,\u2_Display/n2700 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u21  (
    .a(\u2_Display/n2676 ),
    .b(1'b1),
    .c(\u2_Display/add85/c21 ),
    .o({\u2_Display/add85/c22 ,\u2_Display/n2700 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u22  (
    .a(\u2_Display/n2675 ),
    .b(1'b1),
    .c(\u2_Display/add85/c22 ),
    .o({\u2_Display/add85/c23 ,\u2_Display/n2700 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u23  (
    .a(\u2_Display/n2674 ),
    .b(1'b1),
    .c(\u2_Display/add85/c23 ),
    .o({\u2_Display/add85/c24 ,\u2_Display/n2700 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u24  (
    .a(\u2_Display/n2673 ),
    .b(1'b0),
    .c(\u2_Display/add85/c24 ),
    .o({\u2_Display/add85/c25 ,\u2_Display/n2700 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u25  (
    .a(\u2_Display/n2672 ),
    .b(1'b0),
    .c(\u2_Display/add85/c25 ),
    .o({\u2_Display/add85/c26 ,\u2_Display/n2700 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u26  (
    .a(\u2_Display/n2671 ),
    .b(1'b1),
    .c(\u2_Display/add85/c26 ),
    .o({\u2_Display/add85/c27 ,\u2_Display/n2700 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u27  (
    .a(\u2_Display/n2670 ),
    .b(1'b0),
    .c(\u2_Display/add85/c27 ),
    .o({\u2_Display/add85/c28 ,\u2_Display/n2700 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u28  (
    .a(\u2_Display/n2669 ),
    .b(1'b1),
    .c(\u2_Display/add85/c28 ),
    .o({\u2_Display/add85/c29 ,\u2_Display/n2700 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u29  (
    .a(\u2_Display/n2668 ),
    .b(1'b1),
    .c(\u2_Display/add85/c29 ),
    .o({\u2_Display/add85/c30 ,\u2_Display/n2700 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u3  (
    .a(\u2_Display/n2694 ),
    .b(1'b1),
    .c(\u2_Display/add85/c3 ),
    .o({\u2_Display/add85/c4 ,\u2_Display/n2700 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u30  (
    .a(\u2_Display/n2667 ),
    .b(1'b0),
    .c(\u2_Display/add85/c30 ),
    .o({\u2_Display/add85/c31 ,\u2_Display/n2700 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u31  (
    .a(\u2_Display/n2666 ),
    .b(1'b1),
    .c(\u2_Display/add85/c31 ),
    .o({open_n1297,\u2_Display/n2700 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u4  (
    .a(\u2_Display/n2693 ),
    .b(1'b1),
    .c(\u2_Display/add85/c4 ),
    .o({\u2_Display/add85/c5 ,\u2_Display/n2700 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u5  (
    .a(\u2_Display/n2692 ),
    .b(1'b1),
    .c(\u2_Display/add85/c5 ),
    .o({\u2_Display/add85/c6 ,\u2_Display/n2700 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u6  (
    .a(\u2_Display/n2691 ),
    .b(1'b1),
    .c(\u2_Display/add85/c6 ),
    .o({\u2_Display/add85/c7 ,\u2_Display/n2700 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u7  (
    .a(\u2_Display/n2690 ),
    .b(1'b1),
    .c(\u2_Display/add85/c7 ),
    .o({\u2_Display/add85/c8 ,\u2_Display/n2700 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u8  (
    .a(\u2_Display/n2689 ),
    .b(1'b1),
    .c(\u2_Display/add85/c8 ),
    .o({\u2_Display/add85/c9 ,\u2_Display/n2700 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add85/u9  (
    .a(\u2_Display/n2688 ),
    .b(1'b1),
    .c(\u2_Display/add85/c9 ),
    .o({\u2_Display/add85/c10 ,\u2_Display/n2700 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add85/ucin  (
    .a(1'b1),
    .o({\u2_Display/add85/c0 ,open_n1300}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u0  (
    .a(\u2_Display/n2732 ),
    .b(1'b1),
    .c(\u2_Display/add86/c0 ),
    .o({\u2_Display/add86/c1 ,\u2_Display/n2735 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u1  (
    .a(\u2_Display/n2731 ),
    .b(1'b1),
    .c(\u2_Display/add86/c1 ),
    .o({\u2_Display/add86/c2 ,\u2_Display/n2735 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u10  (
    .a(\u2_Display/n2722 ),
    .b(1'b1),
    .c(\u2_Display/add86/c10 ),
    .o({\u2_Display/add86/c11 ,\u2_Display/n2735 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u11  (
    .a(\u2_Display/n2721 ),
    .b(1'b1),
    .c(\u2_Display/add86/c11 ),
    .o({\u2_Display/add86/c12 ,\u2_Display/n2735 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u12  (
    .a(\u2_Display/n2720 ),
    .b(1'b1),
    .c(\u2_Display/add86/c12 ),
    .o({\u2_Display/add86/c13 ,\u2_Display/n2735 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u13  (
    .a(\u2_Display/n2719 ),
    .b(1'b1),
    .c(\u2_Display/add86/c13 ),
    .o({\u2_Display/add86/c14 ,\u2_Display/n2735 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u14  (
    .a(\u2_Display/n2718 ),
    .b(1'b1),
    .c(\u2_Display/add86/c14 ),
    .o({\u2_Display/add86/c15 ,\u2_Display/n2735 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u15  (
    .a(\u2_Display/n2717 ),
    .b(1'b1),
    .c(\u2_Display/add86/c15 ),
    .o({\u2_Display/add86/c16 ,\u2_Display/n2735 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u16  (
    .a(\u2_Display/n2716 ),
    .b(1'b1),
    .c(\u2_Display/add86/c16 ),
    .o({\u2_Display/add86/c17 ,\u2_Display/n2735 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u17  (
    .a(\u2_Display/n2715 ),
    .b(1'b1),
    .c(\u2_Display/add86/c17 ),
    .o({\u2_Display/add86/c18 ,\u2_Display/n2735 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u18  (
    .a(\u2_Display/n2714 ),
    .b(1'b1),
    .c(\u2_Display/add86/c18 ),
    .o({\u2_Display/add86/c19 ,\u2_Display/n2735 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u19  (
    .a(\u2_Display/n2713 ),
    .b(1'b1),
    .c(\u2_Display/add86/c19 ),
    .o({\u2_Display/add86/c20 ,\u2_Display/n2735 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u2  (
    .a(\u2_Display/n2730 ),
    .b(1'b1),
    .c(\u2_Display/add86/c2 ),
    .o({\u2_Display/add86/c3 ,\u2_Display/n2735 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u20  (
    .a(\u2_Display/n2712 ),
    .b(1'b1),
    .c(\u2_Display/add86/c20 ),
    .o({\u2_Display/add86/c21 ,\u2_Display/n2735 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u21  (
    .a(\u2_Display/n2711 ),
    .b(1'b1),
    .c(\u2_Display/add86/c21 ),
    .o({\u2_Display/add86/c22 ,\u2_Display/n2735 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u22  (
    .a(\u2_Display/n2710 ),
    .b(1'b1),
    .c(\u2_Display/add86/c22 ),
    .o({\u2_Display/add86/c23 ,\u2_Display/n2735 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u23  (
    .a(\u2_Display/n2709 ),
    .b(1'b0),
    .c(\u2_Display/add86/c23 ),
    .o({\u2_Display/add86/c24 ,\u2_Display/n2735 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u24  (
    .a(\u2_Display/n2708 ),
    .b(1'b0),
    .c(\u2_Display/add86/c24 ),
    .o({\u2_Display/add86/c25 ,\u2_Display/n2735 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u25  (
    .a(\u2_Display/n2707 ),
    .b(1'b1),
    .c(\u2_Display/add86/c25 ),
    .o({\u2_Display/add86/c26 ,\u2_Display/n2735 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u26  (
    .a(\u2_Display/n2706 ),
    .b(1'b0),
    .c(\u2_Display/add86/c26 ),
    .o({\u2_Display/add86/c27 ,\u2_Display/n2735 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u27  (
    .a(\u2_Display/n2705 ),
    .b(1'b1),
    .c(\u2_Display/add86/c27 ),
    .o({\u2_Display/add86/c28 ,\u2_Display/n2735 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u28  (
    .a(\u2_Display/n2704 ),
    .b(1'b1),
    .c(\u2_Display/add86/c28 ),
    .o({\u2_Display/add86/c29 ,\u2_Display/n2735 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u29  (
    .a(\u2_Display/n2703 ),
    .b(1'b0),
    .c(\u2_Display/add86/c29 ),
    .o({\u2_Display/add86/c30 ,\u2_Display/n2735 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u3  (
    .a(\u2_Display/n2729 ),
    .b(1'b1),
    .c(\u2_Display/add86/c3 ),
    .o({\u2_Display/add86/c4 ,\u2_Display/n2735 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u30  (
    .a(\u2_Display/n2702 ),
    .b(1'b1),
    .c(\u2_Display/add86/c30 ),
    .o({\u2_Display/add86/c31 ,\u2_Display/n2735 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u31  (
    .a(\u2_Display/n2701 ),
    .b(1'b1),
    .c(\u2_Display/add86/c31 ),
    .o({open_n1301,\u2_Display/n2735 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u4  (
    .a(\u2_Display/n2728 ),
    .b(1'b1),
    .c(\u2_Display/add86/c4 ),
    .o({\u2_Display/add86/c5 ,\u2_Display/n2735 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u5  (
    .a(\u2_Display/n2727 ),
    .b(1'b1),
    .c(\u2_Display/add86/c5 ),
    .o({\u2_Display/add86/c6 ,\u2_Display/n2735 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u6  (
    .a(\u2_Display/n2726 ),
    .b(1'b1),
    .c(\u2_Display/add86/c6 ),
    .o({\u2_Display/add86/c7 ,\u2_Display/n2735 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u7  (
    .a(\u2_Display/n2725 ),
    .b(1'b1),
    .c(\u2_Display/add86/c7 ),
    .o({\u2_Display/add86/c8 ,\u2_Display/n2735 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u8  (
    .a(\u2_Display/n2724 ),
    .b(1'b1),
    .c(\u2_Display/add86/c8 ),
    .o({\u2_Display/add86/c9 ,\u2_Display/n2735 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add86/u9  (
    .a(\u2_Display/n2723 ),
    .b(1'b1),
    .c(\u2_Display/add86/c9 ),
    .o({\u2_Display/add86/c10 ,\u2_Display/n2735 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add86/ucin  (
    .a(1'b1),
    .o({\u2_Display/add86/c0 ,open_n1304}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u0  (
    .a(\u2_Display/n2767 ),
    .b(1'b1),
    .c(\u2_Display/add87/c0 ),
    .o({\u2_Display/add87/c1 ,\u2_Display/n2770 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u1  (
    .a(\u2_Display/n2766 ),
    .b(1'b1),
    .c(\u2_Display/add87/c1 ),
    .o({\u2_Display/add87/c2 ,\u2_Display/n2770 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u10  (
    .a(\u2_Display/n2757 ),
    .b(1'b1),
    .c(\u2_Display/add87/c10 ),
    .o({\u2_Display/add87/c11 ,\u2_Display/n2770 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u11  (
    .a(\u2_Display/n2756 ),
    .b(1'b1),
    .c(\u2_Display/add87/c11 ),
    .o({\u2_Display/add87/c12 ,\u2_Display/n2770 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u12  (
    .a(\u2_Display/n2755 ),
    .b(1'b1),
    .c(\u2_Display/add87/c12 ),
    .o({\u2_Display/add87/c13 ,\u2_Display/n2770 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u13  (
    .a(\u2_Display/n2754 ),
    .b(1'b1),
    .c(\u2_Display/add87/c13 ),
    .o({\u2_Display/add87/c14 ,\u2_Display/n2770 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u14  (
    .a(\u2_Display/n2753 ),
    .b(1'b1),
    .c(\u2_Display/add87/c14 ),
    .o({\u2_Display/add87/c15 ,\u2_Display/n2770 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u15  (
    .a(\u2_Display/n2752 ),
    .b(1'b1),
    .c(\u2_Display/add87/c15 ),
    .o({\u2_Display/add87/c16 ,\u2_Display/n2770 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u16  (
    .a(\u2_Display/n2751 ),
    .b(1'b1),
    .c(\u2_Display/add87/c16 ),
    .o({\u2_Display/add87/c17 ,\u2_Display/n2770 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u17  (
    .a(\u2_Display/n2750 ),
    .b(1'b1),
    .c(\u2_Display/add87/c17 ),
    .o({\u2_Display/add87/c18 ,\u2_Display/n2770 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u18  (
    .a(\u2_Display/n2749 ),
    .b(1'b1),
    .c(\u2_Display/add87/c18 ),
    .o({\u2_Display/add87/c19 ,\u2_Display/n2770 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u19  (
    .a(\u2_Display/n2748 ),
    .b(1'b1),
    .c(\u2_Display/add87/c19 ),
    .o({\u2_Display/add87/c20 ,\u2_Display/n2770 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u2  (
    .a(\u2_Display/n2765 ),
    .b(1'b1),
    .c(\u2_Display/add87/c2 ),
    .o({\u2_Display/add87/c3 ,\u2_Display/n2770 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u20  (
    .a(\u2_Display/n2747 ),
    .b(1'b1),
    .c(\u2_Display/add87/c20 ),
    .o({\u2_Display/add87/c21 ,\u2_Display/n2770 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u21  (
    .a(\u2_Display/n2746 ),
    .b(1'b1),
    .c(\u2_Display/add87/c21 ),
    .o({\u2_Display/add87/c22 ,\u2_Display/n2770 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u22  (
    .a(\u2_Display/n2745 ),
    .b(1'b0),
    .c(\u2_Display/add87/c22 ),
    .o({\u2_Display/add87/c23 ,\u2_Display/n2770 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u23  (
    .a(\u2_Display/n2744 ),
    .b(1'b0),
    .c(\u2_Display/add87/c23 ),
    .o({\u2_Display/add87/c24 ,\u2_Display/n2770 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u24  (
    .a(\u2_Display/n2743 ),
    .b(1'b1),
    .c(\u2_Display/add87/c24 ),
    .o({\u2_Display/add87/c25 ,\u2_Display/n2770 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u25  (
    .a(\u2_Display/n2742 ),
    .b(1'b0),
    .c(\u2_Display/add87/c25 ),
    .o({\u2_Display/add87/c26 ,\u2_Display/n2770 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u26  (
    .a(\u2_Display/n2741 ),
    .b(1'b1),
    .c(\u2_Display/add87/c26 ),
    .o({\u2_Display/add87/c27 ,\u2_Display/n2770 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u27  (
    .a(\u2_Display/n2740 ),
    .b(1'b1),
    .c(\u2_Display/add87/c27 ),
    .o({\u2_Display/add87/c28 ,\u2_Display/n2770 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u28  (
    .a(\u2_Display/n2739 ),
    .b(1'b0),
    .c(\u2_Display/add87/c28 ),
    .o({\u2_Display/add87/c29 ,\u2_Display/n2770 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u29  (
    .a(\u2_Display/n2738 ),
    .b(1'b1),
    .c(\u2_Display/add87/c29 ),
    .o({\u2_Display/add87/c30 ,\u2_Display/n2770 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u3  (
    .a(\u2_Display/n2764 ),
    .b(1'b1),
    .c(\u2_Display/add87/c3 ),
    .o({\u2_Display/add87/c4 ,\u2_Display/n2770 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u30  (
    .a(\u2_Display/n2737 ),
    .b(1'b1),
    .c(\u2_Display/add87/c30 ),
    .o({\u2_Display/add87/c31 ,\u2_Display/n2770 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u31  (
    .a(\u2_Display/n2736 ),
    .b(1'b1),
    .c(\u2_Display/add87/c31 ),
    .o({open_n1305,\u2_Display/n2770 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u4  (
    .a(\u2_Display/n2763 ),
    .b(1'b1),
    .c(\u2_Display/add87/c4 ),
    .o({\u2_Display/add87/c5 ,\u2_Display/n2770 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u5  (
    .a(\u2_Display/n2762 ),
    .b(1'b1),
    .c(\u2_Display/add87/c5 ),
    .o({\u2_Display/add87/c6 ,\u2_Display/n2770 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u6  (
    .a(\u2_Display/n2761 ),
    .b(1'b1),
    .c(\u2_Display/add87/c6 ),
    .o({\u2_Display/add87/c7 ,\u2_Display/n2770 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u7  (
    .a(\u2_Display/n2760 ),
    .b(1'b1),
    .c(\u2_Display/add87/c7 ),
    .o({\u2_Display/add87/c8 ,\u2_Display/n2770 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u8  (
    .a(\u2_Display/n2759 ),
    .b(1'b1),
    .c(\u2_Display/add87/c8 ),
    .o({\u2_Display/add87/c9 ,\u2_Display/n2770 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add87/u9  (
    .a(\u2_Display/n2758 ),
    .b(1'b1),
    .c(\u2_Display/add87/c9 ),
    .o({\u2_Display/add87/c10 ,\u2_Display/n2770 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add87/ucin  (
    .a(1'b1),
    .o({\u2_Display/add87/c0 ,open_n1308}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u0  (
    .a(\u2_Display/n2802 ),
    .b(1'b1),
    .c(\u2_Display/add88/c0 ),
    .o({\u2_Display/add88/c1 ,\u2_Display/n2805 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u1  (
    .a(\u2_Display/n2801 ),
    .b(1'b1),
    .c(\u2_Display/add88/c1 ),
    .o({\u2_Display/add88/c2 ,\u2_Display/n2805 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u10  (
    .a(\u2_Display/n2792 ),
    .b(1'b1),
    .c(\u2_Display/add88/c10 ),
    .o({\u2_Display/add88/c11 ,\u2_Display/n2805 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u11  (
    .a(\u2_Display/n2791 ),
    .b(1'b1),
    .c(\u2_Display/add88/c11 ),
    .o({\u2_Display/add88/c12 ,\u2_Display/n2805 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u12  (
    .a(\u2_Display/n2790 ),
    .b(1'b1),
    .c(\u2_Display/add88/c12 ),
    .o({\u2_Display/add88/c13 ,\u2_Display/n2805 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u13  (
    .a(\u2_Display/n2789 ),
    .b(1'b1),
    .c(\u2_Display/add88/c13 ),
    .o({\u2_Display/add88/c14 ,\u2_Display/n2805 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u14  (
    .a(\u2_Display/n2788 ),
    .b(1'b1),
    .c(\u2_Display/add88/c14 ),
    .o({\u2_Display/add88/c15 ,\u2_Display/n2805 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u15  (
    .a(\u2_Display/n2787 ),
    .b(1'b1),
    .c(\u2_Display/add88/c15 ),
    .o({\u2_Display/add88/c16 ,\u2_Display/n2805 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u16  (
    .a(\u2_Display/n2786 ),
    .b(1'b1),
    .c(\u2_Display/add88/c16 ),
    .o({\u2_Display/add88/c17 ,\u2_Display/n2805 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u17  (
    .a(\u2_Display/n2785 ),
    .b(1'b1),
    .c(\u2_Display/add88/c17 ),
    .o({\u2_Display/add88/c18 ,\u2_Display/n2805 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u18  (
    .a(\u2_Display/n2784 ),
    .b(1'b1),
    .c(\u2_Display/add88/c18 ),
    .o({\u2_Display/add88/c19 ,\u2_Display/n2805 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u19  (
    .a(\u2_Display/n2783 ),
    .b(1'b1),
    .c(\u2_Display/add88/c19 ),
    .o({\u2_Display/add88/c20 ,\u2_Display/n2805 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u2  (
    .a(\u2_Display/n2800 ),
    .b(1'b1),
    .c(\u2_Display/add88/c2 ),
    .o({\u2_Display/add88/c3 ,\u2_Display/n2805 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u20  (
    .a(\u2_Display/n2782 ),
    .b(1'b1),
    .c(\u2_Display/add88/c20 ),
    .o({\u2_Display/add88/c21 ,\u2_Display/n2805 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u21  (
    .a(\u2_Display/n2781 ),
    .b(1'b0),
    .c(\u2_Display/add88/c21 ),
    .o({\u2_Display/add88/c22 ,\u2_Display/n2805 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u22  (
    .a(\u2_Display/n2780 ),
    .b(1'b0),
    .c(\u2_Display/add88/c22 ),
    .o({\u2_Display/add88/c23 ,\u2_Display/n2805 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u23  (
    .a(\u2_Display/n2779 ),
    .b(1'b1),
    .c(\u2_Display/add88/c23 ),
    .o({\u2_Display/add88/c24 ,\u2_Display/n2805 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u24  (
    .a(\u2_Display/n2778 ),
    .b(1'b0),
    .c(\u2_Display/add88/c24 ),
    .o({\u2_Display/add88/c25 ,\u2_Display/n2805 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u25  (
    .a(\u2_Display/n2777 ),
    .b(1'b1),
    .c(\u2_Display/add88/c25 ),
    .o({\u2_Display/add88/c26 ,\u2_Display/n2805 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u26  (
    .a(\u2_Display/n2776 ),
    .b(1'b1),
    .c(\u2_Display/add88/c26 ),
    .o({\u2_Display/add88/c27 ,\u2_Display/n2805 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u27  (
    .a(\u2_Display/n2775 ),
    .b(1'b0),
    .c(\u2_Display/add88/c27 ),
    .o({\u2_Display/add88/c28 ,\u2_Display/n2805 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u28  (
    .a(\u2_Display/n2774 ),
    .b(1'b1),
    .c(\u2_Display/add88/c28 ),
    .o({\u2_Display/add88/c29 ,\u2_Display/n2805 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u29  (
    .a(\u2_Display/n2773 ),
    .b(1'b1),
    .c(\u2_Display/add88/c29 ),
    .o({\u2_Display/add88/c30 ,\u2_Display/n2805 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u3  (
    .a(\u2_Display/n2799 ),
    .b(1'b1),
    .c(\u2_Display/add88/c3 ),
    .o({\u2_Display/add88/c4 ,\u2_Display/n2805 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u30  (
    .a(\u2_Display/n2772 ),
    .b(1'b1),
    .c(\u2_Display/add88/c30 ),
    .o({\u2_Display/add88/c31 ,\u2_Display/n2805 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u31  (
    .a(\u2_Display/n2771 ),
    .b(1'b1),
    .c(\u2_Display/add88/c31 ),
    .o({open_n1309,\u2_Display/n2805 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u4  (
    .a(\u2_Display/n2798 ),
    .b(1'b1),
    .c(\u2_Display/add88/c4 ),
    .o({\u2_Display/add88/c5 ,\u2_Display/n2805 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u5  (
    .a(\u2_Display/n2797 ),
    .b(1'b1),
    .c(\u2_Display/add88/c5 ),
    .o({\u2_Display/add88/c6 ,\u2_Display/n2805 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u6  (
    .a(\u2_Display/n2796 ),
    .b(1'b1),
    .c(\u2_Display/add88/c6 ),
    .o({\u2_Display/add88/c7 ,\u2_Display/n2805 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u7  (
    .a(\u2_Display/n2795 ),
    .b(1'b1),
    .c(\u2_Display/add88/c7 ),
    .o({\u2_Display/add88/c8 ,\u2_Display/n2805 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u8  (
    .a(\u2_Display/n2794 ),
    .b(1'b1),
    .c(\u2_Display/add88/c8 ),
    .o({\u2_Display/add88/c9 ,\u2_Display/n2805 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add88/u9  (
    .a(\u2_Display/n2793 ),
    .b(1'b1),
    .c(\u2_Display/add88/c9 ),
    .o({\u2_Display/add88/c10 ,\u2_Display/n2805 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add88/ucin  (
    .a(1'b1),
    .o({\u2_Display/add88/c0 ,open_n1312}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u0  (
    .a(\u2_Display/n2837 ),
    .b(1'b1),
    .c(\u2_Display/add89/c0 ),
    .o({\u2_Display/add89/c1 ,\u2_Display/n2840 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u1  (
    .a(\u2_Display/n2836 ),
    .b(1'b1),
    .c(\u2_Display/add89/c1 ),
    .o({\u2_Display/add89/c2 ,\u2_Display/n2840 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u10  (
    .a(\u2_Display/n2827 ),
    .b(1'b1),
    .c(\u2_Display/add89/c10 ),
    .o({\u2_Display/add89/c11 ,\u2_Display/n2840 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u11  (
    .a(\u2_Display/n2826 ),
    .b(1'b1),
    .c(\u2_Display/add89/c11 ),
    .o({\u2_Display/add89/c12 ,\u2_Display/n2840 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u12  (
    .a(\u2_Display/n2825 ),
    .b(1'b1),
    .c(\u2_Display/add89/c12 ),
    .o({\u2_Display/add89/c13 ,\u2_Display/n2840 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u13  (
    .a(\u2_Display/n2824 ),
    .b(1'b1),
    .c(\u2_Display/add89/c13 ),
    .o({\u2_Display/add89/c14 ,\u2_Display/n2840 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u14  (
    .a(\u2_Display/n2823 ),
    .b(1'b1),
    .c(\u2_Display/add89/c14 ),
    .o({\u2_Display/add89/c15 ,\u2_Display/n2840 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u15  (
    .a(\u2_Display/n2822 ),
    .b(1'b1),
    .c(\u2_Display/add89/c15 ),
    .o({\u2_Display/add89/c16 ,\u2_Display/n2840 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u16  (
    .a(\u2_Display/n2821 ),
    .b(1'b1),
    .c(\u2_Display/add89/c16 ),
    .o({\u2_Display/add89/c17 ,\u2_Display/n2840 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u17  (
    .a(\u2_Display/n2820 ),
    .b(1'b1),
    .c(\u2_Display/add89/c17 ),
    .o({\u2_Display/add89/c18 ,\u2_Display/n2840 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u18  (
    .a(\u2_Display/n2819 ),
    .b(1'b1),
    .c(\u2_Display/add89/c18 ),
    .o({\u2_Display/add89/c19 ,\u2_Display/n2840 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u19  (
    .a(\u2_Display/n2818 ),
    .b(1'b1),
    .c(\u2_Display/add89/c19 ),
    .o({\u2_Display/add89/c20 ,\u2_Display/n2840 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u2  (
    .a(\u2_Display/n2835 ),
    .b(1'b1),
    .c(\u2_Display/add89/c2 ),
    .o({\u2_Display/add89/c3 ,\u2_Display/n2840 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u20  (
    .a(\u2_Display/n2817 ),
    .b(1'b0),
    .c(\u2_Display/add89/c20 ),
    .o({\u2_Display/add89/c21 ,\u2_Display/n2840 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u21  (
    .a(\u2_Display/n2816 ),
    .b(1'b0),
    .c(\u2_Display/add89/c21 ),
    .o({\u2_Display/add89/c22 ,\u2_Display/n2840 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u22  (
    .a(\u2_Display/n2815 ),
    .b(1'b1),
    .c(\u2_Display/add89/c22 ),
    .o({\u2_Display/add89/c23 ,\u2_Display/n2840 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u23  (
    .a(\u2_Display/n2814 ),
    .b(1'b0),
    .c(\u2_Display/add89/c23 ),
    .o({\u2_Display/add89/c24 ,\u2_Display/n2840 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u24  (
    .a(\u2_Display/n2813 ),
    .b(1'b1),
    .c(\u2_Display/add89/c24 ),
    .o({\u2_Display/add89/c25 ,\u2_Display/n2840 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u25  (
    .a(\u2_Display/n2812 ),
    .b(1'b1),
    .c(\u2_Display/add89/c25 ),
    .o({\u2_Display/add89/c26 ,\u2_Display/n2840 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u26  (
    .a(\u2_Display/n2811 ),
    .b(1'b0),
    .c(\u2_Display/add89/c26 ),
    .o({\u2_Display/add89/c27 ,\u2_Display/n2840 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u27  (
    .a(\u2_Display/n2810 ),
    .b(1'b1),
    .c(\u2_Display/add89/c27 ),
    .o({\u2_Display/add89/c28 ,\u2_Display/n2840 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u28  (
    .a(\u2_Display/n2809 ),
    .b(1'b1),
    .c(\u2_Display/add89/c28 ),
    .o({\u2_Display/add89/c29 ,\u2_Display/n2840 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u29  (
    .a(\u2_Display/n2808 ),
    .b(1'b1),
    .c(\u2_Display/add89/c29 ),
    .o({\u2_Display/add89/c30 ,\u2_Display/n2840 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u3  (
    .a(\u2_Display/n2834 ),
    .b(1'b1),
    .c(\u2_Display/add89/c3 ),
    .o({\u2_Display/add89/c4 ,\u2_Display/n2840 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u30  (
    .a(\u2_Display/n2807 ),
    .b(1'b1),
    .c(\u2_Display/add89/c30 ),
    .o({\u2_Display/add89/c31 ,\u2_Display/n2840 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u31  (
    .a(\u2_Display/n2806 ),
    .b(1'b1),
    .c(\u2_Display/add89/c31 ),
    .o({open_n1313,\u2_Display/n2840 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u4  (
    .a(\u2_Display/n2833 ),
    .b(1'b1),
    .c(\u2_Display/add89/c4 ),
    .o({\u2_Display/add89/c5 ,\u2_Display/n2840 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u5  (
    .a(\u2_Display/n2832 ),
    .b(1'b1),
    .c(\u2_Display/add89/c5 ),
    .o({\u2_Display/add89/c6 ,\u2_Display/n2840 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u6  (
    .a(\u2_Display/n2831 ),
    .b(1'b1),
    .c(\u2_Display/add89/c6 ),
    .o({\u2_Display/add89/c7 ,\u2_Display/n2840 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u7  (
    .a(\u2_Display/n2830 ),
    .b(1'b1),
    .c(\u2_Display/add89/c7 ),
    .o({\u2_Display/add89/c8 ,\u2_Display/n2840 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u8  (
    .a(\u2_Display/n2829 ),
    .b(1'b1),
    .c(\u2_Display/add89/c8 ),
    .o({\u2_Display/add89/c9 ,\u2_Display/n2840 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add89/u9  (
    .a(\u2_Display/n2828 ),
    .b(1'b1),
    .c(\u2_Display/add89/c9 ),
    .o({\u2_Display/add89/c10 ,\u2_Display/n2840 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add89/ucin  (
    .a(1'b1),
    .o({\u2_Display/add89/c0 ,open_n1316}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u0  (
    .a(\u2_Display/n2872 ),
    .b(1'b1),
    .c(\u2_Display/add90/c0 ),
    .o({\u2_Display/add90/c1 ,\u2_Display/n2875 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u1  (
    .a(\u2_Display/n2871 ),
    .b(1'b1),
    .c(\u2_Display/add90/c1 ),
    .o({\u2_Display/add90/c2 ,\u2_Display/n2875 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u10  (
    .a(\u2_Display/n2862 ),
    .b(1'b1),
    .c(\u2_Display/add90/c10 ),
    .o({\u2_Display/add90/c11 ,\u2_Display/n2875 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u11  (
    .a(\u2_Display/n2861 ),
    .b(1'b1),
    .c(\u2_Display/add90/c11 ),
    .o({\u2_Display/add90/c12 ,\u2_Display/n2875 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u12  (
    .a(\u2_Display/n2860 ),
    .b(1'b1),
    .c(\u2_Display/add90/c12 ),
    .o({\u2_Display/add90/c13 ,\u2_Display/n2875 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u13  (
    .a(\u2_Display/n2859 ),
    .b(1'b1),
    .c(\u2_Display/add90/c13 ),
    .o({\u2_Display/add90/c14 ,\u2_Display/n2875 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u14  (
    .a(\u2_Display/n2858 ),
    .b(1'b1),
    .c(\u2_Display/add90/c14 ),
    .o({\u2_Display/add90/c15 ,\u2_Display/n2875 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u15  (
    .a(\u2_Display/n2857 ),
    .b(1'b1),
    .c(\u2_Display/add90/c15 ),
    .o({\u2_Display/add90/c16 ,\u2_Display/n2875 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u16  (
    .a(\u2_Display/n2856 ),
    .b(1'b1),
    .c(\u2_Display/add90/c16 ),
    .o({\u2_Display/add90/c17 ,\u2_Display/n2875 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u17  (
    .a(\u2_Display/n2855 ),
    .b(1'b1),
    .c(\u2_Display/add90/c17 ),
    .o({\u2_Display/add90/c18 ,\u2_Display/n2875 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u18  (
    .a(\u2_Display/n2854 ),
    .b(1'b1),
    .c(\u2_Display/add90/c18 ),
    .o({\u2_Display/add90/c19 ,\u2_Display/n2875 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u19  (
    .a(\u2_Display/n2853 ),
    .b(1'b0),
    .c(\u2_Display/add90/c19 ),
    .o({\u2_Display/add90/c20 ,\u2_Display/n2875 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u2  (
    .a(\u2_Display/n2870 ),
    .b(1'b1),
    .c(\u2_Display/add90/c2 ),
    .o({\u2_Display/add90/c3 ,\u2_Display/n2875 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u20  (
    .a(\u2_Display/n2852 ),
    .b(1'b0),
    .c(\u2_Display/add90/c20 ),
    .o({\u2_Display/add90/c21 ,\u2_Display/n2875 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u21  (
    .a(\u2_Display/n2851 ),
    .b(1'b1),
    .c(\u2_Display/add90/c21 ),
    .o({\u2_Display/add90/c22 ,\u2_Display/n2875 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u22  (
    .a(\u2_Display/n2850 ),
    .b(1'b0),
    .c(\u2_Display/add90/c22 ),
    .o({\u2_Display/add90/c23 ,\u2_Display/n2875 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u23  (
    .a(\u2_Display/n2849 ),
    .b(1'b1),
    .c(\u2_Display/add90/c23 ),
    .o({\u2_Display/add90/c24 ,\u2_Display/n2875 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u24  (
    .a(\u2_Display/n2848 ),
    .b(1'b1),
    .c(\u2_Display/add90/c24 ),
    .o({\u2_Display/add90/c25 ,\u2_Display/n2875 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u25  (
    .a(\u2_Display/n2847 ),
    .b(1'b0),
    .c(\u2_Display/add90/c25 ),
    .o({\u2_Display/add90/c26 ,\u2_Display/n2875 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u26  (
    .a(\u2_Display/n2846 ),
    .b(1'b1),
    .c(\u2_Display/add90/c26 ),
    .o({\u2_Display/add90/c27 ,\u2_Display/n2875 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u27  (
    .a(\u2_Display/n2845 ),
    .b(1'b1),
    .c(\u2_Display/add90/c27 ),
    .o({\u2_Display/add90/c28 ,\u2_Display/n2875 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u28  (
    .a(\u2_Display/n2844 ),
    .b(1'b1),
    .c(\u2_Display/add90/c28 ),
    .o({\u2_Display/add90/c29 ,\u2_Display/n2875 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u29  (
    .a(\u2_Display/n2843 ),
    .b(1'b1),
    .c(\u2_Display/add90/c29 ),
    .o({\u2_Display/add90/c30 ,\u2_Display/n2875 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u3  (
    .a(\u2_Display/n2869 ),
    .b(1'b1),
    .c(\u2_Display/add90/c3 ),
    .o({\u2_Display/add90/c4 ,\u2_Display/n2875 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u30  (
    .a(\u2_Display/n2842 ),
    .b(1'b1),
    .c(\u2_Display/add90/c30 ),
    .o({\u2_Display/add90/c31 ,\u2_Display/n2875 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u31  (
    .a(\u2_Display/n2841 ),
    .b(1'b1),
    .c(\u2_Display/add90/c31 ),
    .o({open_n1317,\u2_Display/n2875 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u4  (
    .a(\u2_Display/n2868 ),
    .b(1'b1),
    .c(\u2_Display/add90/c4 ),
    .o({\u2_Display/add90/c5 ,\u2_Display/n2875 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u5  (
    .a(\u2_Display/n2867 ),
    .b(1'b1),
    .c(\u2_Display/add90/c5 ),
    .o({\u2_Display/add90/c6 ,\u2_Display/n2875 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u6  (
    .a(\u2_Display/n2866 ),
    .b(1'b1),
    .c(\u2_Display/add90/c6 ),
    .o({\u2_Display/add90/c7 ,\u2_Display/n2875 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u7  (
    .a(\u2_Display/n2865 ),
    .b(1'b1),
    .c(\u2_Display/add90/c7 ),
    .o({\u2_Display/add90/c8 ,\u2_Display/n2875 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u8  (
    .a(\u2_Display/n2864 ),
    .b(1'b1),
    .c(\u2_Display/add90/c8 ),
    .o({\u2_Display/add90/c9 ,\u2_Display/n2875 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add90/u9  (
    .a(\u2_Display/n2863 ),
    .b(1'b1),
    .c(\u2_Display/add90/c9 ),
    .o({\u2_Display/add90/c10 ,\u2_Display/n2875 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add90/ucin  (
    .a(1'b1),
    .o({\u2_Display/add90/c0 ,open_n1320}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u0  (
    .a(\u2_Display/n2907 ),
    .b(1'b1),
    .c(\u2_Display/add91/c0 ),
    .o({\u2_Display/add91/c1 ,\u2_Display/n2910 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u1  (
    .a(\u2_Display/n2906 ),
    .b(1'b1),
    .c(\u2_Display/add91/c1 ),
    .o({\u2_Display/add91/c2 ,\u2_Display/n2910 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u10  (
    .a(\u2_Display/n2897 ),
    .b(1'b1),
    .c(\u2_Display/add91/c10 ),
    .o({\u2_Display/add91/c11 ,\u2_Display/n2910 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u11  (
    .a(\u2_Display/n2896 ),
    .b(1'b1),
    .c(\u2_Display/add91/c11 ),
    .o({\u2_Display/add91/c12 ,\u2_Display/n2910 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u12  (
    .a(\u2_Display/n2895 ),
    .b(1'b1),
    .c(\u2_Display/add91/c12 ),
    .o({\u2_Display/add91/c13 ,\u2_Display/n2910 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u13  (
    .a(\u2_Display/n2894 ),
    .b(1'b1),
    .c(\u2_Display/add91/c13 ),
    .o({\u2_Display/add91/c14 ,\u2_Display/n2910 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u14  (
    .a(\u2_Display/n2893 ),
    .b(1'b1),
    .c(\u2_Display/add91/c14 ),
    .o({\u2_Display/add91/c15 ,\u2_Display/n2910 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u15  (
    .a(\u2_Display/n2892 ),
    .b(1'b1),
    .c(\u2_Display/add91/c15 ),
    .o({\u2_Display/add91/c16 ,\u2_Display/n2910 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u16  (
    .a(\u2_Display/n2891 ),
    .b(1'b1),
    .c(\u2_Display/add91/c16 ),
    .o({\u2_Display/add91/c17 ,\u2_Display/n2910 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u17  (
    .a(\u2_Display/n2890 ),
    .b(1'b1),
    .c(\u2_Display/add91/c17 ),
    .o({\u2_Display/add91/c18 ,\u2_Display/n2910 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u18  (
    .a(\u2_Display/n2889 ),
    .b(1'b0),
    .c(\u2_Display/add91/c18 ),
    .o({\u2_Display/add91/c19 ,\u2_Display/n2910 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u19  (
    .a(\u2_Display/n2888 ),
    .b(1'b0),
    .c(\u2_Display/add91/c19 ),
    .o({\u2_Display/add91/c20 ,\u2_Display/n2910 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u2  (
    .a(\u2_Display/n2905 ),
    .b(1'b1),
    .c(\u2_Display/add91/c2 ),
    .o({\u2_Display/add91/c3 ,\u2_Display/n2910 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u20  (
    .a(\u2_Display/n2887 ),
    .b(1'b1),
    .c(\u2_Display/add91/c20 ),
    .o({\u2_Display/add91/c21 ,\u2_Display/n2910 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u21  (
    .a(\u2_Display/n2886 ),
    .b(1'b0),
    .c(\u2_Display/add91/c21 ),
    .o({\u2_Display/add91/c22 ,\u2_Display/n2910 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u22  (
    .a(\u2_Display/n2885 ),
    .b(1'b1),
    .c(\u2_Display/add91/c22 ),
    .o({\u2_Display/add91/c23 ,\u2_Display/n2910 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u23  (
    .a(\u2_Display/n2884 ),
    .b(1'b1),
    .c(\u2_Display/add91/c23 ),
    .o({\u2_Display/add91/c24 ,\u2_Display/n2910 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u24  (
    .a(\u2_Display/n2883 ),
    .b(1'b0),
    .c(\u2_Display/add91/c24 ),
    .o({\u2_Display/add91/c25 ,\u2_Display/n2910 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u25  (
    .a(\u2_Display/n2882 ),
    .b(1'b1),
    .c(\u2_Display/add91/c25 ),
    .o({\u2_Display/add91/c26 ,\u2_Display/n2910 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u26  (
    .a(\u2_Display/n2881 ),
    .b(1'b1),
    .c(\u2_Display/add91/c26 ),
    .o({\u2_Display/add91/c27 ,\u2_Display/n2910 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u27  (
    .a(\u2_Display/n2880 ),
    .b(1'b1),
    .c(\u2_Display/add91/c27 ),
    .o({\u2_Display/add91/c28 ,\u2_Display/n2910 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u28  (
    .a(\u2_Display/n2879 ),
    .b(1'b1),
    .c(\u2_Display/add91/c28 ),
    .o({\u2_Display/add91/c29 ,\u2_Display/n2910 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u29  (
    .a(\u2_Display/n2878 ),
    .b(1'b1),
    .c(\u2_Display/add91/c29 ),
    .o({\u2_Display/add91/c30 ,\u2_Display/n2910 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u3  (
    .a(\u2_Display/n2904 ),
    .b(1'b1),
    .c(\u2_Display/add91/c3 ),
    .o({\u2_Display/add91/c4 ,\u2_Display/n2910 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u30  (
    .a(\u2_Display/n2877 ),
    .b(1'b1),
    .c(\u2_Display/add91/c30 ),
    .o({\u2_Display/add91/c31 ,\u2_Display/n2910 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u31  (
    .a(\u2_Display/n2876 ),
    .b(1'b1),
    .c(\u2_Display/add91/c31 ),
    .o({open_n1321,\u2_Display/n2910 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u4  (
    .a(\u2_Display/n2903 ),
    .b(1'b1),
    .c(\u2_Display/add91/c4 ),
    .o({\u2_Display/add91/c5 ,\u2_Display/n2910 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u5  (
    .a(\u2_Display/n2902 ),
    .b(1'b1),
    .c(\u2_Display/add91/c5 ),
    .o({\u2_Display/add91/c6 ,\u2_Display/n2910 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u6  (
    .a(\u2_Display/n2901 ),
    .b(1'b1),
    .c(\u2_Display/add91/c6 ),
    .o({\u2_Display/add91/c7 ,\u2_Display/n2910 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u7  (
    .a(\u2_Display/n2900 ),
    .b(1'b1),
    .c(\u2_Display/add91/c7 ),
    .o({\u2_Display/add91/c8 ,\u2_Display/n2910 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u8  (
    .a(\u2_Display/n2899 ),
    .b(1'b1),
    .c(\u2_Display/add91/c8 ),
    .o({\u2_Display/add91/c9 ,\u2_Display/n2910 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add91/u9  (
    .a(\u2_Display/n2898 ),
    .b(1'b1),
    .c(\u2_Display/add91/c9 ),
    .o({\u2_Display/add91/c10 ,\u2_Display/n2910 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add91/ucin  (
    .a(1'b1),
    .o({\u2_Display/add91/c0 ,open_n1324}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u0  (
    .a(\u2_Display/n2942 ),
    .b(1'b1),
    .c(\u2_Display/add92/c0 ),
    .o({\u2_Display/add92/c1 ,\u2_Display/n2945 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u1  (
    .a(\u2_Display/n2941 ),
    .b(1'b1),
    .c(\u2_Display/add92/c1 ),
    .o({\u2_Display/add92/c2 ,\u2_Display/n2945 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u10  (
    .a(\u2_Display/n2932 ),
    .b(1'b1),
    .c(\u2_Display/add92/c10 ),
    .o({\u2_Display/add92/c11 ,\u2_Display/n2945 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u11  (
    .a(\u2_Display/n2931 ),
    .b(1'b1),
    .c(\u2_Display/add92/c11 ),
    .o({\u2_Display/add92/c12 ,\u2_Display/n2945 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u12  (
    .a(\u2_Display/n2930 ),
    .b(1'b1),
    .c(\u2_Display/add92/c12 ),
    .o({\u2_Display/add92/c13 ,\u2_Display/n2945 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u13  (
    .a(\u2_Display/n2929 ),
    .b(1'b1),
    .c(\u2_Display/add92/c13 ),
    .o({\u2_Display/add92/c14 ,\u2_Display/n2945 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u14  (
    .a(\u2_Display/n2928 ),
    .b(1'b1),
    .c(\u2_Display/add92/c14 ),
    .o({\u2_Display/add92/c15 ,\u2_Display/n2945 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u15  (
    .a(\u2_Display/n2927 ),
    .b(1'b1),
    .c(\u2_Display/add92/c15 ),
    .o({\u2_Display/add92/c16 ,\u2_Display/n2945 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u16  (
    .a(\u2_Display/n2926 ),
    .b(1'b1),
    .c(\u2_Display/add92/c16 ),
    .o({\u2_Display/add92/c17 ,\u2_Display/n2945 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u17  (
    .a(\u2_Display/n2925 ),
    .b(1'b0),
    .c(\u2_Display/add92/c17 ),
    .o({\u2_Display/add92/c18 ,\u2_Display/n2945 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u18  (
    .a(\u2_Display/n2924 ),
    .b(1'b0),
    .c(\u2_Display/add92/c18 ),
    .o({\u2_Display/add92/c19 ,\u2_Display/n2945 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u19  (
    .a(\u2_Display/n2923 ),
    .b(1'b1),
    .c(\u2_Display/add92/c19 ),
    .o({\u2_Display/add92/c20 ,\u2_Display/n2945 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u2  (
    .a(\u2_Display/n2940 ),
    .b(1'b1),
    .c(\u2_Display/add92/c2 ),
    .o({\u2_Display/add92/c3 ,\u2_Display/n2945 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u20  (
    .a(\u2_Display/n2922 ),
    .b(1'b0),
    .c(\u2_Display/add92/c20 ),
    .o({\u2_Display/add92/c21 ,\u2_Display/n2945 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u21  (
    .a(\u2_Display/n2921 ),
    .b(1'b1),
    .c(\u2_Display/add92/c21 ),
    .o({\u2_Display/add92/c22 ,\u2_Display/n2945 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u22  (
    .a(\u2_Display/n2920 ),
    .b(1'b1),
    .c(\u2_Display/add92/c22 ),
    .o({\u2_Display/add92/c23 ,\u2_Display/n2945 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u23  (
    .a(\u2_Display/n2919 ),
    .b(1'b0),
    .c(\u2_Display/add92/c23 ),
    .o({\u2_Display/add92/c24 ,\u2_Display/n2945 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u24  (
    .a(\u2_Display/n2918 ),
    .b(1'b1),
    .c(\u2_Display/add92/c24 ),
    .o({\u2_Display/add92/c25 ,\u2_Display/n2945 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u25  (
    .a(\u2_Display/n2917 ),
    .b(1'b1),
    .c(\u2_Display/add92/c25 ),
    .o({\u2_Display/add92/c26 ,\u2_Display/n2945 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u26  (
    .a(\u2_Display/n2916 ),
    .b(1'b1),
    .c(\u2_Display/add92/c26 ),
    .o({\u2_Display/add92/c27 ,\u2_Display/n2945 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u27  (
    .a(\u2_Display/n2915 ),
    .b(1'b1),
    .c(\u2_Display/add92/c27 ),
    .o({\u2_Display/add92/c28 ,\u2_Display/n2945 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u28  (
    .a(\u2_Display/n2914 ),
    .b(1'b1),
    .c(\u2_Display/add92/c28 ),
    .o({\u2_Display/add92/c29 ,\u2_Display/n2945 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u29  (
    .a(\u2_Display/n2913 ),
    .b(1'b1),
    .c(\u2_Display/add92/c29 ),
    .o({\u2_Display/add92/c30 ,\u2_Display/n2945 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u3  (
    .a(\u2_Display/n2939 ),
    .b(1'b1),
    .c(\u2_Display/add92/c3 ),
    .o({\u2_Display/add92/c4 ,\u2_Display/n2945 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u30  (
    .a(\u2_Display/n2912 ),
    .b(1'b1),
    .c(\u2_Display/add92/c30 ),
    .o({\u2_Display/add92/c31 ,\u2_Display/n2945 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u31  (
    .a(\u2_Display/n2911 ),
    .b(1'b1),
    .c(\u2_Display/add92/c31 ),
    .o({open_n1325,\u2_Display/n2945 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u4  (
    .a(\u2_Display/n2938 ),
    .b(1'b1),
    .c(\u2_Display/add92/c4 ),
    .o({\u2_Display/add92/c5 ,\u2_Display/n2945 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u5  (
    .a(\u2_Display/n2937 ),
    .b(1'b1),
    .c(\u2_Display/add92/c5 ),
    .o({\u2_Display/add92/c6 ,\u2_Display/n2945 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u6  (
    .a(\u2_Display/n2936 ),
    .b(1'b1),
    .c(\u2_Display/add92/c6 ),
    .o({\u2_Display/add92/c7 ,\u2_Display/n2945 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u7  (
    .a(\u2_Display/n2935 ),
    .b(1'b1),
    .c(\u2_Display/add92/c7 ),
    .o({\u2_Display/add92/c8 ,\u2_Display/n2945 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u8  (
    .a(\u2_Display/n2934 ),
    .b(1'b1),
    .c(\u2_Display/add92/c8 ),
    .o({\u2_Display/add92/c9 ,\u2_Display/n2945 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add92/u9  (
    .a(\u2_Display/n2933 ),
    .b(1'b1),
    .c(\u2_Display/add92/c9 ),
    .o({\u2_Display/add92/c10 ,\u2_Display/n2945 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add92/ucin  (
    .a(1'b1),
    .o({\u2_Display/add92/c0 ,open_n1328}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u0  (
    .a(\u2_Display/n2977 ),
    .b(1'b1),
    .c(\u2_Display/add93/c0 ),
    .o({\u2_Display/add93/c1 ,\u2_Display/n2980 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u1  (
    .a(\u2_Display/n2976 ),
    .b(1'b1),
    .c(\u2_Display/add93/c1 ),
    .o({\u2_Display/add93/c2 ,\u2_Display/n2980 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u10  (
    .a(\u2_Display/n2967 ),
    .b(1'b1),
    .c(\u2_Display/add93/c10 ),
    .o({\u2_Display/add93/c11 ,\u2_Display/n2980 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u11  (
    .a(\u2_Display/n2966 ),
    .b(1'b1),
    .c(\u2_Display/add93/c11 ),
    .o({\u2_Display/add93/c12 ,\u2_Display/n2980 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u12  (
    .a(\u2_Display/n2965 ),
    .b(1'b1),
    .c(\u2_Display/add93/c12 ),
    .o({\u2_Display/add93/c13 ,\u2_Display/n2980 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u13  (
    .a(\u2_Display/n2964 ),
    .b(1'b1),
    .c(\u2_Display/add93/c13 ),
    .o({\u2_Display/add93/c14 ,\u2_Display/n2980 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u14  (
    .a(\u2_Display/n2963 ),
    .b(1'b1),
    .c(\u2_Display/add93/c14 ),
    .o({\u2_Display/add93/c15 ,\u2_Display/n2980 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u15  (
    .a(\u2_Display/n2962 ),
    .b(1'b1),
    .c(\u2_Display/add93/c15 ),
    .o({\u2_Display/add93/c16 ,\u2_Display/n2980 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u16  (
    .a(\u2_Display/n2961 ),
    .b(1'b0),
    .c(\u2_Display/add93/c16 ),
    .o({\u2_Display/add93/c17 ,\u2_Display/n2980 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u17  (
    .a(\u2_Display/n2960 ),
    .b(1'b0),
    .c(\u2_Display/add93/c17 ),
    .o({\u2_Display/add93/c18 ,\u2_Display/n2980 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u18  (
    .a(\u2_Display/n2959 ),
    .b(1'b1),
    .c(\u2_Display/add93/c18 ),
    .o({\u2_Display/add93/c19 ,\u2_Display/n2980 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u19  (
    .a(\u2_Display/n2958 ),
    .b(1'b0),
    .c(\u2_Display/add93/c19 ),
    .o({\u2_Display/add93/c20 ,\u2_Display/n2980 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u2  (
    .a(\u2_Display/n2975 ),
    .b(1'b1),
    .c(\u2_Display/add93/c2 ),
    .o({\u2_Display/add93/c3 ,\u2_Display/n2980 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u20  (
    .a(\u2_Display/n2957 ),
    .b(1'b1),
    .c(\u2_Display/add93/c20 ),
    .o({\u2_Display/add93/c21 ,\u2_Display/n2980 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u21  (
    .a(\u2_Display/n2956 ),
    .b(1'b1),
    .c(\u2_Display/add93/c21 ),
    .o({\u2_Display/add93/c22 ,\u2_Display/n2980 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u22  (
    .a(\u2_Display/n2955 ),
    .b(1'b0),
    .c(\u2_Display/add93/c22 ),
    .o({\u2_Display/add93/c23 ,\u2_Display/n2980 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u23  (
    .a(\u2_Display/n2954 ),
    .b(1'b1),
    .c(\u2_Display/add93/c23 ),
    .o({\u2_Display/add93/c24 ,\u2_Display/n2980 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u24  (
    .a(\u2_Display/n2953 ),
    .b(1'b1),
    .c(\u2_Display/add93/c24 ),
    .o({\u2_Display/add93/c25 ,\u2_Display/n2980 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u25  (
    .a(\u2_Display/n2952 ),
    .b(1'b1),
    .c(\u2_Display/add93/c25 ),
    .o({\u2_Display/add93/c26 ,\u2_Display/n2980 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u26  (
    .a(\u2_Display/n2951 ),
    .b(1'b1),
    .c(\u2_Display/add93/c26 ),
    .o({\u2_Display/add93/c27 ,\u2_Display/n2980 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u27  (
    .a(\u2_Display/n2950 ),
    .b(1'b1),
    .c(\u2_Display/add93/c27 ),
    .o({\u2_Display/add93/c28 ,\u2_Display/n2980 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u28  (
    .a(\u2_Display/n2949 ),
    .b(1'b1),
    .c(\u2_Display/add93/c28 ),
    .o({\u2_Display/add93/c29 ,\u2_Display/n2980 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u29  (
    .a(\u2_Display/n2948 ),
    .b(1'b1),
    .c(\u2_Display/add93/c29 ),
    .o({\u2_Display/add93/c30 ,\u2_Display/n2980 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u3  (
    .a(\u2_Display/n2974 ),
    .b(1'b1),
    .c(\u2_Display/add93/c3 ),
    .o({\u2_Display/add93/c4 ,\u2_Display/n2980 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u30  (
    .a(\u2_Display/n2947 ),
    .b(1'b1),
    .c(\u2_Display/add93/c30 ),
    .o({\u2_Display/add93/c31 ,\u2_Display/n2980 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u31  (
    .a(\u2_Display/n2946 ),
    .b(1'b1),
    .c(\u2_Display/add93/c31 ),
    .o({open_n1329,\u2_Display/n2980 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u4  (
    .a(\u2_Display/n2973 ),
    .b(1'b1),
    .c(\u2_Display/add93/c4 ),
    .o({\u2_Display/add93/c5 ,\u2_Display/n2980 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u5  (
    .a(\u2_Display/n2972 ),
    .b(1'b1),
    .c(\u2_Display/add93/c5 ),
    .o({\u2_Display/add93/c6 ,\u2_Display/n2980 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u6  (
    .a(\u2_Display/n2971 ),
    .b(1'b1),
    .c(\u2_Display/add93/c6 ),
    .o({\u2_Display/add93/c7 ,\u2_Display/n2980 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u7  (
    .a(\u2_Display/n2970 ),
    .b(1'b1),
    .c(\u2_Display/add93/c7 ),
    .o({\u2_Display/add93/c8 ,\u2_Display/n2980 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u8  (
    .a(\u2_Display/n2969 ),
    .b(1'b1),
    .c(\u2_Display/add93/c8 ),
    .o({\u2_Display/add93/c9 ,\u2_Display/n2980 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add93/u9  (
    .a(\u2_Display/n2968 ),
    .b(1'b1),
    .c(\u2_Display/add93/c9 ),
    .o({\u2_Display/add93/c10 ,\u2_Display/n2980 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add93/ucin  (
    .a(1'b1),
    .o({\u2_Display/add93/c0 ,open_n1332}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u0  (
    .a(\u2_Display/n3012 ),
    .b(1'b1),
    .c(\u2_Display/add94/c0 ),
    .o({\u2_Display/add94/c1 ,\u2_Display/n3015 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u1  (
    .a(\u2_Display/n3011 ),
    .b(1'b1),
    .c(\u2_Display/add94/c1 ),
    .o({\u2_Display/add94/c2 ,\u2_Display/n3015 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u10  (
    .a(\u2_Display/n3002 ),
    .b(1'b1),
    .c(\u2_Display/add94/c10 ),
    .o({\u2_Display/add94/c11 ,\u2_Display/n3015 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u11  (
    .a(\u2_Display/n3001 ),
    .b(1'b1),
    .c(\u2_Display/add94/c11 ),
    .o({\u2_Display/add94/c12 ,\u2_Display/n3015 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u12  (
    .a(\u2_Display/n3000 ),
    .b(1'b1),
    .c(\u2_Display/add94/c12 ),
    .o({\u2_Display/add94/c13 ,\u2_Display/n3015 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u13  (
    .a(\u2_Display/n2999 ),
    .b(1'b1),
    .c(\u2_Display/add94/c13 ),
    .o({\u2_Display/add94/c14 ,\u2_Display/n3015 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u14  (
    .a(\u2_Display/n2998 ),
    .b(1'b1),
    .c(\u2_Display/add94/c14 ),
    .o({\u2_Display/add94/c15 ,\u2_Display/n3015 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u15  (
    .a(\u2_Display/n2997 ),
    .b(1'b0),
    .c(\u2_Display/add94/c15 ),
    .o({\u2_Display/add94/c16 ,\u2_Display/n3015 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u16  (
    .a(\u2_Display/n2996 ),
    .b(1'b0),
    .c(\u2_Display/add94/c16 ),
    .o({\u2_Display/add94/c17 ,\u2_Display/n3015 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u17  (
    .a(\u2_Display/n2995 ),
    .b(1'b1),
    .c(\u2_Display/add94/c17 ),
    .o({\u2_Display/add94/c18 ,\u2_Display/n3015 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u18  (
    .a(\u2_Display/n2994 ),
    .b(1'b0),
    .c(\u2_Display/add94/c18 ),
    .o({\u2_Display/add94/c19 ,\u2_Display/n3015 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u19  (
    .a(\u2_Display/n2993 ),
    .b(1'b1),
    .c(\u2_Display/add94/c19 ),
    .o({\u2_Display/add94/c20 ,\u2_Display/n3015 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u2  (
    .a(\u2_Display/n3010 ),
    .b(1'b1),
    .c(\u2_Display/add94/c2 ),
    .o({\u2_Display/add94/c3 ,\u2_Display/n3015 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u20  (
    .a(\u2_Display/n2992 ),
    .b(1'b1),
    .c(\u2_Display/add94/c20 ),
    .o({\u2_Display/add94/c21 ,\u2_Display/n3015 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u21  (
    .a(\u2_Display/n2991 ),
    .b(1'b0),
    .c(\u2_Display/add94/c21 ),
    .o({\u2_Display/add94/c22 ,\u2_Display/n3015 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u22  (
    .a(\u2_Display/n2990 ),
    .b(1'b1),
    .c(\u2_Display/add94/c22 ),
    .o({\u2_Display/add94/c23 ,\u2_Display/n3015 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u23  (
    .a(\u2_Display/n2989 ),
    .b(1'b1),
    .c(\u2_Display/add94/c23 ),
    .o({\u2_Display/add94/c24 ,\u2_Display/n3015 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u24  (
    .a(\u2_Display/n2988 ),
    .b(1'b1),
    .c(\u2_Display/add94/c24 ),
    .o({\u2_Display/add94/c25 ,\u2_Display/n3015 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u25  (
    .a(\u2_Display/n2987 ),
    .b(1'b1),
    .c(\u2_Display/add94/c25 ),
    .o({\u2_Display/add94/c26 ,\u2_Display/n3015 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u26  (
    .a(\u2_Display/n2986 ),
    .b(1'b1),
    .c(\u2_Display/add94/c26 ),
    .o({\u2_Display/add94/c27 ,\u2_Display/n3015 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u27  (
    .a(\u2_Display/n2985 ),
    .b(1'b1),
    .c(\u2_Display/add94/c27 ),
    .o({\u2_Display/add94/c28 ,\u2_Display/n3015 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u28  (
    .a(\u2_Display/n2984 ),
    .b(1'b1),
    .c(\u2_Display/add94/c28 ),
    .o({\u2_Display/add94/c29 ,\u2_Display/n3015 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u29  (
    .a(\u2_Display/n2983 ),
    .b(1'b1),
    .c(\u2_Display/add94/c29 ),
    .o({\u2_Display/add94/c30 ,\u2_Display/n3015 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u3  (
    .a(\u2_Display/n3009 ),
    .b(1'b1),
    .c(\u2_Display/add94/c3 ),
    .o({\u2_Display/add94/c4 ,\u2_Display/n3015 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u30  (
    .a(\u2_Display/n2982 ),
    .b(1'b1),
    .c(\u2_Display/add94/c30 ),
    .o({\u2_Display/add94/c31 ,\u2_Display/n3015 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u31  (
    .a(\u2_Display/n2981 ),
    .b(1'b1),
    .c(\u2_Display/add94/c31 ),
    .o({open_n1333,\u2_Display/n3015 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u4  (
    .a(\u2_Display/n3008 ),
    .b(1'b1),
    .c(\u2_Display/add94/c4 ),
    .o({\u2_Display/add94/c5 ,\u2_Display/n3015 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u5  (
    .a(\u2_Display/n3007 ),
    .b(1'b1),
    .c(\u2_Display/add94/c5 ),
    .o({\u2_Display/add94/c6 ,\u2_Display/n3015 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u6  (
    .a(\u2_Display/n3006 ),
    .b(1'b1),
    .c(\u2_Display/add94/c6 ),
    .o({\u2_Display/add94/c7 ,\u2_Display/n3015 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u7  (
    .a(\u2_Display/n3005 ),
    .b(1'b1),
    .c(\u2_Display/add94/c7 ),
    .o({\u2_Display/add94/c8 ,\u2_Display/n3015 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u8  (
    .a(\u2_Display/n3004 ),
    .b(1'b1),
    .c(\u2_Display/add94/c8 ),
    .o({\u2_Display/add94/c9 ,\u2_Display/n3015 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add94/u9  (
    .a(\u2_Display/n3003 ),
    .b(1'b1),
    .c(\u2_Display/add94/c9 ),
    .o({\u2_Display/add94/c10 ,\u2_Display/n3015 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add94/ucin  (
    .a(1'b1),
    .o({\u2_Display/add94/c0 ,open_n1336}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u0  (
    .a(\u2_Display/n3047 ),
    .b(1'b1),
    .c(\u2_Display/add95/c0 ),
    .o({\u2_Display/add95/c1 ,\u2_Display/n3050 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u1  (
    .a(\u2_Display/n3046 ),
    .b(1'b1),
    .c(\u2_Display/add95/c1 ),
    .o({\u2_Display/add95/c2 ,\u2_Display/n3050 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u10  (
    .a(\u2_Display/n3037 ),
    .b(1'b1),
    .c(\u2_Display/add95/c10 ),
    .o({\u2_Display/add95/c11 ,\u2_Display/n3050 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u11  (
    .a(\u2_Display/n3036 ),
    .b(1'b1),
    .c(\u2_Display/add95/c11 ),
    .o({\u2_Display/add95/c12 ,\u2_Display/n3050 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u12  (
    .a(\u2_Display/n3035 ),
    .b(1'b1),
    .c(\u2_Display/add95/c12 ),
    .o({\u2_Display/add95/c13 ,\u2_Display/n3050 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u13  (
    .a(\u2_Display/n3034 ),
    .b(1'b1),
    .c(\u2_Display/add95/c13 ),
    .o({\u2_Display/add95/c14 ,\u2_Display/n3050 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u14  (
    .a(\u2_Display/n3033 ),
    .b(1'b0),
    .c(\u2_Display/add95/c14 ),
    .o({\u2_Display/add95/c15 ,\u2_Display/n3050 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u15  (
    .a(\u2_Display/n3032 ),
    .b(1'b0),
    .c(\u2_Display/add95/c15 ),
    .o({\u2_Display/add95/c16 ,\u2_Display/n3050 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u16  (
    .a(\u2_Display/n3031 ),
    .b(1'b1),
    .c(\u2_Display/add95/c16 ),
    .o({\u2_Display/add95/c17 ,\u2_Display/n3050 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u17  (
    .a(\u2_Display/n3030 ),
    .b(1'b0),
    .c(\u2_Display/add95/c17 ),
    .o({\u2_Display/add95/c18 ,\u2_Display/n3050 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u18  (
    .a(\u2_Display/n3029 ),
    .b(1'b1),
    .c(\u2_Display/add95/c18 ),
    .o({\u2_Display/add95/c19 ,\u2_Display/n3050 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u19  (
    .a(\u2_Display/n3028 ),
    .b(1'b1),
    .c(\u2_Display/add95/c19 ),
    .o({\u2_Display/add95/c20 ,\u2_Display/n3050 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u2  (
    .a(\u2_Display/n3045 ),
    .b(1'b1),
    .c(\u2_Display/add95/c2 ),
    .o({\u2_Display/add95/c3 ,\u2_Display/n3050 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u20  (
    .a(\u2_Display/n3027 ),
    .b(1'b0),
    .c(\u2_Display/add95/c20 ),
    .o({\u2_Display/add95/c21 ,\u2_Display/n3050 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u21  (
    .a(\u2_Display/n3026 ),
    .b(1'b1),
    .c(\u2_Display/add95/c21 ),
    .o({\u2_Display/add95/c22 ,\u2_Display/n3050 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u22  (
    .a(\u2_Display/n3025 ),
    .b(1'b1),
    .c(\u2_Display/add95/c22 ),
    .o({\u2_Display/add95/c23 ,\u2_Display/n3050 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u23  (
    .a(\u2_Display/n3024 ),
    .b(1'b1),
    .c(\u2_Display/add95/c23 ),
    .o({\u2_Display/add95/c24 ,\u2_Display/n3050 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u24  (
    .a(\u2_Display/n3023 ),
    .b(1'b1),
    .c(\u2_Display/add95/c24 ),
    .o({\u2_Display/add95/c25 ,\u2_Display/n3050 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u25  (
    .a(\u2_Display/n3022 ),
    .b(1'b1),
    .c(\u2_Display/add95/c25 ),
    .o({\u2_Display/add95/c26 ,\u2_Display/n3050 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u26  (
    .a(\u2_Display/n3021 ),
    .b(1'b1),
    .c(\u2_Display/add95/c26 ),
    .o({\u2_Display/add95/c27 ,\u2_Display/n3050 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u27  (
    .a(\u2_Display/n3020 ),
    .b(1'b1),
    .c(\u2_Display/add95/c27 ),
    .o({\u2_Display/add95/c28 ,\u2_Display/n3050 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u28  (
    .a(\u2_Display/n3019 ),
    .b(1'b1),
    .c(\u2_Display/add95/c28 ),
    .o({\u2_Display/add95/c29 ,\u2_Display/n3050 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u29  (
    .a(\u2_Display/n3018 ),
    .b(1'b1),
    .c(\u2_Display/add95/c29 ),
    .o({\u2_Display/add95/c30 ,\u2_Display/n3050 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u3  (
    .a(\u2_Display/n3044 ),
    .b(1'b1),
    .c(\u2_Display/add95/c3 ),
    .o({\u2_Display/add95/c4 ,\u2_Display/n3050 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u30  (
    .a(\u2_Display/n3017 ),
    .b(1'b1),
    .c(\u2_Display/add95/c30 ),
    .o({\u2_Display/add95/c31 ,\u2_Display/n3050 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u31  (
    .a(\u2_Display/n3016 ),
    .b(1'b1),
    .c(\u2_Display/add95/c31 ),
    .o({open_n1337,\u2_Display/n3050 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u4  (
    .a(\u2_Display/n3043 ),
    .b(1'b1),
    .c(\u2_Display/add95/c4 ),
    .o({\u2_Display/add95/c5 ,\u2_Display/n3050 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u5  (
    .a(\u2_Display/n3042 ),
    .b(1'b1),
    .c(\u2_Display/add95/c5 ),
    .o({\u2_Display/add95/c6 ,\u2_Display/n3050 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u6  (
    .a(\u2_Display/n3041 ),
    .b(1'b1),
    .c(\u2_Display/add95/c6 ),
    .o({\u2_Display/add95/c7 ,\u2_Display/n3050 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u7  (
    .a(\u2_Display/n3040 ),
    .b(1'b1),
    .c(\u2_Display/add95/c7 ),
    .o({\u2_Display/add95/c8 ,\u2_Display/n3050 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u8  (
    .a(\u2_Display/n3039 ),
    .b(1'b1),
    .c(\u2_Display/add95/c8 ),
    .o({\u2_Display/add95/c9 ,\u2_Display/n3050 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add95/u9  (
    .a(\u2_Display/n3038 ),
    .b(1'b1),
    .c(\u2_Display/add95/c9 ),
    .o({\u2_Display/add95/c10 ,\u2_Display/n3050 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add95/ucin  (
    .a(1'b1),
    .o({\u2_Display/add95/c0 ,open_n1340}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u0  (
    .a(\u2_Display/n3082 ),
    .b(1'b1),
    .c(\u2_Display/add96/c0 ),
    .o({\u2_Display/add96/c1 ,\u2_Display/n3085 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u1  (
    .a(\u2_Display/n3081 ),
    .b(1'b1),
    .c(\u2_Display/add96/c1 ),
    .o({\u2_Display/add96/c2 ,\u2_Display/n3085 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u10  (
    .a(\u2_Display/n3072 ),
    .b(1'b1),
    .c(\u2_Display/add96/c10 ),
    .o({\u2_Display/add96/c11 ,\u2_Display/n3085 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u11  (
    .a(\u2_Display/n3071 ),
    .b(1'b1),
    .c(\u2_Display/add96/c11 ),
    .o({\u2_Display/add96/c12 ,\u2_Display/n3085 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u12  (
    .a(\u2_Display/n3070 ),
    .b(1'b1),
    .c(\u2_Display/add96/c12 ),
    .o({\u2_Display/add96/c13 ,\u2_Display/n3085 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u13  (
    .a(\u2_Display/n3069 ),
    .b(1'b0),
    .c(\u2_Display/add96/c13 ),
    .o({\u2_Display/add96/c14 ,\u2_Display/n3085 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u14  (
    .a(\u2_Display/n3068 ),
    .b(1'b0),
    .c(\u2_Display/add96/c14 ),
    .o({\u2_Display/add96/c15 ,\u2_Display/n3085 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u15  (
    .a(\u2_Display/n3067 ),
    .b(1'b1),
    .c(\u2_Display/add96/c15 ),
    .o({\u2_Display/add96/c16 ,\u2_Display/n3085 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u16  (
    .a(\u2_Display/n3066 ),
    .b(1'b0),
    .c(\u2_Display/add96/c16 ),
    .o({\u2_Display/add96/c17 ,\u2_Display/n3085 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u17  (
    .a(\u2_Display/n3065 ),
    .b(1'b1),
    .c(\u2_Display/add96/c17 ),
    .o({\u2_Display/add96/c18 ,\u2_Display/n3085 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u18  (
    .a(\u2_Display/n3064 ),
    .b(1'b1),
    .c(\u2_Display/add96/c18 ),
    .o({\u2_Display/add96/c19 ,\u2_Display/n3085 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u19  (
    .a(\u2_Display/n3063 ),
    .b(1'b0),
    .c(\u2_Display/add96/c19 ),
    .o({\u2_Display/add96/c20 ,\u2_Display/n3085 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u2  (
    .a(\u2_Display/n3080 ),
    .b(1'b1),
    .c(\u2_Display/add96/c2 ),
    .o({\u2_Display/add96/c3 ,\u2_Display/n3085 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u20  (
    .a(\u2_Display/n3062 ),
    .b(1'b1),
    .c(\u2_Display/add96/c20 ),
    .o({\u2_Display/add96/c21 ,\u2_Display/n3085 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u21  (
    .a(\u2_Display/n3061 ),
    .b(1'b1),
    .c(\u2_Display/add96/c21 ),
    .o({\u2_Display/add96/c22 ,\u2_Display/n3085 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u22  (
    .a(\u2_Display/n3060 ),
    .b(1'b1),
    .c(\u2_Display/add96/c22 ),
    .o({\u2_Display/add96/c23 ,\u2_Display/n3085 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u23  (
    .a(\u2_Display/n3059 ),
    .b(1'b1),
    .c(\u2_Display/add96/c23 ),
    .o({\u2_Display/add96/c24 ,\u2_Display/n3085 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u24  (
    .a(\u2_Display/n3058 ),
    .b(1'b1),
    .c(\u2_Display/add96/c24 ),
    .o({\u2_Display/add96/c25 ,\u2_Display/n3085 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u25  (
    .a(\u2_Display/n3057 ),
    .b(1'b1),
    .c(\u2_Display/add96/c25 ),
    .o({\u2_Display/add96/c26 ,\u2_Display/n3085 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u26  (
    .a(\u2_Display/n3056 ),
    .b(1'b1),
    .c(\u2_Display/add96/c26 ),
    .o({\u2_Display/add96/c27 ,\u2_Display/n3085 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u27  (
    .a(\u2_Display/n3055 ),
    .b(1'b1),
    .c(\u2_Display/add96/c27 ),
    .o({\u2_Display/add96/c28 ,\u2_Display/n3085 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u28  (
    .a(\u2_Display/n3054 ),
    .b(1'b1),
    .c(\u2_Display/add96/c28 ),
    .o({\u2_Display/add96/c29 ,\u2_Display/n3085 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u29  (
    .a(\u2_Display/n3053 ),
    .b(1'b1),
    .c(\u2_Display/add96/c29 ),
    .o({\u2_Display/add96/c30 ,\u2_Display/n3085 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u3  (
    .a(\u2_Display/n3079 ),
    .b(1'b1),
    .c(\u2_Display/add96/c3 ),
    .o({\u2_Display/add96/c4 ,\u2_Display/n3085 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u30  (
    .a(\u2_Display/n3052 ),
    .b(1'b1),
    .c(\u2_Display/add96/c30 ),
    .o({\u2_Display/add96/c31 ,\u2_Display/n3085 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u31  (
    .a(\u2_Display/n3051 ),
    .b(1'b1),
    .c(\u2_Display/add96/c31 ),
    .o({open_n1341,\u2_Display/n3085 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u4  (
    .a(\u2_Display/n3078 ),
    .b(1'b1),
    .c(\u2_Display/add96/c4 ),
    .o({\u2_Display/add96/c5 ,\u2_Display/n3085 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u5  (
    .a(\u2_Display/n3077 ),
    .b(1'b1),
    .c(\u2_Display/add96/c5 ),
    .o({\u2_Display/add96/c6 ,\u2_Display/n3085 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u6  (
    .a(\u2_Display/n3076 ),
    .b(1'b1),
    .c(\u2_Display/add96/c6 ),
    .o({\u2_Display/add96/c7 ,\u2_Display/n3085 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u7  (
    .a(\u2_Display/n3075 ),
    .b(1'b1),
    .c(\u2_Display/add96/c7 ),
    .o({\u2_Display/add96/c8 ,\u2_Display/n3085 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u8  (
    .a(\u2_Display/n3074 ),
    .b(1'b1),
    .c(\u2_Display/add96/c8 ),
    .o({\u2_Display/add96/c9 ,\u2_Display/n3085 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add96/u9  (
    .a(\u2_Display/n3073 ),
    .b(1'b1),
    .c(\u2_Display/add96/c9 ),
    .o({\u2_Display/add96/c10 ,\u2_Display/n3085 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add96/ucin  (
    .a(1'b1),
    .o({\u2_Display/add96/c0 ,open_n1344}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u0  (
    .a(\u2_Display/n3117 ),
    .b(1'b1),
    .c(\u2_Display/add97/c0 ),
    .o({\u2_Display/add97/c1 ,\u2_Display/n3120 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u1  (
    .a(\u2_Display/n3116 ),
    .b(1'b1),
    .c(\u2_Display/add97/c1 ),
    .o({\u2_Display/add97/c2 ,\u2_Display/n3120 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u10  (
    .a(\u2_Display/n3107 ),
    .b(1'b1),
    .c(\u2_Display/add97/c10 ),
    .o({\u2_Display/add97/c11 ,\u2_Display/n3120 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u11  (
    .a(\u2_Display/n3106 ),
    .b(1'b1),
    .c(\u2_Display/add97/c11 ),
    .o({\u2_Display/add97/c12 ,\u2_Display/n3120 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u12  (
    .a(\u2_Display/n3105 ),
    .b(1'b0),
    .c(\u2_Display/add97/c12 ),
    .o({\u2_Display/add97/c13 ,\u2_Display/n3120 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u13  (
    .a(\u2_Display/n3104 ),
    .b(1'b0),
    .c(\u2_Display/add97/c13 ),
    .o({\u2_Display/add97/c14 ,\u2_Display/n3120 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u14  (
    .a(\u2_Display/n3103 ),
    .b(1'b1),
    .c(\u2_Display/add97/c14 ),
    .o({\u2_Display/add97/c15 ,\u2_Display/n3120 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u15  (
    .a(\u2_Display/n3102 ),
    .b(1'b0),
    .c(\u2_Display/add97/c15 ),
    .o({\u2_Display/add97/c16 ,\u2_Display/n3120 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u16  (
    .a(\u2_Display/n3101 ),
    .b(1'b1),
    .c(\u2_Display/add97/c16 ),
    .o({\u2_Display/add97/c17 ,\u2_Display/n3120 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u17  (
    .a(\u2_Display/n3100 ),
    .b(1'b1),
    .c(\u2_Display/add97/c17 ),
    .o({\u2_Display/add97/c18 ,\u2_Display/n3120 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u18  (
    .a(\u2_Display/n3099 ),
    .b(1'b0),
    .c(\u2_Display/add97/c18 ),
    .o({\u2_Display/add97/c19 ,\u2_Display/n3120 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u19  (
    .a(\u2_Display/n3098 ),
    .b(1'b1),
    .c(\u2_Display/add97/c19 ),
    .o({\u2_Display/add97/c20 ,\u2_Display/n3120 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u2  (
    .a(\u2_Display/n3115 ),
    .b(1'b1),
    .c(\u2_Display/add97/c2 ),
    .o({\u2_Display/add97/c3 ,\u2_Display/n3120 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u20  (
    .a(\u2_Display/n3097 ),
    .b(1'b1),
    .c(\u2_Display/add97/c20 ),
    .o({\u2_Display/add97/c21 ,\u2_Display/n3120 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u21  (
    .a(\u2_Display/n3096 ),
    .b(1'b1),
    .c(\u2_Display/add97/c21 ),
    .o({\u2_Display/add97/c22 ,\u2_Display/n3120 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u22  (
    .a(\u2_Display/n3095 ),
    .b(1'b1),
    .c(\u2_Display/add97/c22 ),
    .o({\u2_Display/add97/c23 ,\u2_Display/n3120 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u23  (
    .a(\u2_Display/n3094 ),
    .b(1'b1),
    .c(\u2_Display/add97/c23 ),
    .o({\u2_Display/add97/c24 ,\u2_Display/n3120 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u24  (
    .a(\u2_Display/n3093 ),
    .b(1'b1),
    .c(\u2_Display/add97/c24 ),
    .o({\u2_Display/add97/c25 ,\u2_Display/n3120 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u25  (
    .a(\u2_Display/n3092 ),
    .b(1'b1),
    .c(\u2_Display/add97/c25 ),
    .o({\u2_Display/add97/c26 ,\u2_Display/n3120 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u26  (
    .a(\u2_Display/n3091 ),
    .b(1'b1),
    .c(\u2_Display/add97/c26 ),
    .o({\u2_Display/add97/c27 ,\u2_Display/n3120 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u27  (
    .a(\u2_Display/n3090 ),
    .b(1'b1),
    .c(\u2_Display/add97/c27 ),
    .o({\u2_Display/add97/c28 ,\u2_Display/n3120 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u28  (
    .a(\u2_Display/n3089 ),
    .b(1'b1),
    .c(\u2_Display/add97/c28 ),
    .o({\u2_Display/add97/c29 ,\u2_Display/n3120 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u29  (
    .a(\u2_Display/n3088 ),
    .b(1'b1),
    .c(\u2_Display/add97/c29 ),
    .o({\u2_Display/add97/c30 ,\u2_Display/n3120 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u3  (
    .a(\u2_Display/n3114 ),
    .b(1'b1),
    .c(\u2_Display/add97/c3 ),
    .o({\u2_Display/add97/c4 ,\u2_Display/n3120 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u30  (
    .a(\u2_Display/n3087 ),
    .b(1'b1),
    .c(\u2_Display/add97/c30 ),
    .o({\u2_Display/add97/c31 ,\u2_Display/n3120 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u31  (
    .a(\u2_Display/n3086 ),
    .b(1'b1),
    .c(\u2_Display/add97/c31 ),
    .o({open_n1345,\u2_Display/n3120 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u4  (
    .a(\u2_Display/n3113 ),
    .b(1'b1),
    .c(\u2_Display/add97/c4 ),
    .o({\u2_Display/add97/c5 ,\u2_Display/n3120 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u5  (
    .a(\u2_Display/n3112 ),
    .b(1'b1),
    .c(\u2_Display/add97/c5 ),
    .o({\u2_Display/add97/c6 ,\u2_Display/n3120 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u6  (
    .a(\u2_Display/n3111 ),
    .b(1'b1),
    .c(\u2_Display/add97/c6 ),
    .o({\u2_Display/add97/c7 ,\u2_Display/n3120 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u7  (
    .a(\u2_Display/n3110 ),
    .b(1'b1),
    .c(\u2_Display/add97/c7 ),
    .o({\u2_Display/add97/c8 ,\u2_Display/n3120 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u8  (
    .a(\u2_Display/n3109 ),
    .b(1'b1),
    .c(\u2_Display/add97/c8 ),
    .o({\u2_Display/add97/c9 ,\u2_Display/n3120 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add97/u9  (
    .a(\u2_Display/n3108 ),
    .b(1'b1),
    .c(\u2_Display/add97/c9 ),
    .o({\u2_Display/add97/c10 ,\u2_Display/n3120 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add97/ucin  (
    .a(1'b1),
    .o({\u2_Display/add97/c0 ,open_n1348}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u0  (
    .a(\u2_Display/n3152 ),
    .b(1'b1),
    .c(\u2_Display/add98/c0 ),
    .o({\u2_Display/add98/c1 ,\u2_Display/n3155 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u1  (
    .a(\u2_Display/n3151 ),
    .b(1'b1),
    .c(\u2_Display/add98/c1 ),
    .o({\u2_Display/add98/c2 ,\u2_Display/n3155 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u10  (
    .a(\u2_Display/n3142 ),
    .b(1'b1),
    .c(\u2_Display/add98/c10 ),
    .o({\u2_Display/add98/c11 ,\u2_Display/n3155 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u11  (
    .a(\u2_Display/n3141 ),
    .b(1'b0),
    .c(\u2_Display/add98/c11 ),
    .o({\u2_Display/add98/c12 ,\u2_Display/n3155 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u12  (
    .a(\u2_Display/n3140 ),
    .b(1'b0),
    .c(\u2_Display/add98/c12 ),
    .o({\u2_Display/add98/c13 ,\u2_Display/n3155 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u13  (
    .a(\u2_Display/n3139 ),
    .b(1'b1),
    .c(\u2_Display/add98/c13 ),
    .o({\u2_Display/add98/c14 ,\u2_Display/n3155 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u14  (
    .a(\u2_Display/n3138 ),
    .b(1'b0),
    .c(\u2_Display/add98/c14 ),
    .o({\u2_Display/add98/c15 ,\u2_Display/n3155 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u15  (
    .a(\u2_Display/n3137 ),
    .b(1'b1),
    .c(\u2_Display/add98/c15 ),
    .o({\u2_Display/add98/c16 ,\u2_Display/n3155 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u16  (
    .a(\u2_Display/n3136 ),
    .b(1'b1),
    .c(\u2_Display/add98/c16 ),
    .o({\u2_Display/add98/c17 ,\u2_Display/n3155 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u17  (
    .a(\u2_Display/n3135 ),
    .b(1'b0),
    .c(\u2_Display/add98/c17 ),
    .o({\u2_Display/add98/c18 ,\u2_Display/n3155 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u18  (
    .a(\u2_Display/n3134 ),
    .b(1'b1),
    .c(\u2_Display/add98/c18 ),
    .o({\u2_Display/add98/c19 ,\u2_Display/n3155 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u19  (
    .a(\u2_Display/n3133 ),
    .b(1'b1),
    .c(\u2_Display/add98/c19 ),
    .o({\u2_Display/add98/c20 ,\u2_Display/n3155 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u2  (
    .a(\u2_Display/n3150 ),
    .b(1'b1),
    .c(\u2_Display/add98/c2 ),
    .o({\u2_Display/add98/c3 ,\u2_Display/n3155 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u20  (
    .a(\u2_Display/n3132 ),
    .b(1'b1),
    .c(\u2_Display/add98/c20 ),
    .o({\u2_Display/add98/c21 ,\u2_Display/n3155 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u21  (
    .a(\u2_Display/n3131 ),
    .b(1'b1),
    .c(\u2_Display/add98/c21 ),
    .o({\u2_Display/add98/c22 ,\u2_Display/n3155 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u22  (
    .a(\u2_Display/n3130 ),
    .b(1'b1),
    .c(\u2_Display/add98/c22 ),
    .o({\u2_Display/add98/c23 ,\u2_Display/n3155 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u23  (
    .a(\u2_Display/n3129 ),
    .b(1'b1),
    .c(\u2_Display/add98/c23 ),
    .o({\u2_Display/add98/c24 ,\u2_Display/n3155 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u24  (
    .a(\u2_Display/n3128 ),
    .b(1'b1),
    .c(\u2_Display/add98/c24 ),
    .o({\u2_Display/add98/c25 ,\u2_Display/n3155 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u25  (
    .a(\u2_Display/n3127 ),
    .b(1'b1),
    .c(\u2_Display/add98/c25 ),
    .o({\u2_Display/add98/c26 ,\u2_Display/n3155 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u26  (
    .a(\u2_Display/n3126 ),
    .b(1'b1),
    .c(\u2_Display/add98/c26 ),
    .o({\u2_Display/add98/c27 ,\u2_Display/n3155 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u27  (
    .a(\u2_Display/n3125 ),
    .b(1'b1),
    .c(\u2_Display/add98/c27 ),
    .o({\u2_Display/add98/c28 ,\u2_Display/n3155 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u28  (
    .a(\u2_Display/n3124 ),
    .b(1'b1),
    .c(\u2_Display/add98/c28 ),
    .o({\u2_Display/add98/c29 ,\u2_Display/n3155 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u29  (
    .a(\u2_Display/n3123 ),
    .b(1'b1),
    .c(\u2_Display/add98/c29 ),
    .o({\u2_Display/add98/c30 ,\u2_Display/n3155 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u3  (
    .a(\u2_Display/n3149 ),
    .b(1'b1),
    .c(\u2_Display/add98/c3 ),
    .o({\u2_Display/add98/c4 ,\u2_Display/n3155 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u30  (
    .a(\u2_Display/n3122 ),
    .b(1'b1),
    .c(\u2_Display/add98/c30 ),
    .o({\u2_Display/add98/c31 ,\u2_Display/n3155 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u31  (
    .a(\u2_Display/n3121 ),
    .b(1'b1),
    .c(\u2_Display/add98/c31 ),
    .o({open_n1349,\u2_Display/n3155 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u4  (
    .a(\u2_Display/n3148 ),
    .b(1'b1),
    .c(\u2_Display/add98/c4 ),
    .o({\u2_Display/add98/c5 ,\u2_Display/n3155 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u5  (
    .a(\u2_Display/n3147 ),
    .b(1'b1),
    .c(\u2_Display/add98/c5 ),
    .o({\u2_Display/add98/c6 ,\u2_Display/n3155 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u6  (
    .a(\u2_Display/n3146 ),
    .b(1'b1),
    .c(\u2_Display/add98/c6 ),
    .o({\u2_Display/add98/c7 ,\u2_Display/n3155 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u7  (
    .a(\u2_Display/n3145 ),
    .b(1'b1),
    .c(\u2_Display/add98/c7 ),
    .o({\u2_Display/add98/c8 ,\u2_Display/n3155 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u8  (
    .a(\u2_Display/n3144 ),
    .b(1'b1),
    .c(\u2_Display/add98/c8 ),
    .o({\u2_Display/add98/c9 ,\u2_Display/n3155 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add98/u9  (
    .a(\u2_Display/n3143 ),
    .b(1'b1),
    .c(\u2_Display/add98/c9 ),
    .o({\u2_Display/add98/c10 ,\u2_Display/n3155 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add98/ucin  (
    .a(1'b1),
    .o({\u2_Display/add98/c0 ,open_n1352}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u0  (
    .a(\u2_Display/n3187 ),
    .b(1'b1),
    .c(\u2_Display/add99/c0 ),
    .o({\u2_Display/add99/c1 ,\u2_Display/n3190 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u1  (
    .a(\u2_Display/n3186 ),
    .b(1'b1),
    .c(\u2_Display/add99/c1 ),
    .o({\u2_Display/add99/c2 ,\u2_Display/n3190 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u10  (
    .a(\u2_Display/n3177 ),
    .b(1'b0),
    .c(\u2_Display/add99/c10 ),
    .o({\u2_Display/add99/c11 ,\u2_Display/n3190 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u11  (
    .a(\u2_Display/n3176 ),
    .b(1'b0),
    .c(\u2_Display/add99/c11 ),
    .o({\u2_Display/add99/c12 ,\u2_Display/n3190 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u12  (
    .a(\u2_Display/n3175 ),
    .b(1'b1),
    .c(\u2_Display/add99/c12 ),
    .o({\u2_Display/add99/c13 ,\u2_Display/n3190 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u13  (
    .a(\u2_Display/n3174 ),
    .b(1'b0),
    .c(\u2_Display/add99/c13 ),
    .o({\u2_Display/add99/c14 ,\u2_Display/n3190 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u14  (
    .a(\u2_Display/n3173 ),
    .b(1'b1),
    .c(\u2_Display/add99/c14 ),
    .o({\u2_Display/add99/c15 ,\u2_Display/n3190 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u15  (
    .a(\u2_Display/n3172 ),
    .b(1'b1),
    .c(\u2_Display/add99/c15 ),
    .o({\u2_Display/add99/c16 ,\u2_Display/n3190 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u16  (
    .a(\u2_Display/n3171 ),
    .b(1'b0),
    .c(\u2_Display/add99/c16 ),
    .o({\u2_Display/add99/c17 ,\u2_Display/n3190 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u17  (
    .a(\u2_Display/n3170 ),
    .b(1'b1),
    .c(\u2_Display/add99/c17 ),
    .o({\u2_Display/add99/c18 ,\u2_Display/n3190 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u18  (
    .a(\u2_Display/n3169 ),
    .b(1'b1),
    .c(\u2_Display/add99/c18 ),
    .o({\u2_Display/add99/c19 ,\u2_Display/n3190 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u19  (
    .a(\u2_Display/n3168 ),
    .b(1'b1),
    .c(\u2_Display/add99/c19 ),
    .o({\u2_Display/add99/c20 ,\u2_Display/n3190 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u2  (
    .a(\u2_Display/n3185 ),
    .b(1'b1),
    .c(\u2_Display/add99/c2 ),
    .o({\u2_Display/add99/c3 ,\u2_Display/n3190 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u20  (
    .a(\u2_Display/n3167 ),
    .b(1'b1),
    .c(\u2_Display/add99/c20 ),
    .o({\u2_Display/add99/c21 ,\u2_Display/n3190 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u21  (
    .a(\u2_Display/n3166 ),
    .b(1'b1),
    .c(\u2_Display/add99/c21 ),
    .o({\u2_Display/add99/c22 ,\u2_Display/n3190 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u22  (
    .a(\u2_Display/n3165 ),
    .b(1'b1),
    .c(\u2_Display/add99/c22 ),
    .o({\u2_Display/add99/c23 ,\u2_Display/n3190 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u23  (
    .a(\u2_Display/n3164 ),
    .b(1'b1),
    .c(\u2_Display/add99/c23 ),
    .o({\u2_Display/add99/c24 ,\u2_Display/n3190 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u24  (
    .a(\u2_Display/n3163 ),
    .b(1'b1),
    .c(\u2_Display/add99/c24 ),
    .o({\u2_Display/add99/c25 ,\u2_Display/n3190 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u25  (
    .a(\u2_Display/n3162 ),
    .b(1'b1),
    .c(\u2_Display/add99/c25 ),
    .o({\u2_Display/add99/c26 ,\u2_Display/n3190 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u26  (
    .a(\u2_Display/n3161 ),
    .b(1'b1),
    .c(\u2_Display/add99/c26 ),
    .o({\u2_Display/add99/c27 ,\u2_Display/n3190 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u27  (
    .a(\u2_Display/n3160 ),
    .b(1'b1),
    .c(\u2_Display/add99/c27 ),
    .o({\u2_Display/add99/c28 ,\u2_Display/n3190 [27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u28  (
    .a(\u2_Display/n3159 ),
    .b(1'b1),
    .c(\u2_Display/add99/c28 ),
    .o({\u2_Display/add99/c29 ,\u2_Display/n3190 [28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u29  (
    .a(\u2_Display/n3158 ),
    .b(1'b1),
    .c(\u2_Display/add99/c29 ),
    .o({\u2_Display/add99/c30 ,\u2_Display/n3190 [29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u3  (
    .a(\u2_Display/n3184 ),
    .b(1'b1),
    .c(\u2_Display/add99/c3 ),
    .o({\u2_Display/add99/c4 ,\u2_Display/n3190 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u30  (
    .a(\u2_Display/n3157 ),
    .b(1'b1),
    .c(\u2_Display/add99/c30 ),
    .o({\u2_Display/add99/c31 ,\u2_Display/n3190 [30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u31  (
    .a(\u2_Display/n3156 ),
    .b(1'b1),
    .c(\u2_Display/add99/c31 ),
    .o({open_n1353,\u2_Display/n3190 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u4  (
    .a(\u2_Display/n3183 ),
    .b(1'b1),
    .c(\u2_Display/add99/c4 ),
    .o({\u2_Display/add99/c5 ,\u2_Display/n3190 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u5  (
    .a(\u2_Display/n3182 ),
    .b(1'b1),
    .c(\u2_Display/add99/c5 ),
    .o({\u2_Display/add99/c6 ,\u2_Display/n3190 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u6  (
    .a(\u2_Display/n3181 ),
    .b(1'b1),
    .c(\u2_Display/add99/c6 ),
    .o({\u2_Display/add99/c7 ,\u2_Display/n3190 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u7  (
    .a(\u2_Display/n3180 ),
    .b(1'b1),
    .c(\u2_Display/add99/c7 ),
    .o({\u2_Display/add99/c8 ,\u2_Display/n3190 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u8  (
    .a(\u2_Display/n3179 ),
    .b(1'b1),
    .c(\u2_Display/add99/c8 ),
    .o({\u2_Display/add99/c9 ,\u2_Display/n3190 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u2_Display/add99/u9  (
    .a(\u2_Display/n3178 ),
    .b(1'b1),
    .c(\u2_Display/add99/c9 ),
    .o({\u2_Display/add99/c10 ,\u2_Display/n3190 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u2_Display/add99/ucin  (
    .a(1'b1),
    .o({\u2_Display/add99/c0 ,open_n1356}));
  reg_ar_as_w1 \u2_Display/clk1s_reg  (
    .clk(clk_vga),
    .d(\u2_Display/n36 ),
    .en(\u2_Display/n35 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/clk1s ));  // source/rtl/Display.v(61)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt0_2_0  (
    .a(lcd_xpos[0]),
    .b(\u2_Display/i [0]),
    .c(\u2_Display/lt0_2_c0 ),
    .o({\u2_Display/lt0_2_c1 ,open_n1357}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt0_2_1  (
    .a(lcd_xpos[1]),
    .b(\u2_Display/i [1]),
    .c(\u2_Display/lt0_2_c1 ),
    .o({\u2_Display/lt0_2_c2 ,open_n1358}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt0_2_10  (
    .a(lcd_xpos[10]),
    .b(\u2_Display/n43 [2]),
    .c(\u2_Display/lt0_2_c10 ),
    .o({\u2_Display/lt0_2_c11 ,open_n1359}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt0_2_11  (
    .a(lcd_xpos[11]),
    .b(\u2_Display/add2_2_co ),
    .c(\u2_Display/lt0_2_c11 ),
    .o({\u2_Display/lt0_2_c12 ,open_n1360}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt0_2_2  (
    .a(lcd_xpos[2]),
    .b(\u2_Display/i [2]),
    .c(\u2_Display/lt0_2_c2 ),
    .o({\u2_Display/lt0_2_c3 ,open_n1361}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt0_2_3  (
    .a(lcd_xpos[3]),
    .b(\u2_Display/i [3]),
    .c(\u2_Display/lt0_2_c3 ),
    .o({\u2_Display/lt0_2_c4 ,open_n1362}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt0_2_4  (
    .a(lcd_xpos[4]),
    .b(\u2_Display/i [4]),
    .c(\u2_Display/lt0_2_c4 ),
    .o({\u2_Display/lt0_2_c5 ,open_n1363}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt0_2_5  (
    .a(lcd_xpos[5]),
    .b(\u2_Display/i [5]),
    .c(\u2_Display/lt0_2_c5 ),
    .o({\u2_Display/lt0_2_c6 ,open_n1364}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt0_2_6  (
    .a(lcd_xpos[6]),
    .b(\u2_Display/i [6]),
    .c(\u2_Display/lt0_2_c6 ),
    .o({\u2_Display/lt0_2_c7 ,open_n1365}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt0_2_7  (
    .a(lcd_xpos[7]),
    .b(\u2_Display/i [7]),
    .c(\u2_Display/lt0_2_c7 ),
    .o({\u2_Display/lt0_2_c8 ,open_n1366}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt0_2_8  (
    .a(lcd_xpos[8]),
    .b(\u2_Display/n43 [0]),
    .c(\u2_Display/lt0_2_c8 ),
    .o({\u2_Display/lt0_2_c9 ,open_n1367}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt0_2_9  (
    .a(lcd_xpos[9]),
    .b(\u2_Display/n43 [1]),
    .c(\u2_Display/lt0_2_c9 ),
    .o({\u2_Display/lt0_2_c10 ,open_n1368}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt0_2_cin  (
    .a(1'b0),
    .o({\u2_Display/lt0_2_c0 ,open_n1371}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt0_2_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt0_2_c12 ),
    .o({open_n1372,\u2_Display/n44 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_0  (
    .a(\u2_Display/n3082 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c0 ),
    .o({\u2_Display/lt100_c1 ,open_n1373}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_1  (
    .a(\u2_Display/n3081 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c1 ),
    .o({\u2_Display/lt100_c2 ,open_n1374}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_10  (
    .a(\u2_Display/n3072 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c10 ),
    .o({\u2_Display/lt100_c11 ,open_n1375}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_11  (
    .a(\u2_Display/n3071 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c11 ),
    .o({\u2_Display/lt100_c12 ,open_n1376}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_12  (
    .a(\u2_Display/n3070 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c12 ),
    .o({\u2_Display/lt100_c13 ,open_n1377}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_13  (
    .a(\u2_Display/n3069 ),
    .b(1'b1),
    .c(\u2_Display/lt100_c13 ),
    .o({\u2_Display/lt100_c14 ,open_n1378}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_14  (
    .a(\u2_Display/n3068 ),
    .b(1'b1),
    .c(\u2_Display/lt100_c14 ),
    .o({\u2_Display/lt100_c15 ,open_n1379}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_15  (
    .a(\u2_Display/n3067 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c15 ),
    .o({\u2_Display/lt100_c16 ,open_n1380}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_16  (
    .a(\u2_Display/n3066 ),
    .b(1'b1),
    .c(\u2_Display/lt100_c16 ),
    .o({\u2_Display/lt100_c17 ,open_n1381}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_17  (
    .a(\u2_Display/n3065 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c17 ),
    .o({\u2_Display/lt100_c18 ,open_n1382}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_18  (
    .a(\u2_Display/n3064 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c18 ),
    .o({\u2_Display/lt100_c19 ,open_n1383}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_19  (
    .a(\u2_Display/n3063 ),
    .b(1'b1),
    .c(\u2_Display/lt100_c19 ),
    .o({\u2_Display/lt100_c20 ,open_n1384}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_2  (
    .a(\u2_Display/n3080 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c2 ),
    .o({\u2_Display/lt100_c3 ,open_n1385}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_20  (
    .a(\u2_Display/n3062 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c20 ),
    .o({\u2_Display/lt100_c21 ,open_n1386}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_21  (
    .a(\u2_Display/n3061 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c21 ),
    .o({\u2_Display/lt100_c22 ,open_n1387}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_22  (
    .a(\u2_Display/n3060 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c22 ),
    .o({\u2_Display/lt100_c23 ,open_n1388}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_23  (
    .a(\u2_Display/n3059 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c23 ),
    .o({\u2_Display/lt100_c24 ,open_n1389}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_24  (
    .a(\u2_Display/n3058 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c24 ),
    .o({\u2_Display/lt100_c25 ,open_n1390}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_25  (
    .a(\u2_Display/n3057 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c25 ),
    .o({\u2_Display/lt100_c26 ,open_n1391}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_26  (
    .a(\u2_Display/n3056 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c26 ),
    .o({\u2_Display/lt100_c27 ,open_n1392}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_27  (
    .a(\u2_Display/n3055 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c27 ),
    .o({\u2_Display/lt100_c28 ,open_n1393}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_28  (
    .a(\u2_Display/n3054 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c28 ),
    .o({\u2_Display/lt100_c29 ,open_n1394}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_29  (
    .a(\u2_Display/n3053 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c29 ),
    .o({\u2_Display/lt100_c30 ,open_n1395}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_3  (
    .a(\u2_Display/n3079 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c3 ),
    .o({\u2_Display/lt100_c4 ,open_n1396}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_30  (
    .a(\u2_Display/n3052 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c30 ),
    .o({\u2_Display/lt100_c31 ,open_n1397}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_31  (
    .a(\u2_Display/n3051 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c31 ),
    .o({\u2_Display/lt100_c32 ,open_n1398}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_4  (
    .a(\u2_Display/n3078 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c4 ),
    .o({\u2_Display/lt100_c5 ,open_n1399}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_5  (
    .a(\u2_Display/n3077 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c5 ),
    .o({\u2_Display/lt100_c6 ,open_n1400}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_6  (
    .a(\u2_Display/n3076 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c6 ),
    .o({\u2_Display/lt100_c7 ,open_n1401}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_7  (
    .a(\u2_Display/n3075 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c7 ),
    .o({\u2_Display/lt100_c8 ,open_n1402}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_8  (
    .a(\u2_Display/n3074 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c8 ),
    .o({\u2_Display/lt100_c9 ,open_n1403}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_9  (
    .a(\u2_Display/n3073 ),
    .b(1'b0),
    .c(\u2_Display/lt100_c9 ),
    .o({\u2_Display/lt100_c10 ,open_n1404}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt100_cin  (
    .a(1'b0),
    .o({\u2_Display/lt100_c0 ,open_n1407}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt100_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt100_c32 ),
    .o({open_n1408,\u2_Display/n3083 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_0  (
    .a(\u2_Display/n3117 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c0 ),
    .o({\u2_Display/lt101_c1 ,open_n1409}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_1  (
    .a(\u2_Display/n3116 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c1 ),
    .o({\u2_Display/lt101_c2 ,open_n1410}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_10  (
    .a(\u2_Display/n3107 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c10 ),
    .o({\u2_Display/lt101_c11 ,open_n1411}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_11  (
    .a(\u2_Display/n3106 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c11 ),
    .o({\u2_Display/lt101_c12 ,open_n1412}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_12  (
    .a(\u2_Display/n3105 ),
    .b(1'b1),
    .c(\u2_Display/lt101_c12 ),
    .o({\u2_Display/lt101_c13 ,open_n1413}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_13  (
    .a(\u2_Display/n3104 ),
    .b(1'b1),
    .c(\u2_Display/lt101_c13 ),
    .o({\u2_Display/lt101_c14 ,open_n1414}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_14  (
    .a(\u2_Display/n3103 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c14 ),
    .o({\u2_Display/lt101_c15 ,open_n1415}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_15  (
    .a(\u2_Display/n3102 ),
    .b(1'b1),
    .c(\u2_Display/lt101_c15 ),
    .o({\u2_Display/lt101_c16 ,open_n1416}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_16  (
    .a(\u2_Display/n3101 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c16 ),
    .o({\u2_Display/lt101_c17 ,open_n1417}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_17  (
    .a(\u2_Display/n3100 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c17 ),
    .o({\u2_Display/lt101_c18 ,open_n1418}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_18  (
    .a(\u2_Display/n3099 ),
    .b(1'b1),
    .c(\u2_Display/lt101_c18 ),
    .o({\u2_Display/lt101_c19 ,open_n1419}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_19  (
    .a(\u2_Display/n3098 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c19 ),
    .o({\u2_Display/lt101_c20 ,open_n1420}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_2  (
    .a(\u2_Display/n3115 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c2 ),
    .o({\u2_Display/lt101_c3 ,open_n1421}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_20  (
    .a(\u2_Display/n3097 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c20 ),
    .o({\u2_Display/lt101_c21 ,open_n1422}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_21  (
    .a(\u2_Display/n3096 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c21 ),
    .o({\u2_Display/lt101_c22 ,open_n1423}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_22  (
    .a(\u2_Display/n3095 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c22 ),
    .o({\u2_Display/lt101_c23 ,open_n1424}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_23  (
    .a(\u2_Display/n3094 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c23 ),
    .o({\u2_Display/lt101_c24 ,open_n1425}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_24  (
    .a(\u2_Display/n3093 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c24 ),
    .o({\u2_Display/lt101_c25 ,open_n1426}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_25  (
    .a(\u2_Display/n3092 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c25 ),
    .o({\u2_Display/lt101_c26 ,open_n1427}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_26  (
    .a(\u2_Display/n3091 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c26 ),
    .o({\u2_Display/lt101_c27 ,open_n1428}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_27  (
    .a(\u2_Display/n3090 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c27 ),
    .o({\u2_Display/lt101_c28 ,open_n1429}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_28  (
    .a(\u2_Display/n3089 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c28 ),
    .o({\u2_Display/lt101_c29 ,open_n1430}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_29  (
    .a(\u2_Display/n3088 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c29 ),
    .o({\u2_Display/lt101_c30 ,open_n1431}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_3  (
    .a(\u2_Display/n3114 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c3 ),
    .o({\u2_Display/lt101_c4 ,open_n1432}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_30  (
    .a(\u2_Display/n3087 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c30 ),
    .o({\u2_Display/lt101_c31 ,open_n1433}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_31  (
    .a(\u2_Display/n3086 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c31 ),
    .o({\u2_Display/lt101_c32 ,open_n1434}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_4  (
    .a(\u2_Display/n3113 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c4 ),
    .o({\u2_Display/lt101_c5 ,open_n1435}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_5  (
    .a(\u2_Display/n3112 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c5 ),
    .o({\u2_Display/lt101_c6 ,open_n1436}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_6  (
    .a(\u2_Display/n3111 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c6 ),
    .o({\u2_Display/lt101_c7 ,open_n1437}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_7  (
    .a(\u2_Display/n3110 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c7 ),
    .o({\u2_Display/lt101_c8 ,open_n1438}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_8  (
    .a(\u2_Display/n3109 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c8 ),
    .o({\u2_Display/lt101_c9 ,open_n1439}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_9  (
    .a(\u2_Display/n3108 ),
    .b(1'b0),
    .c(\u2_Display/lt101_c9 ),
    .o({\u2_Display/lt101_c10 ,open_n1440}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt101_cin  (
    .a(1'b0),
    .o({\u2_Display/lt101_c0 ,open_n1443}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt101_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt101_c32 ),
    .o({open_n1444,\u2_Display/n3118 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_0  (
    .a(\u2_Display/n3152 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c0 ),
    .o({\u2_Display/lt102_c1 ,open_n1445}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_1  (
    .a(\u2_Display/n3151 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c1 ),
    .o({\u2_Display/lt102_c2 ,open_n1446}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_10  (
    .a(\u2_Display/n3142 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c10 ),
    .o({\u2_Display/lt102_c11 ,open_n1447}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_11  (
    .a(\u2_Display/n3141 ),
    .b(1'b1),
    .c(\u2_Display/lt102_c11 ),
    .o({\u2_Display/lt102_c12 ,open_n1448}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_12  (
    .a(\u2_Display/n3140 ),
    .b(1'b1),
    .c(\u2_Display/lt102_c12 ),
    .o({\u2_Display/lt102_c13 ,open_n1449}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_13  (
    .a(\u2_Display/n3139 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c13 ),
    .o({\u2_Display/lt102_c14 ,open_n1450}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_14  (
    .a(\u2_Display/n3138 ),
    .b(1'b1),
    .c(\u2_Display/lt102_c14 ),
    .o({\u2_Display/lt102_c15 ,open_n1451}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_15  (
    .a(\u2_Display/n3137 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c15 ),
    .o({\u2_Display/lt102_c16 ,open_n1452}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_16  (
    .a(\u2_Display/n3136 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c16 ),
    .o({\u2_Display/lt102_c17 ,open_n1453}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_17  (
    .a(\u2_Display/n3135 ),
    .b(1'b1),
    .c(\u2_Display/lt102_c17 ),
    .o({\u2_Display/lt102_c18 ,open_n1454}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_18  (
    .a(\u2_Display/n3134 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c18 ),
    .o({\u2_Display/lt102_c19 ,open_n1455}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_19  (
    .a(\u2_Display/n3133 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c19 ),
    .o({\u2_Display/lt102_c20 ,open_n1456}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_2  (
    .a(\u2_Display/n3150 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c2 ),
    .o({\u2_Display/lt102_c3 ,open_n1457}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_20  (
    .a(\u2_Display/n3132 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c20 ),
    .o({\u2_Display/lt102_c21 ,open_n1458}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_21  (
    .a(\u2_Display/n3131 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c21 ),
    .o({\u2_Display/lt102_c22 ,open_n1459}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_22  (
    .a(\u2_Display/n3130 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c22 ),
    .o({\u2_Display/lt102_c23 ,open_n1460}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_23  (
    .a(\u2_Display/n3129 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c23 ),
    .o({\u2_Display/lt102_c24 ,open_n1461}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_24  (
    .a(\u2_Display/n3128 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c24 ),
    .o({\u2_Display/lt102_c25 ,open_n1462}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_25  (
    .a(\u2_Display/n3127 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c25 ),
    .o({\u2_Display/lt102_c26 ,open_n1463}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_26  (
    .a(\u2_Display/n3126 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c26 ),
    .o({\u2_Display/lt102_c27 ,open_n1464}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_27  (
    .a(\u2_Display/n3125 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c27 ),
    .o({\u2_Display/lt102_c28 ,open_n1465}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_28  (
    .a(\u2_Display/n3124 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c28 ),
    .o({\u2_Display/lt102_c29 ,open_n1466}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_29  (
    .a(\u2_Display/n3123 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c29 ),
    .o({\u2_Display/lt102_c30 ,open_n1467}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_3  (
    .a(\u2_Display/n3149 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c3 ),
    .o({\u2_Display/lt102_c4 ,open_n1468}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_30  (
    .a(\u2_Display/n3122 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c30 ),
    .o({\u2_Display/lt102_c31 ,open_n1469}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_31  (
    .a(\u2_Display/n3121 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c31 ),
    .o({\u2_Display/lt102_c32 ,open_n1470}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_4  (
    .a(\u2_Display/n3148 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c4 ),
    .o({\u2_Display/lt102_c5 ,open_n1471}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_5  (
    .a(\u2_Display/n3147 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c5 ),
    .o({\u2_Display/lt102_c6 ,open_n1472}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_6  (
    .a(\u2_Display/n3146 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c6 ),
    .o({\u2_Display/lt102_c7 ,open_n1473}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_7  (
    .a(\u2_Display/n3145 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c7 ),
    .o({\u2_Display/lt102_c8 ,open_n1474}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_8  (
    .a(\u2_Display/n3144 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c8 ),
    .o({\u2_Display/lt102_c9 ,open_n1475}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_9  (
    .a(\u2_Display/n3143 ),
    .b(1'b0),
    .c(\u2_Display/lt102_c9 ),
    .o({\u2_Display/lt102_c10 ,open_n1476}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt102_cin  (
    .a(1'b0),
    .o({\u2_Display/lt102_c0 ,open_n1479}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt102_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt102_c32 ),
    .o({open_n1480,\u2_Display/n3153 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_0  (
    .a(\u2_Display/n3187 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c0 ),
    .o({\u2_Display/lt103_c1 ,open_n1481}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_1  (
    .a(\u2_Display/n3186 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c1 ),
    .o({\u2_Display/lt103_c2 ,open_n1482}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_10  (
    .a(\u2_Display/n3177 ),
    .b(1'b1),
    .c(\u2_Display/lt103_c10 ),
    .o({\u2_Display/lt103_c11 ,open_n1483}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_11  (
    .a(\u2_Display/n3176 ),
    .b(1'b1),
    .c(\u2_Display/lt103_c11 ),
    .o({\u2_Display/lt103_c12 ,open_n1484}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_12  (
    .a(\u2_Display/n3175 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c12 ),
    .o({\u2_Display/lt103_c13 ,open_n1485}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_13  (
    .a(\u2_Display/n3174 ),
    .b(1'b1),
    .c(\u2_Display/lt103_c13 ),
    .o({\u2_Display/lt103_c14 ,open_n1486}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_14  (
    .a(\u2_Display/n3173 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c14 ),
    .o({\u2_Display/lt103_c15 ,open_n1487}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_15  (
    .a(\u2_Display/n3172 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c15 ),
    .o({\u2_Display/lt103_c16 ,open_n1488}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_16  (
    .a(\u2_Display/n3171 ),
    .b(1'b1),
    .c(\u2_Display/lt103_c16 ),
    .o({\u2_Display/lt103_c17 ,open_n1489}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_17  (
    .a(\u2_Display/n3170 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c17 ),
    .o({\u2_Display/lt103_c18 ,open_n1490}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_18  (
    .a(\u2_Display/n3169 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c18 ),
    .o({\u2_Display/lt103_c19 ,open_n1491}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_19  (
    .a(\u2_Display/n3168 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c19 ),
    .o({\u2_Display/lt103_c20 ,open_n1492}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_2  (
    .a(\u2_Display/n3185 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c2 ),
    .o({\u2_Display/lt103_c3 ,open_n1493}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_20  (
    .a(\u2_Display/n3167 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c20 ),
    .o({\u2_Display/lt103_c21 ,open_n1494}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_21  (
    .a(\u2_Display/n3166 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c21 ),
    .o({\u2_Display/lt103_c22 ,open_n1495}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_22  (
    .a(\u2_Display/n3165 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c22 ),
    .o({\u2_Display/lt103_c23 ,open_n1496}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_23  (
    .a(\u2_Display/n3164 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c23 ),
    .o({\u2_Display/lt103_c24 ,open_n1497}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_24  (
    .a(\u2_Display/n3163 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c24 ),
    .o({\u2_Display/lt103_c25 ,open_n1498}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_25  (
    .a(\u2_Display/n3162 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c25 ),
    .o({\u2_Display/lt103_c26 ,open_n1499}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_26  (
    .a(\u2_Display/n3161 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c26 ),
    .o({\u2_Display/lt103_c27 ,open_n1500}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_27  (
    .a(\u2_Display/n3160 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c27 ),
    .o({\u2_Display/lt103_c28 ,open_n1501}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_28  (
    .a(\u2_Display/n3159 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c28 ),
    .o({\u2_Display/lt103_c29 ,open_n1502}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_29  (
    .a(\u2_Display/n3158 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c29 ),
    .o({\u2_Display/lt103_c30 ,open_n1503}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_3  (
    .a(\u2_Display/n3184 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c3 ),
    .o({\u2_Display/lt103_c4 ,open_n1504}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_30  (
    .a(\u2_Display/n3157 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c30 ),
    .o({\u2_Display/lt103_c31 ,open_n1505}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_31  (
    .a(\u2_Display/n3156 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c31 ),
    .o({\u2_Display/lt103_c32 ,open_n1506}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_4  (
    .a(\u2_Display/n3183 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c4 ),
    .o({\u2_Display/lt103_c5 ,open_n1507}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_5  (
    .a(\u2_Display/n3182 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c5 ),
    .o({\u2_Display/lt103_c6 ,open_n1508}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_6  (
    .a(\u2_Display/n3181 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c6 ),
    .o({\u2_Display/lt103_c7 ,open_n1509}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_7  (
    .a(\u2_Display/n3180 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c7 ),
    .o({\u2_Display/lt103_c8 ,open_n1510}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_8  (
    .a(\u2_Display/n3179 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c8 ),
    .o({\u2_Display/lt103_c9 ,open_n1511}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_9  (
    .a(\u2_Display/n3178 ),
    .b(1'b0),
    .c(\u2_Display/lt103_c9 ),
    .o({\u2_Display/lt103_c10 ,open_n1512}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt103_cin  (
    .a(1'b0),
    .o({\u2_Display/lt103_c0 ,open_n1515}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt103_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt103_c32 ),
    .o({open_n1516,\u2_Display/n3188 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_0  (
    .a(\u2_Display/n3222 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c0 ),
    .o({\u2_Display/lt104_c1 ,open_n1517}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_1  (
    .a(\u2_Display/n3221 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c1 ),
    .o({\u2_Display/lt104_c2 ,open_n1518}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_10  (
    .a(\u2_Display/n3212 ),
    .b(1'b1),
    .c(\u2_Display/lt104_c10 ),
    .o({\u2_Display/lt104_c11 ,open_n1519}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_11  (
    .a(\u2_Display/n3211 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c11 ),
    .o({\u2_Display/lt104_c12 ,open_n1520}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_12  (
    .a(\u2_Display/n3210 ),
    .b(1'b1),
    .c(\u2_Display/lt104_c12 ),
    .o({\u2_Display/lt104_c13 ,open_n1521}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_13  (
    .a(\u2_Display/n3209 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c13 ),
    .o({\u2_Display/lt104_c14 ,open_n1522}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_14  (
    .a(\u2_Display/n3208 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c14 ),
    .o({\u2_Display/lt104_c15 ,open_n1523}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_15  (
    .a(\u2_Display/n3207 ),
    .b(1'b1),
    .c(\u2_Display/lt104_c15 ),
    .o({\u2_Display/lt104_c16 ,open_n1524}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_16  (
    .a(\u2_Display/n3206 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c16 ),
    .o({\u2_Display/lt104_c17 ,open_n1525}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_17  (
    .a(\u2_Display/n3205 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c17 ),
    .o({\u2_Display/lt104_c18 ,open_n1526}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_18  (
    .a(\u2_Display/n3204 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c18 ),
    .o({\u2_Display/lt104_c19 ,open_n1527}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_19  (
    .a(\u2_Display/n3203 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c19 ),
    .o({\u2_Display/lt104_c20 ,open_n1528}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_2  (
    .a(\u2_Display/n3220 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c2 ),
    .o({\u2_Display/lt104_c3 ,open_n1529}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_20  (
    .a(\u2_Display/n3202 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c20 ),
    .o({\u2_Display/lt104_c21 ,open_n1530}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_21  (
    .a(\u2_Display/n3201 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c21 ),
    .o({\u2_Display/lt104_c22 ,open_n1531}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_22  (
    .a(\u2_Display/n3200 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c22 ),
    .o({\u2_Display/lt104_c23 ,open_n1532}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_23  (
    .a(\u2_Display/n3199 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c23 ),
    .o({\u2_Display/lt104_c24 ,open_n1533}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_24  (
    .a(\u2_Display/n3198 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c24 ),
    .o({\u2_Display/lt104_c25 ,open_n1534}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_25  (
    .a(\u2_Display/n3197 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c25 ),
    .o({\u2_Display/lt104_c26 ,open_n1535}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_26  (
    .a(\u2_Display/n3196 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c26 ),
    .o({\u2_Display/lt104_c27 ,open_n1536}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_27  (
    .a(\u2_Display/n3195 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c27 ),
    .o({\u2_Display/lt104_c28 ,open_n1537}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_28  (
    .a(\u2_Display/n3194 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c28 ),
    .o({\u2_Display/lt104_c29 ,open_n1538}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_29  (
    .a(\u2_Display/n3193 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c29 ),
    .o({\u2_Display/lt104_c30 ,open_n1539}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_3  (
    .a(\u2_Display/n3219 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c3 ),
    .o({\u2_Display/lt104_c4 ,open_n1540}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_30  (
    .a(\u2_Display/n3192 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c30 ),
    .o({\u2_Display/lt104_c31 ,open_n1541}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_31  (
    .a(\u2_Display/n3191 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c31 ),
    .o({\u2_Display/lt104_c32 ,open_n1542}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_4  (
    .a(\u2_Display/n3218 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c4 ),
    .o({\u2_Display/lt104_c5 ,open_n1543}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_5  (
    .a(\u2_Display/n3217 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c5 ),
    .o({\u2_Display/lt104_c6 ,open_n1544}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_6  (
    .a(\u2_Display/n3216 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c6 ),
    .o({\u2_Display/lt104_c7 ,open_n1545}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_7  (
    .a(\u2_Display/n3215 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c7 ),
    .o({\u2_Display/lt104_c8 ,open_n1546}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_8  (
    .a(\u2_Display/n3214 ),
    .b(1'b0),
    .c(\u2_Display/lt104_c8 ),
    .o({\u2_Display/lt104_c9 ,open_n1547}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_9  (
    .a(\u2_Display/n3213 ),
    .b(1'b1),
    .c(\u2_Display/lt104_c9 ),
    .o({\u2_Display/lt104_c10 ,open_n1548}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt104_cin  (
    .a(1'b0),
    .o({\u2_Display/lt104_c0 ,open_n1551}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt104_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt104_c32 ),
    .o({open_n1552,\u2_Display/n3223 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_0  (
    .a(\u2_Display/n3257 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c0 ),
    .o({\u2_Display/lt105_c1 ,open_n1553}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_1  (
    .a(\u2_Display/n3256 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c1 ),
    .o({\u2_Display/lt105_c2 ,open_n1554}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_10  (
    .a(\u2_Display/n3247 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c10 ),
    .o({\u2_Display/lt105_c11 ,open_n1555}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_11  (
    .a(\u2_Display/n3246 ),
    .b(1'b1),
    .c(\u2_Display/lt105_c11 ),
    .o({\u2_Display/lt105_c12 ,open_n1556}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_12  (
    .a(\u2_Display/n3245 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c12 ),
    .o({\u2_Display/lt105_c13 ,open_n1557}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_13  (
    .a(\u2_Display/n3244 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c13 ),
    .o({\u2_Display/lt105_c14 ,open_n1558}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_14  (
    .a(\u2_Display/n3243 ),
    .b(1'b1),
    .c(\u2_Display/lt105_c14 ),
    .o({\u2_Display/lt105_c15 ,open_n1559}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_15  (
    .a(\u2_Display/n3242 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c15 ),
    .o({\u2_Display/lt105_c16 ,open_n1560}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_16  (
    .a(\u2_Display/n3241 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c16 ),
    .o({\u2_Display/lt105_c17 ,open_n1561}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_17  (
    .a(\u2_Display/n3240 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c17 ),
    .o({\u2_Display/lt105_c18 ,open_n1562}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_18  (
    .a(\u2_Display/n3239 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c18 ),
    .o({\u2_Display/lt105_c19 ,open_n1563}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_19  (
    .a(\u2_Display/n3238 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c19 ),
    .o({\u2_Display/lt105_c20 ,open_n1564}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_2  (
    .a(\u2_Display/n3255 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c2 ),
    .o({\u2_Display/lt105_c3 ,open_n1565}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_20  (
    .a(\u2_Display/n3237 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c20 ),
    .o({\u2_Display/lt105_c21 ,open_n1566}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_21  (
    .a(\u2_Display/n3236 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c21 ),
    .o({\u2_Display/lt105_c22 ,open_n1567}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_22  (
    .a(\u2_Display/n3235 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c22 ),
    .o({\u2_Display/lt105_c23 ,open_n1568}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_23  (
    .a(\u2_Display/n3234 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c23 ),
    .o({\u2_Display/lt105_c24 ,open_n1569}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_24  (
    .a(\u2_Display/n3233 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c24 ),
    .o({\u2_Display/lt105_c25 ,open_n1570}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_25  (
    .a(\u2_Display/n3232 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c25 ),
    .o({\u2_Display/lt105_c26 ,open_n1571}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_26  (
    .a(\u2_Display/n3231 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c26 ),
    .o({\u2_Display/lt105_c27 ,open_n1572}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_27  (
    .a(\u2_Display/n3230 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c27 ),
    .o({\u2_Display/lt105_c28 ,open_n1573}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_28  (
    .a(\u2_Display/n3229 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c28 ),
    .o({\u2_Display/lt105_c29 ,open_n1574}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_29  (
    .a(\u2_Display/n3228 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c29 ),
    .o({\u2_Display/lt105_c30 ,open_n1575}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_3  (
    .a(\u2_Display/n3254 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c3 ),
    .o({\u2_Display/lt105_c4 ,open_n1576}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_30  (
    .a(\u2_Display/n3227 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c30 ),
    .o({\u2_Display/lt105_c31 ,open_n1577}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_31  (
    .a(\u2_Display/n3226 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c31 ),
    .o({\u2_Display/lt105_c32 ,open_n1578}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_4  (
    .a(\u2_Display/n3253 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c4 ),
    .o({\u2_Display/lt105_c5 ,open_n1579}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_5  (
    .a(\u2_Display/n3252 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c5 ),
    .o({\u2_Display/lt105_c6 ,open_n1580}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_6  (
    .a(\u2_Display/n3251 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c6 ),
    .o({\u2_Display/lt105_c7 ,open_n1581}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_7  (
    .a(\u2_Display/n3250 ),
    .b(1'b0),
    .c(\u2_Display/lt105_c7 ),
    .o({\u2_Display/lt105_c8 ,open_n1582}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_8  (
    .a(\u2_Display/n3249 ),
    .b(1'b1),
    .c(\u2_Display/lt105_c8 ),
    .o({\u2_Display/lt105_c9 ,open_n1583}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_9  (
    .a(\u2_Display/n3248 ),
    .b(1'b1),
    .c(\u2_Display/lt105_c9 ),
    .o({\u2_Display/lt105_c10 ,open_n1584}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt105_cin  (
    .a(1'b0),
    .o({\u2_Display/lt105_c0 ,open_n1587}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt105_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt105_c32 ),
    .o({open_n1588,\u2_Display/n3258 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_0  (
    .a(\u2_Display/n3292 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c0 ),
    .o({\u2_Display/lt106_c1 ,open_n1589}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_1  (
    .a(\u2_Display/n3291 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c1 ),
    .o({\u2_Display/lt106_c2 ,open_n1590}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_10  (
    .a(\u2_Display/n3282 ),
    .b(1'b1),
    .c(\u2_Display/lt106_c10 ),
    .o({\u2_Display/lt106_c11 ,open_n1591}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_11  (
    .a(\u2_Display/n3281 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c11 ),
    .o({\u2_Display/lt106_c12 ,open_n1592}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_12  (
    .a(\u2_Display/n3280 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c12 ),
    .o({\u2_Display/lt106_c13 ,open_n1593}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_13  (
    .a(\u2_Display/n3279 ),
    .b(1'b1),
    .c(\u2_Display/lt106_c13 ),
    .o({\u2_Display/lt106_c14 ,open_n1594}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_14  (
    .a(\u2_Display/n3278 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c14 ),
    .o({\u2_Display/lt106_c15 ,open_n1595}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_15  (
    .a(\u2_Display/n3277 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c15 ),
    .o({\u2_Display/lt106_c16 ,open_n1596}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_16  (
    .a(\u2_Display/n3276 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c16 ),
    .o({\u2_Display/lt106_c17 ,open_n1597}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_17  (
    .a(\u2_Display/n3275 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c17 ),
    .o({\u2_Display/lt106_c18 ,open_n1598}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_18  (
    .a(\u2_Display/n3274 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c18 ),
    .o({\u2_Display/lt106_c19 ,open_n1599}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_19  (
    .a(\u2_Display/n3273 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c19 ),
    .o({\u2_Display/lt106_c20 ,open_n1600}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_2  (
    .a(\u2_Display/n3290 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c2 ),
    .o({\u2_Display/lt106_c3 ,open_n1601}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_20  (
    .a(\u2_Display/n3272 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c20 ),
    .o({\u2_Display/lt106_c21 ,open_n1602}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_21  (
    .a(\u2_Display/n3271 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c21 ),
    .o({\u2_Display/lt106_c22 ,open_n1603}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_22  (
    .a(\u2_Display/n3270 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c22 ),
    .o({\u2_Display/lt106_c23 ,open_n1604}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_23  (
    .a(\u2_Display/n3269 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c23 ),
    .o({\u2_Display/lt106_c24 ,open_n1605}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_24  (
    .a(\u2_Display/n3268 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c24 ),
    .o({\u2_Display/lt106_c25 ,open_n1606}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_25  (
    .a(\u2_Display/n3267 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c25 ),
    .o({\u2_Display/lt106_c26 ,open_n1607}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_26  (
    .a(\u2_Display/n3266 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c26 ),
    .o({\u2_Display/lt106_c27 ,open_n1608}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_27  (
    .a(\u2_Display/n3265 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c27 ),
    .o({\u2_Display/lt106_c28 ,open_n1609}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_28  (
    .a(\u2_Display/n3264 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c28 ),
    .o({\u2_Display/lt106_c29 ,open_n1610}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_29  (
    .a(\u2_Display/n3263 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c29 ),
    .o({\u2_Display/lt106_c30 ,open_n1611}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_3  (
    .a(\u2_Display/n3289 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c3 ),
    .o({\u2_Display/lt106_c4 ,open_n1612}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_30  (
    .a(\u2_Display/n3262 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c30 ),
    .o({\u2_Display/lt106_c31 ,open_n1613}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_31  (
    .a(\u2_Display/n3261 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c31 ),
    .o({\u2_Display/lt106_c32 ,open_n1614}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_4  (
    .a(\u2_Display/n3288 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c4 ),
    .o({\u2_Display/lt106_c5 ,open_n1615}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_5  (
    .a(\u2_Display/n3287 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c5 ),
    .o({\u2_Display/lt106_c6 ,open_n1616}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_6  (
    .a(\u2_Display/n3286 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c6 ),
    .o({\u2_Display/lt106_c7 ,open_n1617}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_7  (
    .a(\u2_Display/n3285 ),
    .b(1'b1),
    .c(\u2_Display/lt106_c7 ),
    .o({\u2_Display/lt106_c8 ,open_n1618}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_8  (
    .a(\u2_Display/n3284 ),
    .b(1'b1),
    .c(\u2_Display/lt106_c8 ),
    .o({\u2_Display/lt106_c9 ,open_n1619}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_9  (
    .a(\u2_Display/n3283 ),
    .b(1'b0),
    .c(\u2_Display/lt106_c9 ),
    .o({\u2_Display/lt106_c10 ,open_n1620}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt106_cin  (
    .a(1'b0),
    .o({\u2_Display/lt106_c0 ,open_n1623}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt106_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt106_c32 ),
    .o({open_n1624,\u2_Display/n3293 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_0  (
    .a(\u2_Display/n3327 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c0 ),
    .o({\u2_Display/lt107_c1 ,open_n1625}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_1  (
    .a(\u2_Display/n3326 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c1 ),
    .o({\u2_Display/lt107_c2 ,open_n1626}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_10  (
    .a(\u2_Display/n3317 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c10 ),
    .o({\u2_Display/lt107_c11 ,open_n1627}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_11  (
    .a(\u2_Display/n3316 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c11 ),
    .o({\u2_Display/lt107_c12 ,open_n1628}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_12  (
    .a(\u2_Display/n3315 ),
    .b(1'b1),
    .c(\u2_Display/lt107_c12 ),
    .o({\u2_Display/lt107_c13 ,open_n1629}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_13  (
    .a(\u2_Display/n3314 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c13 ),
    .o({\u2_Display/lt107_c14 ,open_n1630}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_14  (
    .a(\u2_Display/n3313 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c14 ),
    .o({\u2_Display/lt107_c15 ,open_n1631}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_15  (
    .a(\u2_Display/n3312 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c15 ),
    .o({\u2_Display/lt107_c16 ,open_n1632}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_16  (
    .a(\u2_Display/n3311 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c16 ),
    .o({\u2_Display/lt107_c17 ,open_n1633}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_17  (
    .a(\u2_Display/n3310 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c17 ),
    .o({\u2_Display/lt107_c18 ,open_n1634}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_18  (
    .a(\u2_Display/n3309 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c18 ),
    .o({\u2_Display/lt107_c19 ,open_n1635}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_19  (
    .a(\u2_Display/n3308 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c19 ),
    .o({\u2_Display/lt107_c20 ,open_n1636}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_2  (
    .a(\u2_Display/n3325 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c2 ),
    .o({\u2_Display/lt107_c3 ,open_n1637}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_20  (
    .a(\u2_Display/n3307 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c20 ),
    .o({\u2_Display/lt107_c21 ,open_n1638}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_21  (
    .a(\u2_Display/n3306 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c21 ),
    .o({\u2_Display/lt107_c22 ,open_n1639}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_22  (
    .a(\u2_Display/n3305 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c22 ),
    .o({\u2_Display/lt107_c23 ,open_n1640}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_23  (
    .a(\u2_Display/n3304 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c23 ),
    .o({\u2_Display/lt107_c24 ,open_n1641}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_24  (
    .a(\u2_Display/n3303 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c24 ),
    .o({\u2_Display/lt107_c25 ,open_n1642}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_25  (
    .a(\u2_Display/n3302 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c25 ),
    .o({\u2_Display/lt107_c26 ,open_n1643}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_26  (
    .a(\u2_Display/n3301 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c26 ),
    .o({\u2_Display/lt107_c27 ,open_n1644}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_27  (
    .a(\u2_Display/n3300 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c27 ),
    .o({\u2_Display/lt107_c28 ,open_n1645}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_28  (
    .a(\u2_Display/n3299 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c28 ),
    .o({\u2_Display/lt107_c29 ,open_n1646}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_29  (
    .a(\u2_Display/n3298 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c29 ),
    .o({\u2_Display/lt107_c30 ,open_n1647}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_3  (
    .a(\u2_Display/n3324 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c3 ),
    .o({\u2_Display/lt107_c4 ,open_n1648}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_30  (
    .a(\u2_Display/n3297 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c30 ),
    .o({\u2_Display/lt107_c31 ,open_n1649}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_31  (
    .a(\u2_Display/n3296 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c31 ),
    .o({\u2_Display/lt107_c32 ,open_n1650}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_4  (
    .a(\u2_Display/n3323 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c4 ),
    .o({\u2_Display/lt107_c5 ,open_n1651}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_5  (
    .a(\u2_Display/n3322 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c5 ),
    .o({\u2_Display/lt107_c6 ,open_n1652}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_6  (
    .a(\u2_Display/n3321 ),
    .b(1'b1),
    .c(\u2_Display/lt107_c6 ),
    .o({\u2_Display/lt107_c7 ,open_n1653}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_7  (
    .a(\u2_Display/n3320 ),
    .b(1'b1),
    .c(\u2_Display/lt107_c7 ),
    .o({\u2_Display/lt107_c8 ,open_n1654}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_8  (
    .a(\u2_Display/n3319 ),
    .b(1'b0),
    .c(\u2_Display/lt107_c8 ),
    .o({\u2_Display/lt107_c9 ,open_n1655}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_9  (
    .a(\u2_Display/n3318 ),
    .b(1'b1),
    .c(\u2_Display/lt107_c9 ),
    .o({\u2_Display/lt107_c10 ,open_n1656}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt107_cin  (
    .a(1'b0),
    .o({\u2_Display/lt107_c0 ,open_n1659}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt107_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt107_c32 ),
    .o({open_n1660,\u2_Display/n3328 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_0  (
    .a(\u2_Display/n3362 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c0 ),
    .o({\u2_Display/lt108_c1 ,open_n1661}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_1  (
    .a(\u2_Display/n3361 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c1 ),
    .o({\u2_Display/lt108_c2 ,open_n1662}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_10  (
    .a(\u2_Display/n3352 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c10 ),
    .o({\u2_Display/lt108_c11 ,open_n1663}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_11  (
    .a(\u2_Display/n3351 ),
    .b(1'b1),
    .c(\u2_Display/lt108_c11 ),
    .o({\u2_Display/lt108_c12 ,open_n1664}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_12  (
    .a(\u2_Display/n3350 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c12 ),
    .o({\u2_Display/lt108_c13 ,open_n1665}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_13  (
    .a(\u2_Display/n3349 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c13 ),
    .o({\u2_Display/lt108_c14 ,open_n1666}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_14  (
    .a(\u2_Display/n3348 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c14 ),
    .o({\u2_Display/lt108_c15 ,open_n1667}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_15  (
    .a(\u2_Display/n3347 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c15 ),
    .o({\u2_Display/lt108_c16 ,open_n1668}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_16  (
    .a(\u2_Display/n3346 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c16 ),
    .o({\u2_Display/lt108_c17 ,open_n1669}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_17  (
    .a(\u2_Display/n3345 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c17 ),
    .o({\u2_Display/lt108_c18 ,open_n1670}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_18  (
    .a(\u2_Display/n3344 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c18 ),
    .o({\u2_Display/lt108_c19 ,open_n1671}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_19  (
    .a(\u2_Display/n3343 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c19 ),
    .o({\u2_Display/lt108_c20 ,open_n1672}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_2  (
    .a(\u2_Display/n3360 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c2 ),
    .o({\u2_Display/lt108_c3 ,open_n1673}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_20  (
    .a(\u2_Display/n3342 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c20 ),
    .o({\u2_Display/lt108_c21 ,open_n1674}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_21  (
    .a(\u2_Display/n3341 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c21 ),
    .o({\u2_Display/lt108_c22 ,open_n1675}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_22  (
    .a(\u2_Display/n3340 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c22 ),
    .o({\u2_Display/lt108_c23 ,open_n1676}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_23  (
    .a(\u2_Display/n3339 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c23 ),
    .o({\u2_Display/lt108_c24 ,open_n1677}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_24  (
    .a(\u2_Display/n3338 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c24 ),
    .o({\u2_Display/lt108_c25 ,open_n1678}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_25  (
    .a(\u2_Display/n3337 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c25 ),
    .o({\u2_Display/lt108_c26 ,open_n1679}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_26  (
    .a(\u2_Display/n3336 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c26 ),
    .o({\u2_Display/lt108_c27 ,open_n1680}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_27  (
    .a(\u2_Display/n3335 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c27 ),
    .o({\u2_Display/lt108_c28 ,open_n1681}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_28  (
    .a(\u2_Display/n3334 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c28 ),
    .o({\u2_Display/lt108_c29 ,open_n1682}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_29  (
    .a(\u2_Display/n3333 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c29 ),
    .o({\u2_Display/lt108_c30 ,open_n1683}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_3  (
    .a(\u2_Display/n3359 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c3 ),
    .o({\u2_Display/lt108_c4 ,open_n1684}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_30  (
    .a(\u2_Display/n3332 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c30 ),
    .o({\u2_Display/lt108_c31 ,open_n1685}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_31  (
    .a(\u2_Display/n3331 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c31 ),
    .o({\u2_Display/lt108_c32 ,open_n1686}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_4  (
    .a(\u2_Display/n3358 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c4 ),
    .o({\u2_Display/lt108_c5 ,open_n1687}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_5  (
    .a(\u2_Display/n3357 ),
    .b(1'b1),
    .c(\u2_Display/lt108_c5 ),
    .o({\u2_Display/lt108_c6 ,open_n1688}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_6  (
    .a(\u2_Display/n3356 ),
    .b(1'b1),
    .c(\u2_Display/lt108_c6 ),
    .o({\u2_Display/lt108_c7 ,open_n1689}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_7  (
    .a(\u2_Display/n3355 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c7 ),
    .o({\u2_Display/lt108_c8 ,open_n1690}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_8  (
    .a(\u2_Display/n3354 ),
    .b(1'b1),
    .c(\u2_Display/lt108_c8 ),
    .o({\u2_Display/lt108_c9 ,open_n1691}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_9  (
    .a(\u2_Display/n3353 ),
    .b(1'b0),
    .c(\u2_Display/lt108_c9 ),
    .o({\u2_Display/lt108_c10 ,open_n1692}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt108_cin  (
    .a(1'b0),
    .o({\u2_Display/lt108_c0 ,open_n1695}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt108_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt108_c32 ),
    .o({open_n1696,\u2_Display/n3363 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_0  (
    .a(\u2_Display/n3397 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c0 ),
    .o({\u2_Display/lt109_c1 ,open_n1697}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_1  (
    .a(\u2_Display/n3396 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c1 ),
    .o({\u2_Display/lt109_c2 ,open_n1698}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_10  (
    .a(\u2_Display/n3387 ),
    .b(1'b1),
    .c(\u2_Display/lt109_c10 ),
    .o({\u2_Display/lt109_c11 ,open_n1699}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_11  (
    .a(\u2_Display/n3386 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c11 ),
    .o({\u2_Display/lt109_c12 ,open_n1700}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_12  (
    .a(\u2_Display/n3385 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c12 ),
    .o({\u2_Display/lt109_c13 ,open_n1701}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_13  (
    .a(\u2_Display/n3384 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c13 ),
    .o({\u2_Display/lt109_c14 ,open_n1702}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_14  (
    .a(\u2_Display/n3383 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c14 ),
    .o({\u2_Display/lt109_c15 ,open_n1703}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_15  (
    .a(\u2_Display/n3382 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c15 ),
    .o({\u2_Display/lt109_c16 ,open_n1704}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_16  (
    .a(\u2_Display/n3381 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c16 ),
    .o({\u2_Display/lt109_c17 ,open_n1705}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_17  (
    .a(\u2_Display/n3380 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c17 ),
    .o({\u2_Display/lt109_c18 ,open_n1706}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_18  (
    .a(\u2_Display/n3379 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c18 ),
    .o({\u2_Display/lt109_c19 ,open_n1707}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_19  (
    .a(\u2_Display/n3378 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c19 ),
    .o({\u2_Display/lt109_c20 ,open_n1708}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_2  (
    .a(\u2_Display/n3395 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c2 ),
    .o({\u2_Display/lt109_c3 ,open_n1709}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_20  (
    .a(\u2_Display/n3377 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c20 ),
    .o({\u2_Display/lt109_c21 ,open_n1710}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_21  (
    .a(\u2_Display/n3376 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c21 ),
    .o({\u2_Display/lt109_c22 ,open_n1711}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_22  (
    .a(\u2_Display/n3375 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c22 ),
    .o({\u2_Display/lt109_c23 ,open_n1712}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_23  (
    .a(\u2_Display/n3374 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c23 ),
    .o({\u2_Display/lt109_c24 ,open_n1713}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_24  (
    .a(\u2_Display/n3373 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c24 ),
    .o({\u2_Display/lt109_c25 ,open_n1714}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_25  (
    .a(\u2_Display/n3372 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c25 ),
    .o({\u2_Display/lt109_c26 ,open_n1715}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_26  (
    .a(\u2_Display/n3371 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c26 ),
    .o({\u2_Display/lt109_c27 ,open_n1716}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_27  (
    .a(\u2_Display/n3370 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c27 ),
    .o({\u2_Display/lt109_c28 ,open_n1717}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_28  (
    .a(\u2_Display/n3369 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c28 ),
    .o({\u2_Display/lt109_c29 ,open_n1718}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_29  (
    .a(\u2_Display/n3368 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c29 ),
    .o({\u2_Display/lt109_c30 ,open_n1719}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_3  (
    .a(\u2_Display/n3394 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c3 ),
    .o({\u2_Display/lt109_c4 ,open_n1720}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_30  (
    .a(\u2_Display/n3367 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c30 ),
    .o({\u2_Display/lt109_c31 ,open_n1721}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_31  (
    .a(\u2_Display/n3366 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c31 ),
    .o({\u2_Display/lt109_c32 ,open_n1722}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_4  (
    .a(\u2_Display/n3393 ),
    .b(1'b1),
    .c(\u2_Display/lt109_c4 ),
    .o({\u2_Display/lt109_c5 ,open_n1723}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_5  (
    .a(\u2_Display/n3392 ),
    .b(1'b1),
    .c(\u2_Display/lt109_c5 ),
    .o({\u2_Display/lt109_c6 ,open_n1724}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_6  (
    .a(\u2_Display/n3391 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c6 ),
    .o({\u2_Display/lt109_c7 ,open_n1725}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_7  (
    .a(\u2_Display/n3390 ),
    .b(1'b1),
    .c(\u2_Display/lt109_c7 ),
    .o({\u2_Display/lt109_c8 ,open_n1726}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_8  (
    .a(\u2_Display/n3389 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c8 ),
    .o({\u2_Display/lt109_c9 ,open_n1727}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_9  (
    .a(\u2_Display/n3388 ),
    .b(1'b0),
    .c(\u2_Display/lt109_c9 ),
    .o({\u2_Display/lt109_c10 ,open_n1728}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt109_cin  (
    .a(1'b0),
    .o({\u2_Display/lt109_c0 ,open_n1731}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt109_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt109_c32 ),
    .o({open_n1732,\u2_Display/n3398 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt10_2_0  (
    .a(lcd_ypos[0]),
    .b(\u2_Display/i [0]),
    .c(\u2_Display/lt10_2_c0 ),
    .o({\u2_Display/lt10_2_c1 ,open_n1733}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt10_2_1  (
    .a(lcd_ypos[1]),
    .b(\u2_Display/i [1]),
    .c(\u2_Display/lt10_2_c1 ),
    .o({\u2_Display/lt10_2_c2 ,open_n1734}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt10_2_10  (
    .a(lcd_ypos[10]),
    .b(\u2_Display/n140 [1]),
    .c(\u2_Display/lt10_2_c10 ),
    .o({\u2_Display/lt10_2_c11 ,open_n1735}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt10_2_11  (
    .a(lcd_ypos[11]),
    .b(\u2_Display/add7_2_co ),
    .c(\u2_Display/lt10_2_c11 ),
    .o({\u2_Display/lt10_2_c12 ,open_n1736}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt10_2_2  (
    .a(lcd_ypos[2]),
    .b(\u2_Display/i [2]),
    .c(\u2_Display/lt10_2_c2 ),
    .o({\u2_Display/lt10_2_c3 ,open_n1737}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt10_2_3  (
    .a(lcd_ypos[3]),
    .b(\u2_Display/i [3]),
    .c(\u2_Display/lt10_2_c3 ),
    .o({\u2_Display/lt10_2_c4 ,open_n1738}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt10_2_4  (
    .a(lcd_ypos[4]),
    .b(\u2_Display/i [4]),
    .c(\u2_Display/lt10_2_c4 ),
    .o({\u2_Display/lt10_2_c5 ,open_n1739}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt10_2_5  (
    .a(lcd_ypos[5]),
    .b(\u2_Display/i [5]),
    .c(\u2_Display/lt10_2_c5 ),
    .o({\u2_Display/lt10_2_c6 ,open_n1740}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt10_2_6  (
    .a(lcd_ypos[6]),
    .b(\u2_Display/i [6]),
    .c(\u2_Display/lt10_2_c6 ),
    .o({\u2_Display/lt10_2_c7 ,open_n1741}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt10_2_7  (
    .a(lcd_ypos[7]),
    .b(\u2_Display/i [7]),
    .c(\u2_Display/lt10_2_c7 ),
    .o({\u2_Display/lt10_2_c8 ,open_n1742}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt10_2_8  (
    .a(lcd_ypos[8]),
    .b(\u2_Display/i [8]),
    .c(\u2_Display/lt10_2_c8 ),
    .o({\u2_Display/lt10_2_c9 ,open_n1743}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt10_2_9  (
    .a(lcd_ypos[9]),
    .b(\u2_Display/n140 [0]),
    .c(\u2_Display/lt10_2_c9 ),
    .o({\u2_Display/lt10_2_c10 ,open_n1744}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt10_2_cin  (
    .a(1'b0),
    .o({\u2_Display/lt10_2_c0 ,open_n1747}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt10_2_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt10_2_c12 ),
    .o({open_n1748,\u2_Display/n141 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_0  (
    .a(\u2_Display/n3432 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c0 ),
    .o({\u2_Display/lt110_c1 ,open_n1749}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_1  (
    .a(\u2_Display/n3431 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c1 ),
    .o({\u2_Display/lt110_c2 ,open_n1750}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_10  (
    .a(\u2_Display/n3422 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c10 ),
    .o({\u2_Display/lt110_c11 ,open_n1751}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_11  (
    .a(\u2_Display/n3421 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c11 ),
    .o({\u2_Display/lt110_c12 ,open_n1752}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_12  (
    .a(\u2_Display/n3420 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c12 ),
    .o({\u2_Display/lt110_c13 ,open_n1753}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_13  (
    .a(\u2_Display/n3419 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c13 ),
    .o({\u2_Display/lt110_c14 ,open_n1754}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_14  (
    .a(\u2_Display/n3418 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c14 ),
    .o({\u2_Display/lt110_c15 ,open_n1755}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_15  (
    .a(\u2_Display/n3417 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c15 ),
    .o({\u2_Display/lt110_c16 ,open_n1756}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_16  (
    .a(\u2_Display/n3416 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c16 ),
    .o({\u2_Display/lt110_c17 ,open_n1757}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_17  (
    .a(\u2_Display/n3415 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c17 ),
    .o({\u2_Display/lt110_c18 ,open_n1758}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_18  (
    .a(\u2_Display/n3414 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c18 ),
    .o({\u2_Display/lt110_c19 ,open_n1759}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_19  (
    .a(\u2_Display/n3413 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c19 ),
    .o({\u2_Display/lt110_c20 ,open_n1760}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_2  (
    .a(\u2_Display/n3430 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c2 ),
    .o({\u2_Display/lt110_c3 ,open_n1761}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_20  (
    .a(\u2_Display/n3412 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c20 ),
    .o({\u2_Display/lt110_c21 ,open_n1762}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_21  (
    .a(\u2_Display/n3411 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c21 ),
    .o({\u2_Display/lt110_c22 ,open_n1763}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_22  (
    .a(\u2_Display/n3410 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c22 ),
    .o({\u2_Display/lt110_c23 ,open_n1764}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_23  (
    .a(\u2_Display/n3409 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c23 ),
    .o({\u2_Display/lt110_c24 ,open_n1765}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_24  (
    .a(\u2_Display/n3408 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c24 ),
    .o({\u2_Display/lt110_c25 ,open_n1766}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_25  (
    .a(\u2_Display/n3407 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c25 ),
    .o({\u2_Display/lt110_c26 ,open_n1767}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_26  (
    .a(\u2_Display/n3406 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c26 ),
    .o({\u2_Display/lt110_c27 ,open_n1768}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_27  (
    .a(\u2_Display/n3405 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c27 ),
    .o({\u2_Display/lt110_c28 ,open_n1769}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_28  (
    .a(\u2_Display/n3404 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c28 ),
    .o({\u2_Display/lt110_c29 ,open_n1770}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_29  (
    .a(\u2_Display/n3403 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c29 ),
    .o({\u2_Display/lt110_c30 ,open_n1771}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_3  (
    .a(\u2_Display/n3429 ),
    .b(1'b1),
    .c(\u2_Display/lt110_c3 ),
    .o({\u2_Display/lt110_c4 ,open_n1772}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_30  (
    .a(\u2_Display/n3402 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c30 ),
    .o({\u2_Display/lt110_c31 ,open_n1773}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_31  (
    .a(\u2_Display/n3401 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c31 ),
    .o({\u2_Display/lt110_c32 ,open_n1774}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_4  (
    .a(\u2_Display/n3428 ),
    .b(1'b1),
    .c(\u2_Display/lt110_c4 ),
    .o({\u2_Display/lt110_c5 ,open_n1775}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_5  (
    .a(\u2_Display/n3427 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c5 ),
    .o({\u2_Display/lt110_c6 ,open_n1776}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_6  (
    .a(\u2_Display/n3426 ),
    .b(1'b1),
    .c(\u2_Display/lt110_c6 ),
    .o({\u2_Display/lt110_c7 ,open_n1777}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_7  (
    .a(\u2_Display/n3425 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c7 ),
    .o({\u2_Display/lt110_c8 ,open_n1778}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_8  (
    .a(\u2_Display/n3424 ),
    .b(1'b0),
    .c(\u2_Display/lt110_c8 ),
    .o({\u2_Display/lt110_c9 ,open_n1779}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_9  (
    .a(\u2_Display/n3423 ),
    .b(1'b1),
    .c(\u2_Display/lt110_c9 ),
    .o({\u2_Display/lt110_c10 ,open_n1780}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt110_cin  (
    .a(1'b0),
    .o({\u2_Display/lt110_c0 ,open_n1783}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt110_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt110_c32 ),
    .o({open_n1784,\u2_Display/n3433 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_0  (
    .a(\u2_Display/n143 [0]),
    .b(lcd_ypos[0]),
    .c(\u2_Display/lt11_2_c0 ),
    .o({\u2_Display/lt11_2_c1 ,open_n1785}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_1  (
    .a(\u2_Display/n143 [1]),
    .b(lcd_ypos[1]),
    .c(\u2_Display/lt11_2_c1 ),
    .o({\u2_Display/lt11_2_c2 ,open_n1786}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_10  (
    .a(\u2_Display/n143 [10]),
    .b(lcd_ypos[10]),
    .c(\u2_Display/lt11_2_c10 ),
    .o({\u2_Display/lt11_2_c11 ,open_n1787}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_11  (
    .a(\u2_Display/n143 [31]),
    .b(lcd_ypos[11]),
    .c(\u2_Display/lt11_2_c11 ),
    .o({\u2_Display/lt11_2_c12 ,open_n1788}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_12  (
    .a(\u2_Display/n143 [31]),
    .b(1'b0),
    .c(\u2_Display/lt11_2_c12 ),
    .o({\u2_Display/lt11_2_c13 ,open_n1789}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_2  (
    .a(\u2_Display/n143 [2]),
    .b(lcd_ypos[2]),
    .c(\u2_Display/lt11_2_c2 ),
    .o({\u2_Display/lt11_2_c3 ,open_n1790}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_3  (
    .a(\u2_Display/n143 [3]),
    .b(lcd_ypos[3]),
    .c(\u2_Display/lt11_2_c3 ),
    .o({\u2_Display/lt11_2_c4 ,open_n1791}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_4  (
    .a(\u2_Display/n143 [4]),
    .b(lcd_ypos[4]),
    .c(\u2_Display/lt11_2_c4 ),
    .o({\u2_Display/lt11_2_c5 ,open_n1792}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_5  (
    .a(\u2_Display/n143 [5]),
    .b(lcd_ypos[5]),
    .c(\u2_Display/lt11_2_c5 ),
    .o({\u2_Display/lt11_2_c6 ,open_n1793}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_6  (
    .a(\u2_Display/n143 [6]),
    .b(lcd_ypos[6]),
    .c(\u2_Display/lt11_2_c6 ),
    .o({\u2_Display/lt11_2_c7 ,open_n1794}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_7  (
    .a(\u2_Display/n143 [7]),
    .b(lcd_ypos[7]),
    .c(\u2_Display/lt11_2_c7 ),
    .o({\u2_Display/lt11_2_c8 ,open_n1795}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_8  (
    .a(\u2_Display/n143 [8]),
    .b(lcd_ypos[8]),
    .c(\u2_Display/lt11_2_c8 ),
    .o({\u2_Display/lt11_2_c9 ,open_n1796}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_9  (
    .a(\u2_Display/n143 [9]),
    .b(lcd_ypos[9]),
    .c(\u2_Display/lt11_2_c9 ),
    .o({\u2_Display/lt11_2_c10 ,open_n1797}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt11_2_cin  (
    .a(1'b0),
    .o({\u2_Display/lt11_2_c0 ,open_n1800}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt11_2_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt11_2_c13 ),
    .o({open_n1801,\u2_Display/n144 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_0  (
    .a(\u2_Display/counta [0]),
    .b(1'b0),
    .c(\u2_Display/lt121_c0 ),
    .o({\u2_Display/lt121_c1 ,open_n1802}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_1  (
    .a(\u2_Display/counta [1]),
    .b(1'b0),
    .c(\u2_Display/lt121_c1 ),
    .o({\u2_Display/lt121_c2 ,open_n1803}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_10  (
    .a(\u2_Display/counta [10]),
    .b(1'b0),
    .c(\u2_Display/lt121_c10 ),
    .o({\u2_Display/lt121_c11 ,open_n1804}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_11  (
    .a(\u2_Display/counta [11]),
    .b(1'b0),
    .c(\u2_Display/lt121_c11 ),
    .o({\u2_Display/lt121_c12 ,open_n1805}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_12  (
    .a(\u2_Display/counta [12]),
    .b(1'b0),
    .c(\u2_Display/lt121_c12 ),
    .o({\u2_Display/lt121_c13 ,open_n1806}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_13  (
    .a(\u2_Display/counta [13]),
    .b(1'b0),
    .c(\u2_Display/lt121_c13 ),
    .o({\u2_Display/lt121_c14 ,open_n1807}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_14  (
    .a(\u2_Display/counta [14]),
    .b(1'b0),
    .c(\u2_Display/lt121_c14 ),
    .o({\u2_Display/lt121_c15 ,open_n1808}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_15  (
    .a(\u2_Display/counta [15]),
    .b(1'b0),
    .c(\u2_Display/lt121_c15 ),
    .o({\u2_Display/lt121_c16 ,open_n1809}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_16  (
    .a(\u2_Display/counta [16]),
    .b(1'b0),
    .c(\u2_Display/lt121_c16 ),
    .o({\u2_Display/lt121_c17 ,open_n1810}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_17  (
    .a(\u2_Display/counta [17]),
    .b(1'b0),
    .c(\u2_Display/lt121_c17 ),
    .o({\u2_Display/lt121_c18 ,open_n1811}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_18  (
    .a(\u2_Display/counta [18]),
    .b(1'b0),
    .c(\u2_Display/lt121_c18 ),
    .o({\u2_Display/lt121_c19 ,open_n1812}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_19  (
    .a(\u2_Display/counta [19]),
    .b(1'b0),
    .c(\u2_Display/lt121_c19 ),
    .o({\u2_Display/lt121_c20 ,open_n1813}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_2  (
    .a(\u2_Display/counta [2]),
    .b(1'b0),
    .c(\u2_Display/lt121_c2 ),
    .o({\u2_Display/lt121_c3 ,open_n1814}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_20  (
    .a(\u2_Display/counta [20]),
    .b(1'b0),
    .c(\u2_Display/lt121_c20 ),
    .o({\u2_Display/lt121_c21 ,open_n1815}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_21  (
    .a(\u2_Display/counta [21]),
    .b(1'b0),
    .c(\u2_Display/lt121_c21 ),
    .o({\u2_Display/lt121_c22 ,open_n1816}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_22  (
    .a(\u2_Display/counta [22]),
    .b(1'b0),
    .c(\u2_Display/lt121_c22 ),
    .o({\u2_Display/lt121_c23 ,open_n1817}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_23  (
    .a(\u2_Display/counta [23]),
    .b(1'b0),
    .c(\u2_Display/lt121_c23 ),
    .o({\u2_Display/lt121_c24 ,open_n1818}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_24  (
    .a(\u2_Display/counta [24]),
    .b(1'b0),
    .c(\u2_Display/lt121_c24 ),
    .o({\u2_Display/lt121_c25 ,open_n1819}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_25  (
    .a(\u2_Display/counta [25]),
    .b(1'b0),
    .c(\u2_Display/lt121_c25 ),
    .o({\u2_Display/lt121_c26 ,open_n1820}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_26  (
    .a(\u2_Display/counta [26]),
    .b(1'b0),
    .c(\u2_Display/lt121_c26 ),
    .o({\u2_Display/lt121_c27 ,open_n1821}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_27  (
    .a(\u2_Display/counta [27]),
    .b(1'b1),
    .c(\u2_Display/lt121_c27 ),
    .o({\u2_Display/lt121_c28 ,open_n1822}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_28  (
    .a(\u2_Display/counta [28]),
    .b(1'b0),
    .c(\u2_Display/lt121_c28 ),
    .o({\u2_Display/lt121_c29 ,open_n1823}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_29  (
    .a(\u2_Display/counta [29]),
    .b(1'b0),
    .c(\u2_Display/lt121_c29 ),
    .o({\u2_Display/lt121_c30 ,open_n1824}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_3  (
    .a(\u2_Display/counta [3]),
    .b(1'b0),
    .c(\u2_Display/lt121_c3 ),
    .o({\u2_Display/lt121_c4 ,open_n1825}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_30  (
    .a(\u2_Display/counta [30]),
    .b(1'b1),
    .c(\u2_Display/lt121_c30 ),
    .o({\u2_Display/lt121_c31 ,open_n1826}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_31  (
    .a(\u2_Display/counta [31]),
    .b(1'b1),
    .c(\u2_Display/lt121_c31 ),
    .o({\u2_Display/lt121_c32 ,open_n1827}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_4  (
    .a(\u2_Display/counta [4]),
    .b(1'b0),
    .c(\u2_Display/lt121_c4 ),
    .o({\u2_Display/lt121_c5 ,open_n1828}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_5  (
    .a(\u2_Display/counta [5]),
    .b(1'b0),
    .c(\u2_Display/lt121_c5 ),
    .o({\u2_Display/lt121_c6 ,open_n1829}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_6  (
    .a(\u2_Display/counta [6]),
    .b(1'b0),
    .c(\u2_Display/lt121_c6 ),
    .o({\u2_Display/lt121_c7 ,open_n1830}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_7  (
    .a(\u2_Display/counta [7]),
    .b(1'b0),
    .c(\u2_Display/lt121_c7 ),
    .o({\u2_Display/lt121_c8 ,open_n1831}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_8  (
    .a(\u2_Display/counta [8]),
    .b(1'b0),
    .c(\u2_Display/lt121_c8 ),
    .o({\u2_Display/lt121_c9 ,open_n1832}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_9  (
    .a(\u2_Display/counta [9]),
    .b(1'b0),
    .c(\u2_Display/lt121_c9 ),
    .o({\u2_Display/lt121_c10 ,open_n1833}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt121_cin  (
    .a(1'b0),
    .o({\u2_Display/lt121_c0 ,open_n1836}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt121_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt121_c32 ),
    .o({open_n1837,\u2_Display/n3786 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_0  (
    .a(\u2_Display/n3820 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c0 ),
    .o({\u2_Display/lt122_c1 ,open_n1838}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_1  (
    .a(\u2_Display/n3819 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c1 ),
    .o({\u2_Display/lt122_c2 ,open_n1839}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_10  (
    .a(\u2_Display/n3810 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c10 ),
    .o({\u2_Display/lt122_c11 ,open_n1840}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_11  (
    .a(\u2_Display/n3809 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c11 ),
    .o({\u2_Display/lt122_c12 ,open_n1841}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_12  (
    .a(\u2_Display/n3808 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c12 ),
    .o({\u2_Display/lt122_c13 ,open_n1842}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_13  (
    .a(\u2_Display/n3807 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c13 ),
    .o({\u2_Display/lt122_c14 ,open_n1843}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_14  (
    .a(\u2_Display/n3806 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c14 ),
    .o({\u2_Display/lt122_c15 ,open_n1844}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_15  (
    .a(\u2_Display/n3805 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c15 ),
    .o({\u2_Display/lt122_c16 ,open_n1845}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_16  (
    .a(\u2_Display/n3804 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c16 ),
    .o({\u2_Display/lt122_c17 ,open_n1846}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_17  (
    .a(\u2_Display/n3803 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c17 ),
    .o({\u2_Display/lt122_c18 ,open_n1847}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_18  (
    .a(\u2_Display/n3802 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c18 ),
    .o({\u2_Display/lt122_c19 ,open_n1848}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_19  (
    .a(\u2_Display/n3801 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c19 ),
    .o({\u2_Display/lt122_c20 ,open_n1849}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_2  (
    .a(\u2_Display/n3818 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c2 ),
    .o({\u2_Display/lt122_c3 ,open_n1850}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_20  (
    .a(\u2_Display/n3800 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c20 ),
    .o({\u2_Display/lt122_c21 ,open_n1851}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_21  (
    .a(\u2_Display/n3799 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c21 ),
    .o({\u2_Display/lt122_c22 ,open_n1852}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_22  (
    .a(\u2_Display/n3798 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c22 ),
    .o({\u2_Display/lt122_c23 ,open_n1853}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_23  (
    .a(\u2_Display/n3797 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c23 ),
    .o({\u2_Display/lt122_c24 ,open_n1854}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_24  (
    .a(\u2_Display/n3796 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c24 ),
    .o({\u2_Display/lt122_c25 ,open_n1855}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_25  (
    .a(\u2_Display/n3795 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c25 ),
    .o({\u2_Display/lt122_c26 ,open_n1856}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_26  (
    .a(\u2_Display/n3794 ),
    .b(1'b1),
    .c(\u2_Display/lt122_c26 ),
    .o({\u2_Display/lt122_c27 ,open_n1857}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_27  (
    .a(\u2_Display/n3793 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c27 ),
    .o({\u2_Display/lt122_c28 ,open_n1858}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_28  (
    .a(\u2_Display/n3792 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c28 ),
    .o({\u2_Display/lt122_c29 ,open_n1859}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_29  (
    .a(\u2_Display/n3791 ),
    .b(1'b1),
    .c(\u2_Display/lt122_c29 ),
    .o({\u2_Display/lt122_c30 ,open_n1860}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_3  (
    .a(\u2_Display/n3817 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c3 ),
    .o({\u2_Display/lt122_c4 ,open_n1861}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_30  (
    .a(\u2_Display/n3790 ),
    .b(1'b1),
    .c(\u2_Display/lt122_c30 ),
    .o({\u2_Display/lt122_c31 ,open_n1862}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_31  (
    .a(\u2_Display/n3789 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c31 ),
    .o({\u2_Display/lt122_c32 ,open_n1863}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_4  (
    .a(\u2_Display/n3816 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c4 ),
    .o({\u2_Display/lt122_c5 ,open_n1864}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_5  (
    .a(\u2_Display/n3815 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c5 ),
    .o({\u2_Display/lt122_c6 ,open_n1865}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_6  (
    .a(\u2_Display/n3814 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c6 ),
    .o({\u2_Display/lt122_c7 ,open_n1866}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_7  (
    .a(\u2_Display/n3813 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c7 ),
    .o({\u2_Display/lt122_c8 ,open_n1867}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_8  (
    .a(\u2_Display/n3812 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c8 ),
    .o({\u2_Display/lt122_c9 ,open_n1868}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_9  (
    .a(\u2_Display/n3811 ),
    .b(1'b0),
    .c(\u2_Display/lt122_c9 ),
    .o({\u2_Display/lt122_c10 ,open_n1869}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt122_cin  (
    .a(1'b0),
    .o({\u2_Display/lt122_c0 ,open_n1872}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt122_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt122_c32 ),
    .o({open_n1873,\u2_Display/n3821 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_0  (
    .a(\u2_Display/n3855 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c0 ),
    .o({\u2_Display/lt123_c1 ,open_n1874}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_1  (
    .a(\u2_Display/n3854 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c1 ),
    .o({\u2_Display/lt123_c2 ,open_n1875}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_10  (
    .a(\u2_Display/n3845 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c10 ),
    .o({\u2_Display/lt123_c11 ,open_n1876}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_11  (
    .a(\u2_Display/n3844 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c11 ),
    .o({\u2_Display/lt123_c12 ,open_n1877}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_12  (
    .a(\u2_Display/n3843 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c12 ),
    .o({\u2_Display/lt123_c13 ,open_n1878}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_13  (
    .a(\u2_Display/n3842 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c13 ),
    .o({\u2_Display/lt123_c14 ,open_n1879}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_14  (
    .a(\u2_Display/n3841 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c14 ),
    .o({\u2_Display/lt123_c15 ,open_n1880}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_15  (
    .a(\u2_Display/n3840 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c15 ),
    .o({\u2_Display/lt123_c16 ,open_n1881}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_16  (
    .a(\u2_Display/n3839 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c16 ),
    .o({\u2_Display/lt123_c17 ,open_n1882}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_17  (
    .a(\u2_Display/n3838 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c17 ),
    .o({\u2_Display/lt123_c18 ,open_n1883}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_18  (
    .a(\u2_Display/n3837 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c18 ),
    .o({\u2_Display/lt123_c19 ,open_n1884}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_19  (
    .a(\u2_Display/n3836 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c19 ),
    .o({\u2_Display/lt123_c20 ,open_n1885}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_2  (
    .a(\u2_Display/n3853 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c2 ),
    .o({\u2_Display/lt123_c3 ,open_n1886}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_20  (
    .a(\u2_Display/n3835 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c20 ),
    .o({\u2_Display/lt123_c21 ,open_n1887}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_21  (
    .a(\u2_Display/n3834 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c21 ),
    .o({\u2_Display/lt123_c22 ,open_n1888}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_22  (
    .a(\u2_Display/n3833 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c22 ),
    .o({\u2_Display/lt123_c23 ,open_n1889}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_23  (
    .a(\u2_Display/n3832 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c23 ),
    .o({\u2_Display/lt123_c24 ,open_n1890}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_24  (
    .a(\u2_Display/n3831 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c24 ),
    .o({\u2_Display/lt123_c25 ,open_n1891}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_25  (
    .a(\u2_Display/n3830 ),
    .b(1'b1),
    .c(\u2_Display/lt123_c25 ),
    .o({\u2_Display/lt123_c26 ,open_n1892}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_26  (
    .a(\u2_Display/n3829 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c26 ),
    .o({\u2_Display/lt123_c27 ,open_n1893}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_27  (
    .a(\u2_Display/n3828 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c27 ),
    .o({\u2_Display/lt123_c28 ,open_n1894}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_28  (
    .a(\u2_Display/n3827 ),
    .b(1'b1),
    .c(\u2_Display/lt123_c28 ),
    .o({\u2_Display/lt123_c29 ,open_n1895}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_29  (
    .a(\u2_Display/n3826 ),
    .b(1'b1),
    .c(\u2_Display/lt123_c29 ),
    .o({\u2_Display/lt123_c30 ,open_n1896}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_3  (
    .a(\u2_Display/n3852 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c3 ),
    .o({\u2_Display/lt123_c4 ,open_n1897}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_30  (
    .a(\u2_Display/n3825 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c30 ),
    .o({\u2_Display/lt123_c31 ,open_n1898}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_31  (
    .a(\u2_Display/n3824 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c31 ),
    .o({\u2_Display/lt123_c32 ,open_n1899}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_4  (
    .a(\u2_Display/n3851 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c4 ),
    .o({\u2_Display/lt123_c5 ,open_n1900}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_5  (
    .a(\u2_Display/n3850 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c5 ),
    .o({\u2_Display/lt123_c6 ,open_n1901}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_6  (
    .a(\u2_Display/n3849 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c6 ),
    .o({\u2_Display/lt123_c7 ,open_n1902}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_7  (
    .a(\u2_Display/n3848 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c7 ),
    .o({\u2_Display/lt123_c8 ,open_n1903}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_8  (
    .a(\u2_Display/n3847 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c8 ),
    .o({\u2_Display/lt123_c9 ,open_n1904}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_9  (
    .a(\u2_Display/n3846 ),
    .b(1'b0),
    .c(\u2_Display/lt123_c9 ),
    .o({\u2_Display/lt123_c10 ,open_n1905}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt123_cin  (
    .a(1'b0),
    .o({\u2_Display/lt123_c0 ,open_n1908}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt123_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt123_c32 ),
    .o({open_n1909,\u2_Display/n3856 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_0  (
    .a(\u2_Display/n3890 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c0 ),
    .o({\u2_Display/lt124_c1 ,open_n1910}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_1  (
    .a(\u2_Display/n3889 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c1 ),
    .o({\u2_Display/lt124_c2 ,open_n1911}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_10  (
    .a(\u2_Display/n3880 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c10 ),
    .o({\u2_Display/lt124_c11 ,open_n1912}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_11  (
    .a(\u2_Display/n3879 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c11 ),
    .o({\u2_Display/lt124_c12 ,open_n1913}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_12  (
    .a(\u2_Display/n3878 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c12 ),
    .o({\u2_Display/lt124_c13 ,open_n1914}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_13  (
    .a(\u2_Display/n3877 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c13 ),
    .o({\u2_Display/lt124_c14 ,open_n1915}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_14  (
    .a(\u2_Display/n3876 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c14 ),
    .o({\u2_Display/lt124_c15 ,open_n1916}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_15  (
    .a(\u2_Display/n3875 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c15 ),
    .o({\u2_Display/lt124_c16 ,open_n1917}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_16  (
    .a(\u2_Display/n3874 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c16 ),
    .o({\u2_Display/lt124_c17 ,open_n1918}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_17  (
    .a(\u2_Display/n3873 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c17 ),
    .o({\u2_Display/lt124_c18 ,open_n1919}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_18  (
    .a(\u2_Display/n3872 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c18 ),
    .o({\u2_Display/lt124_c19 ,open_n1920}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_19  (
    .a(\u2_Display/n3871 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c19 ),
    .o({\u2_Display/lt124_c20 ,open_n1921}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_2  (
    .a(\u2_Display/n3888 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c2 ),
    .o({\u2_Display/lt124_c3 ,open_n1922}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_20  (
    .a(\u2_Display/n3870 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c20 ),
    .o({\u2_Display/lt124_c21 ,open_n1923}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_21  (
    .a(\u2_Display/n3869 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c21 ),
    .o({\u2_Display/lt124_c22 ,open_n1924}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_22  (
    .a(\u2_Display/n3868 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c22 ),
    .o({\u2_Display/lt124_c23 ,open_n1925}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_23  (
    .a(\u2_Display/n3867 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c23 ),
    .o({\u2_Display/lt124_c24 ,open_n1926}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_24  (
    .a(\u2_Display/n3866 ),
    .b(1'b1),
    .c(\u2_Display/lt124_c24 ),
    .o({\u2_Display/lt124_c25 ,open_n1927}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_25  (
    .a(\u2_Display/n3865 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c25 ),
    .o({\u2_Display/lt124_c26 ,open_n1928}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_26  (
    .a(\u2_Display/n3864 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c26 ),
    .o({\u2_Display/lt124_c27 ,open_n1929}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_27  (
    .a(\u2_Display/n3863 ),
    .b(1'b1),
    .c(\u2_Display/lt124_c27 ),
    .o({\u2_Display/lt124_c28 ,open_n1930}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_28  (
    .a(\u2_Display/n3862 ),
    .b(1'b1),
    .c(\u2_Display/lt124_c28 ),
    .o({\u2_Display/lt124_c29 ,open_n1931}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_29  (
    .a(\u2_Display/n3861 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c29 ),
    .o({\u2_Display/lt124_c30 ,open_n1932}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_3  (
    .a(\u2_Display/n3887 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c3 ),
    .o({\u2_Display/lt124_c4 ,open_n1933}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_30  (
    .a(\u2_Display/n3860 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c30 ),
    .o({\u2_Display/lt124_c31 ,open_n1934}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_31  (
    .a(\u2_Display/n3859 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c31 ),
    .o({\u2_Display/lt124_c32 ,open_n1935}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_4  (
    .a(\u2_Display/n3886 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c4 ),
    .o({\u2_Display/lt124_c5 ,open_n1936}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_5  (
    .a(\u2_Display/n3885 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c5 ),
    .o({\u2_Display/lt124_c6 ,open_n1937}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_6  (
    .a(\u2_Display/n3884 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c6 ),
    .o({\u2_Display/lt124_c7 ,open_n1938}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_7  (
    .a(\u2_Display/n3883 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c7 ),
    .o({\u2_Display/lt124_c8 ,open_n1939}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_8  (
    .a(\u2_Display/n3882 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c8 ),
    .o({\u2_Display/lt124_c9 ,open_n1940}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_9  (
    .a(\u2_Display/n3881 ),
    .b(1'b0),
    .c(\u2_Display/lt124_c9 ),
    .o({\u2_Display/lt124_c10 ,open_n1941}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt124_cin  (
    .a(1'b0),
    .o({\u2_Display/lt124_c0 ,open_n1944}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt124_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt124_c32 ),
    .o({open_n1945,\u2_Display/n3891 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_0  (
    .a(\u2_Display/n3925 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c0 ),
    .o({\u2_Display/lt125_c1 ,open_n1946}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_1  (
    .a(\u2_Display/n3924 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c1 ),
    .o({\u2_Display/lt125_c2 ,open_n1947}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_10  (
    .a(\u2_Display/n3915 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c10 ),
    .o({\u2_Display/lt125_c11 ,open_n1948}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_11  (
    .a(\u2_Display/n3914 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c11 ),
    .o({\u2_Display/lt125_c12 ,open_n1949}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_12  (
    .a(\u2_Display/n3913 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c12 ),
    .o({\u2_Display/lt125_c13 ,open_n1950}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_13  (
    .a(\u2_Display/n3912 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c13 ),
    .o({\u2_Display/lt125_c14 ,open_n1951}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_14  (
    .a(\u2_Display/n3911 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c14 ),
    .o({\u2_Display/lt125_c15 ,open_n1952}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_15  (
    .a(\u2_Display/n3910 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c15 ),
    .o({\u2_Display/lt125_c16 ,open_n1953}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_16  (
    .a(\u2_Display/n3909 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c16 ),
    .o({\u2_Display/lt125_c17 ,open_n1954}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_17  (
    .a(\u2_Display/n3908 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c17 ),
    .o({\u2_Display/lt125_c18 ,open_n1955}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_18  (
    .a(\u2_Display/n3907 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c18 ),
    .o({\u2_Display/lt125_c19 ,open_n1956}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_19  (
    .a(\u2_Display/n3906 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c19 ),
    .o({\u2_Display/lt125_c20 ,open_n1957}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_2  (
    .a(\u2_Display/n3923 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c2 ),
    .o({\u2_Display/lt125_c3 ,open_n1958}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_20  (
    .a(\u2_Display/n3905 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c20 ),
    .o({\u2_Display/lt125_c21 ,open_n1959}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_21  (
    .a(\u2_Display/n3904 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c21 ),
    .o({\u2_Display/lt125_c22 ,open_n1960}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_22  (
    .a(\u2_Display/n3903 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c22 ),
    .o({\u2_Display/lt125_c23 ,open_n1961}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_23  (
    .a(\u2_Display/n3902 ),
    .b(1'b1),
    .c(\u2_Display/lt125_c23 ),
    .o({\u2_Display/lt125_c24 ,open_n1962}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_24  (
    .a(\u2_Display/n3901 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c24 ),
    .o({\u2_Display/lt125_c25 ,open_n1963}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_25  (
    .a(\u2_Display/n3900 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c25 ),
    .o({\u2_Display/lt125_c26 ,open_n1964}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_26  (
    .a(\u2_Display/n3899 ),
    .b(1'b1),
    .c(\u2_Display/lt125_c26 ),
    .o({\u2_Display/lt125_c27 ,open_n1965}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_27  (
    .a(\u2_Display/n3898 ),
    .b(1'b1),
    .c(\u2_Display/lt125_c27 ),
    .o({\u2_Display/lt125_c28 ,open_n1966}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_28  (
    .a(\u2_Display/n3897 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c28 ),
    .o({\u2_Display/lt125_c29 ,open_n1967}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_29  (
    .a(\u2_Display/n3896 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c29 ),
    .o({\u2_Display/lt125_c30 ,open_n1968}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_3  (
    .a(\u2_Display/n3922 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c3 ),
    .o({\u2_Display/lt125_c4 ,open_n1969}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_30  (
    .a(\u2_Display/n3895 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c30 ),
    .o({\u2_Display/lt125_c31 ,open_n1970}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_31  (
    .a(\u2_Display/n3894 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c31 ),
    .o({\u2_Display/lt125_c32 ,open_n1971}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_4  (
    .a(\u2_Display/n3921 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c4 ),
    .o({\u2_Display/lt125_c5 ,open_n1972}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_5  (
    .a(\u2_Display/n3920 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c5 ),
    .o({\u2_Display/lt125_c6 ,open_n1973}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_6  (
    .a(\u2_Display/n3919 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c6 ),
    .o({\u2_Display/lt125_c7 ,open_n1974}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_7  (
    .a(\u2_Display/n3918 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c7 ),
    .o({\u2_Display/lt125_c8 ,open_n1975}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_8  (
    .a(\u2_Display/n3917 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c8 ),
    .o({\u2_Display/lt125_c9 ,open_n1976}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_9  (
    .a(\u2_Display/n3916 ),
    .b(1'b0),
    .c(\u2_Display/lt125_c9 ),
    .o({\u2_Display/lt125_c10 ,open_n1977}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt125_cin  (
    .a(1'b0),
    .o({\u2_Display/lt125_c0 ,open_n1980}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt125_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt125_c32 ),
    .o({open_n1981,\u2_Display/n3926 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_0  (
    .a(\u2_Display/n3960 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c0 ),
    .o({\u2_Display/lt126_c1 ,open_n1982}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_1  (
    .a(\u2_Display/n3959 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c1 ),
    .o({\u2_Display/lt126_c2 ,open_n1983}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_10  (
    .a(\u2_Display/n3950 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c10 ),
    .o({\u2_Display/lt126_c11 ,open_n1984}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_11  (
    .a(\u2_Display/n3949 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c11 ),
    .o({\u2_Display/lt126_c12 ,open_n1985}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_12  (
    .a(\u2_Display/n3948 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c12 ),
    .o({\u2_Display/lt126_c13 ,open_n1986}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_13  (
    .a(\u2_Display/n3947 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c13 ),
    .o({\u2_Display/lt126_c14 ,open_n1987}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_14  (
    .a(\u2_Display/n3946 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c14 ),
    .o({\u2_Display/lt126_c15 ,open_n1988}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_15  (
    .a(\u2_Display/n3945 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c15 ),
    .o({\u2_Display/lt126_c16 ,open_n1989}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_16  (
    .a(\u2_Display/n3944 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c16 ),
    .o({\u2_Display/lt126_c17 ,open_n1990}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_17  (
    .a(\u2_Display/n3943 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c17 ),
    .o({\u2_Display/lt126_c18 ,open_n1991}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_18  (
    .a(\u2_Display/n3942 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c18 ),
    .o({\u2_Display/lt126_c19 ,open_n1992}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_19  (
    .a(\u2_Display/n3941 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c19 ),
    .o({\u2_Display/lt126_c20 ,open_n1993}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_2  (
    .a(\u2_Display/n3958 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c2 ),
    .o({\u2_Display/lt126_c3 ,open_n1994}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_20  (
    .a(\u2_Display/n3940 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c20 ),
    .o({\u2_Display/lt126_c21 ,open_n1995}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_21  (
    .a(\u2_Display/n3939 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c21 ),
    .o({\u2_Display/lt126_c22 ,open_n1996}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_22  (
    .a(\u2_Display/n3938 ),
    .b(1'b1),
    .c(\u2_Display/lt126_c22 ),
    .o({\u2_Display/lt126_c23 ,open_n1997}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_23  (
    .a(\u2_Display/n3937 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c23 ),
    .o({\u2_Display/lt126_c24 ,open_n1998}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_24  (
    .a(\u2_Display/n3936 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c24 ),
    .o({\u2_Display/lt126_c25 ,open_n1999}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_25  (
    .a(\u2_Display/n3935 ),
    .b(1'b1),
    .c(\u2_Display/lt126_c25 ),
    .o({\u2_Display/lt126_c26 ,open_n2000}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_26  (
    .a(\u2_Display/n3934 ),
    .b(1'b1),
    .c(\u2_Display/lt126_c26 ),
    .o({\u2_Display/lt126_c27 ,open_n2001}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_27  (
    .a(\u2_Display/n3933 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c27 ),
    .o({\u2_Display/lt126_c28 ,open_n2002}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_28  (
    .a(\u2_Display/n3932 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c28 ),
    .o({\u2_Display/lt126_c29 ,open_n2003}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_29  (
    .a(\u2_Display/n3931 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c29 ),
    .o({\u2_Display/lt126_c30 ,open_n2004}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_3  (
    .a(\u2_Display/n3957 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c3 ),
    .o({\u2_Display/lt126_c4 ,open_n2005}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_30  (
    .a(\u2_Display/n3930 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c30 ),
    .o({\u2_Display/lt126_c31 ,open_n2006}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_31  (
    .a(\u2_Display/n3929 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c31 ),
    .o({\u2_Display/lt126_c32 ,open_n2007}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_4  (
    .a(\u2_Display/n3956 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c4 ),
    .o({\u2_Display/lt126_c5 ,open_n2008}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_5  (
    .a(\u2_Display/n3955 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c5 ),
    .o({\u2_Display/lt126_c6 ,open_n2009}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_6  (
    .a(\u2_Display/n3954 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c6 ),
    .o({\u2_Display/lt126_c7 ,open_n2010}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_7  (
    .a(\u2_Display/n3953 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c7 ),
    .o({\u2_Display/lt126_c8 ,open_n2011}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_8  (
    .a(\u2_Display/n3952 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c8 ),
    .o({\u2_Display/lt126_c9 ,open_n2012}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_9  (
    .a(\u2_Display/n3951 ),
    .b(1'b0),
    .c(\u2_Display/lt126_c9 ),
    .o({\u2_Display/lt126_c10 ,open_n2013}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt126_cin  (
    .a(1'b0),
    .o({\u2_Display/lt126_c0 ,open_n2016}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt126_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt126_c32 ),
    .o({open_n2017,\u2_Display/n3961 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_0  (
    .a(\u2_Display/n3995 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c0 ),
    .o({\u2_Display/lt127_c1 ,open_n2018}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_1  (
    .a(\u2_Display/n3994 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c1 ),
    .o({\u2_Display/lt127_c2 ,open_n2019}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_10  (
    .a(\u2_Display/n3985 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c10 ),
    .o({\u2_Display/lt127_c11 ,open_n2020}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_11  (
    .a(\u2_Display/n3984 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c11 ),
    .o({\u2_Display/lt127_c12 ,open_n2021}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_12  (
    .a(\u2_Display/n3983 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c12 ),
    .o({\u2_Display/lt127_c13 ,open_n2022}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_13  (
    .a(\u2_Display/n3982 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c13 ),
    .o({\u2_Display/lt127_c14 ,open_n2023}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_14  (
    .a(\u2_Display/n3981 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c14 ),
    .o({\u2_Display/lt127_c15 ,open_n2024}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_15  (
    .a(\u2_Display/n3980 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c15 ),
    .o({\u2_Display/lt127_c16 ,open_n2025}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_16  (
    .a(\u2_Display/n3979 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c16 ),
    .o({\u2_Display/lt127_c17 ,open_n2026}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_17  (
    .a(\u2_Display/n3978 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c17 ),
    .o({\u2_Display/lt127_c18 ,open_n2027}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_18  (
    .a(\u2_Display/n3977 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c18 ),
    .o({\u2_Display/lt127_c19 ,open_n2028}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_19  (
    .a(\u2_Display/n3976 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c19 ),
    .o({\u2_Display/lt127_c20 ,open_n2029}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_2  (
    .a(\u2_Display/n3993 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c2 ),
    .o({\u2_Display/lt127_c3 ,open_n2030}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_20  (
    .a(\u2_Display/n3975 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c20 ),
    .o({\u2_Display/lt127_c21 ,open_n2031}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_21  (
    .a(\u2_Display/n3974 ),
    .b(1'b1),
    .c(\u2_Display/lt127_c21 ),
    .o({\u2_Display/lt127_c22 ,open_n2032}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_22  (
    .a(\u2_Display/n3973 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c22 ),
    .o({\u2_Display/lt127_c23 ,open_n2033}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_23  (
    .a(\u2_Display/n3972 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c23 ),
    .o({\u2_Display/lt127_c24 ,open_n2034}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_24  (
    .a(\u2_Display/n3971 ),
    .b(1'b1),
    .c(\u2_Display/lt127_c24 ),
    .o({\u2_Display/lt127_c25 ,open_n2035}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_25  (
    .a(\u2_Display/n3970 ),
    .b(1'b1),
    .c(\u2_Display/lt127_c25 ),
    .o({\u2_Display/lt127_c26 ,open_n2036}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_26  (
    .a(\u2_Display/n3969 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c26 ),
    .o({\u2_Display/lt127_c27 ,open_n2037}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_27  (
    .a(\u2_Display/n3968 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c27 ),
    .o({\u2_Display/lt127_c28 ,open_n2038}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_28  (
    .a(\u2_Display/n3967 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c28 ),
    .o({\u2_Display/lt127_c29 ,open_n2039}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_29  (
    .a(\u2_Display/n3966 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c29 ),
    .o({\u2_Display/lt127_c30 ,open_n2040}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_3  (
    .a(\u2_Display/n3992 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c3 ),
    .o({\u2_Display/lt127_c4 ,open_n2041}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_30  (
    .a(\u2_Display/n3965 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c30 ),
    .o({\u2_Display/lt127_c31 ,open_n2042}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_31  (
    .a(\u2_Display/n3964 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c31 ),
    .o({\u2_Display/lt127_c32 ,open_n2043}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_4  (
    .a(\u2_Display/n3991 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c4 ),
    .o({\u2_Display/lt127_c5 ,open_n2044}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_5  (
    .a(\u2_Display/n3990 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c5 ),
    .o({\u2_Display/lt127_c6 ,open_n2045}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_6  (
    .a(\u2_Display/n3989 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c6 ),
    .o({\u2_Display/lt127_c7 ,open_n2046}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_7  (
    .a(\u2_Display/n3988 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c7 ),
    .o({\u2_Display/lt127_c8 ,open_n2047}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_8  (
    .a(\u2_Display/n3987 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c8 ),
    .o({\u2_Display/lt127_c9 ,open_n2048}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_9  (
    .a(\u2_Display/n3986 ),
    .b(1'b0),
    .c(\u2_Display/lt127_c9 ),
    .o({\u2_Display/lt127_c10 ,open_n2049}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt127_cin  (
    .a(1'b0),
    .o({\u2_Display/lt127_c0 ,open_n2052}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt127_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt127_c32 ),
    .o({open_n2053,\u2_Display/n3996 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_0  (
    .a(\u2_Display/n4030 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c0 ),
    .o({\u2_Display/lt128_c1 ,open_n2054}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_1  (
    .a(\u2_Display/n4029 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c1 ),
    .o({\u2_Display/lt128_c2 ,open_n2055}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_10  (
    .a(\u2_Display/n4020 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c10 ),
    .o({\u2_Display/lt128_c11 ,open_n2056}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_11  (
    .a(\u2_Display/n4019 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c11 ),
    .o({\u2_Display/lt128_c12 ,open_n2057}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_12  (
    .a(\u2_Display/n4018 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c12 ),
    .o({\u2_Display/lt128_c13 ,open_n2058}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_13  (
    .a(\u2_Display/n4017 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c13 ),
    .o({\u2_Display/lt128_c14 ,open_n2059}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_14  (
    .a(\u2_Display/n4016 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c14 ),
    .o({\u2_Display/lt128_c15 ,open_n2060}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_15  (
    .a(\u2_Display/n4015 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c15 ),
    .o({\u2_Display/lt128_c16 ,open_n2061}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_16  (
    .a(\u2_Display/n4014 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c16 ),
    .o({\u2_Display/lt128_c17 ,open_n2062}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_17  (
    .a(\u2_Display/n4013 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c17 ),
    .o({\u2_Display/lt128_c18 ,open_n2063}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_18  (
    .a(\u2_Display/n4012 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c18 ),
    .o({\u2_Display/lt128_c19 ,open_n2064}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_19  (
    .a(\u2_Display/n4011 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c19 ),
    .o({\u2_Display/lt128_c20 ,open_n2065}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_2  (
    .a(\u2_Display/n4028 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c2 ),
    .o({\u2_Display/lt128_c3 ,open_n2066}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_20  (
    .a(\u2_Display/n4010 ),
    .b(1'b1),
    .c(\u2_Display/lt128_c20 ),
    .o({\u2_Display/lt128_c21 ,open_n2067}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_21  (
    .a(\u2_Display/n4009 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c21 ),
    .o({\u2_Display/lt128_c22 ,open_n2068}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_22  (
    .a(\u2_Display/n4008 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c22 ),
    .o({\u2_Display/lt128_c23 ,open_n2069}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_23  (
    .a(\u2_Display/n4007 ),
    .b(1'b1),
    .c(\u2_Display/lt128_c23 ),
    .o({\u2_Display/lt128_c24 ,open_n2070}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_24  (
    .a(\u2_Display/n4006 ),
    .b(1'b1),
    .c(\u2_Display/lt128_c24 ),
    .o({\u2_Display/lt128_c25 ,open_n2071}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_25  (
    .a(\u2_Display/n4005 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c25 ),
    .o({\u2_Display/lt128_c26 ,open_n2072}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_26  (
    .a(\u2_Display/n4004 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c26 ),
    .o({\u2_Display/lt128_c27 ,open_n2073}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_27  (
    .a(\u2_Display/n4003 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c27 ),
    .o({\u2_Display/lt128_c28 ,open_n2074}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_28  (
    .a(\u2_Display/n4002 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c28 ),
    .o({\u2_Display/lt128_c29 ,open_n2075}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_29  (
    .a(\u2_Display/n4001 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c29 ),
    .o({\u2_Display/lt128_c30 ,open_n2076}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_3  (
    .a(\u2_Display/n4027 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c3 ),
    .o({\u2_Display/lt128_c4 ,open_n2077}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_30  (
    .a(\u2_Display/n4000 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c30 ),
    .o({\u2_Display/lt128_c31 ,open_n2078}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_31  (
    .a(\u2_Display/n3999 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c31 ),
    .o({\u2_Display/lt128_c32 ,open_n2079}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_4  (
    .a(\u2_Display/n4026 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c4 ),
    .o({\u2_Display/lt128_c5 ,open_n2080}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_5  (
    .a(\u2_Display/n4025 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c5 ),
    .o({\u2_Display/lt128_c6 ,open_n2081}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_6  (
    .a(\u2_Display/n4024 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c6 ),
    .o({\u2_Display/lt128_c7 ,open_n2082}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_7  (
    .a(\u2_Display/n4023 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c7 ),
    .o({\u2_Display/lt128_c8 ,open_n2083}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_8  (
    .a(\u2_Display/n4022 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c8 ),
    .o({\u2_Display/lt128_c9 ,open_n2084}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_9  (
    .a(\u2_Display/n4021 ),
    .b(1'b0),
    .c(\u2_Display/lt128_c9 ),
    .o({\u2_Display/lt128_c10 ,open_n2085}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt128_cin  (
    .a(1'b0),
    .o({\u2_Display/lt128_c0 ,open_n2088}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt128_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt128_c32 ),
    .o({open_n2089,\u2_Display/n4031 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_0  (
    .a(\u2_Display/n4065 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c0 ),
    .o({\u2_Display/lt129_c1 ,open_n2090}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_1  (
    .a(\u2_Display/n4064 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c1 ),
    .o({\u2_Display/lt129_c2 ,open_n2091}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_10  (
    .a(\u2_Display/n4055 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c10 ),
    .o({\u2_Display/lt129_c11 ,open_n2092}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_11  (
    .a(\u2_Display/n4054 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c11 ),
    .o({\u2_Display/lt129_c12 ,open_n2093}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_12  (
    .a(\u2_Display/n4053 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c12 ),
    .o({\u2_Display/lt129_c13 ,open_n2094}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_13  (
    .a(\u2_Display/n4052 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c13 ),
    .o({\u2_Display/lt129_c14 ,open_n2095}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_14  (
    .a(\u2_Display/n4051 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c14 ),
    .o({\u2_Display/lt129_c15 ,open_n2096}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_15  (
    .a(\u2_Display/n4050 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c15 ),
    .o({\u2_Display/lt129_c16 ,open_n2097}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_16  (
    .a(\u2_Display/n4049 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c16 ),
    .o({\u2_Display/lt129_c17 ,open_n2098}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_17  (
    .a(\u2_Display/n4048 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c17 ),
    .o({\u2_Display/lt129_c18 ,open_n2099}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_18  (
    .a(\u2_Display/n4047 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c18 ),
    .o({\u2_Display/lt129_c19 ,open_n2100}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_19  (
    .a(\u2_Display/n4046 ),
    .b(1'b1),
    .c(\u2_Display/lt129_c19 ),
    .o({\u2_Display/lt129_c20 ,open_n2101}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_2  (
    .a(\u2_Display/n4063 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c2 ),
    .o({\u2_Display/lt129_c3 ,open_n2102}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_20  (
    .a(\u2_Display/n4045 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c20 ),
    .o({\u2_Display/lt129_c21 ,open_n2103}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_21  (
    .a(\u2_Display/n4044 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c21 ),
    .o({\u2_Display/lt129_c22 ,open_n2104}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_22  (
    .a(\u2_Display/n4043 ),
    .b(1'b1),
    .c(\u2_Display/lt129_c22 ),
    .o({\u2_Display/lt129_c23 ,open_n2105}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_23  (
    .a(\u2_Display/n4042 ),
    .b(1'b1),
    .c(\u2_Display/lt129_c23 ),
    .o({\u2_Display/lt129_c24 ,open_n2106}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_24  (
    .a(\u2_Display/n4041 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c24 ),
    .o({\u2_Display/lt129_c25 ,open_n2107}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_25  (
    .a(\u2_Display/n4040 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c25 ),
    .o({\u2_Display/lt129_c26 ,open_n2108}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_26  (
    .a(\u2_Display/n4039 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c26 ),
    .o({\u2_Display/lt129_c27 ,open_n2109}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_27  (
    .a(\u2_Display/n4038 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c27 ),
    .o({\u2_Display/lt129_c28 ,open_n2110}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_28  (
    .a(\u2_Display/n4037 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c28 ),
    .o({\u2_Display/lt129_c29 ,open_n2111}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_29  (
    .a(\u2_Display/n4036 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c29 ),
    .o({\u2_Display/lt129_c30 ,open_n2112}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_3  (
    .a(\u2_Display/n4062 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c3 ),
    .o({\u2_Display/lt129_c4 ,open_n2113}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_30  (
    .a(\u2_Display/n4035 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c30 ),
    .o({\u2_Display/lt129_c31 ,open_n2114}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_31  (
    .a(\u2_Display/n4034 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c31 ),
    .o({\u2_Display/lt129_c32 ,open_n2115}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_4  (
    .a(\u2_Display/n4061 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c4 ),
    .o({\u2_Display/lt129_c5 ,open_n2116}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_5  (
    .a(\u2_Display/n4060 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c5 ),
    .o({\u2_Display/lt129_c6 ,open_n2117}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_6  (
    .a(\u2_Display/n4059 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c6 ),
    .o({\u2_Display/lt129_c7 ,open_n2118}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_7  (
    .a(\u2_Display/n4058 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c7 ),
    .o({\u2_Display/lt129_c8 ,open_n2119}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_8  (
    .a(\u2_Display/n4057 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c8 ),
    .o({\u2_Display/lt129_c9 ,open_n2120}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_9  (
    .a(\u2_Display/n4056 ),
    .b(1'b0),
    .c(\u2_Display/lt129_c9 ),
    .o({\u2_Display/lt129_c10 ,open_n2121}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt129_cin  (
    .a(1'b0),
    .o({\u2_Display/lt129_c0 ,open_n2124}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt129_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt129_c32 ),
    .o({open_n2125,\u2_Display/n4066 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_0  (
    .a(\u2_Display/n4100 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c0 ),
    .o({\u2_Display/lt130_c1 ,open_n2126}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_1  (
    .a(\u2_Display/n4099 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c1 ),
    .o({\u2_Display/lt130_c2 ,open_n2127}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_10  (
    .a(\u2_Display/n4090 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c10 ),
    .o({\u2_Display/lt130_c11 ,open_n2128}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_11  (
    .a(\u2_Display/n4089 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c11 ),
    .o({\u2_Display/lt130_c12 ,open_n2129}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_12  (
    .a(\u2_Display/n4088 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c12 ),
    .o({\u2_Display/lt130_c13 ,open_n2130}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_13  (
    .a(\u2_Display/n4087 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c13 ),
    .o({\u2_Display/lt130_c14 ,open_n2131}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_14  (
    .a(\u2_Display/n4086 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c14 ),
    .o({\u2_Display/lt130_c15 ,open_n2132}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_15  (
    .a(\u2_Display/n4085 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c15 ),
    .o({\u2_Display/lt130_c16 ,open_n2133}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_16  (
    .a(\u2_Display/n4084 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c16 ),
    .o({\u2_Display/lt130_c17 ,open_n2134}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_17  (
    .a(\u2_Display/n4083 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c17 ),
    .o({\u2_Display/lt130_c18 ,open_n2135}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_18  (
    .a(\u2_Display/n4082 ),
    .b(1'b1),
    .c(\u2_Display/lt130_c18 ),
    .o({\u2_Display/lt130_c19 ,open_n2136}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_19  (
    .a(\u2_Display/n4081 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c19 ),
    .o({\u2_Display/lt130_c20 ,open_n2137}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_2  (
    .a(\u2_Display/n4098 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c2 ),
    .o({\u2_Display/lt130_c3 ,open_n2138}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_20  (
    .a(\u2_Display/n4080 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c20 ),
    .o({\u2_Display/lt130_c21 ,open_n2139}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_21  (
    .a(\u2_Display/n4079 ),
    .b(1'b1),
    .c(\u2_Display/lt130_c21 ),
    .o({\u2_Display/lt130_c22 ,open_n2140}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_22  (
    .a(\u2_Display/n4078 ),
    .b(1'b1),
    .c(\u2_Display/lt130_c22 ),
    .o({\u2_Display/lt130_c23 ,open_n2141}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_23  (
    .a(\u2_Display/n4077 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c23 ),
    .o({\u2_Display/lt130_c24 ,open_n2142}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_24  (
    .a(\u2_Display/n4076 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c24 ),
    .o({\u2_Display/lt130_c25 ,open_n2143}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_25  (
    .a(\u2_Display/n4075 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c25 ),
    .o({\u2_Display/lt130_c26 ,open_n2144}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_26  (
    .a(\u2_Display/n4074 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c26 ),
    .o({\u2_Display/lt130_c27 ,open_n2145}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_27  (
    .a(\u2_Display/n4073 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c27 ),
    .o({\u2_Display/lt130_c28 ,open_n2146}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_28  (
    .a(\u2_Display/n4072 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c28 ),
    .o({\u2_Display/lt130_c29 ,open_n2147}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_29  (
    .a(\u2_Display/n4071 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c29 ),
    .o({\u2_Display/lt130_c30 ,open_n2148}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_3  (
    .a(\u2_Display/n4097 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c3 ),
    .o({\u2_Display/lt130_c4 ,open_n2149}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_30  (
    .a(\u2_Display/n4070 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c30 ),
    .o({\u2_Display/lt130_c31 ,open_n2150}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_31  (
    .a(\u2_Display/n4069 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c31 ),
    .o({\u2_Display/lt130_c32 ,open_n2151}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_4  (
    .a(\u2_Display/n4096 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c4 ),
    .o({\u2_Display/lt130_c5 ,open_n2152}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_5  (
    .a(\u2_Display/n4095 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c5 ),
    .o({\u2_Display/lt130_c6 ,open_n2153}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_6  (
    .a(\u2_Display/n4094 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c6 ),
    .o({\u2_Display/lt130_c7 ,open_n2154}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_7  (
    .a(\u2_Display/n4093 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c7 ),
    .o({\u2_Display/lt130_c8 ,open_n2155}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_8  (
    .a(\u2_Display/n4092 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c8 ),
    .o({\u2_Display/lt130_c9 ,open_n2156}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_9  (
    .a(\u2_Display/n4091 ),
    .b(1'b0),
    .c(\u2_Display/lt130_c9 ),
    .o({\u2_Display/lt130_c10 ,open_n2157}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt130_cin  (
    .a(1'b0),
    .o({\u2_Display/lt130_c0 ,open_n2160}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt130_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt130_c32 ),
    .o({open_n2161,\u2_Display/n4101 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_0  (
    .a(\u2_Display/n4135 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c0 ),
    .o({\u2_Display/lt131_c1 ,open_n2162}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_1  (
    .a(\u2_Display/n4134 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c1 ),
    .o({\u2_Display/lt131_c2 ,open_n2163}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_10  (
    .a(\u2_Display/n4125 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c10 ),
    .o({\u2_Display/lt131_c11 ,open_n2164}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_11  (
    .a(\u2_Display/n4124 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c11 ),
    .o({\u2_Display/lt131_c12 ,open_n2165}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_12  (
    .a(\u2_Display/n4123 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c12 ),
    .o({\u2_Display/lt131_c13 ,open_n2166}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_13  (
    .a(\u2_Display/n4122 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c13 ),
    .o({\u2_Display/lt131_c14 ,open_n2167}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_14  (
    .a(\u2_Display/n4121 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c14 ),
    .o({\u2_Display/lt131_c15 ,open_n2168}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_15  (
    .a(\u2_Display/n4120 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c15 ),
    .o({\u2_Display/lt131_c16 ,open_n2169}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_16  (
    .a(\u2_Display/n4119 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c16 ),
    .o({\u2_Display/lt131_c17 ,open_n2170}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_17  (
    .a(\u2_Display/n4118 ),
    .b(1'b1),
    .c(\u2_Display/lt131_c17 ),
    .o({\u2_Display/lt131_c18 ,open_n2171}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_18  (
    .a(\u2_Display/n4117 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c18 ),
    .o({\u2_Display/lt131_c19 ,open_n2172}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_19  (
    .a(\u2_Display/n4116 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c19 ),
    .o({\u2_Display/lt131_c20 ,open_n2173}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_2  (
    .a(\u2_Display/n4133 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c2 ),
    .o({\u2_Display/lt131_c3 ,open_n2174}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_20  (
    .a(\u2_Display/n4115 ),
    .b(1'b1),
    .c(\u2_Display/lt131_c20 ),
    .o({\u2_Display/lt131_c21 ,open_n2175}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_21  (
    .a(\u2_Display/n4114 ),
    .b(1'b1),
    .c(\u2_Display/lt131_c21 ),
    .o({\u2_Display/lt131_c22 ,open_n2176}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_22  (
    .a(\u2_Display/n4113 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c22 ),
    .o({\u2_Display/lt131_c23 ,open_n2177}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_23  (
    .a(\u2_Display/n4112 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c23 ),
    .o({\u2_Display/lt131_c24 ,open_n2178}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_24  (
    .a(\u2_Display/n4111 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c24 ),
    .o({\u2_Display/lt131_c25 ,open_n2179}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_25  (
    .a(\u2_Display/n4110 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c25 ),
    .o({\u2_Display/lt131_c26 ,open_n2180}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_26  (
    .a(\u2_Display/n4109 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c26 ),
    .o({\u2_Display/lt131_c27 ,open_n2181}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_27  (
    .a(\u2_Display/n4108 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c27 ),
    .o({\u2_Display/lt131_c28 ,open_n2182}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_28  (
    .a(\u2_Display/n4107 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c28 ),
    .o({\u2_Display/lt131_c29 ,open_n2183}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_29  (
    .a(\u2_Display/n4106 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c29 ),
    .o({\u2_Display/lt131_c30 ,open_n2184}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_3  (
    .a(\u2_Display/n4132 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c3 ),
    .o({\u2_Display/lt131_c4 ,open_n2185}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_30  (
    .a(\u2_Display/n4105 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c30 ),
    .o({\u2_Display/lt131_c31 ,open_n2186}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_31  (
    .a(\u2_Display/n4104 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c31 ),
    .o({\u2_Display/lt131_c32 ,open_n2187}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_4  (
    .a(\u2_Display/n4131 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c4 ),
    .o({\u2_Display/lt131_c5 ,open_n2188}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_5  (
    .a(\u2_Display/n4130 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c5 ),
    .o({\u2_Display/lt131_c6 ,open_n2189}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_6  (
    .a(\u2_Display/n4129 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c6 ),
    .o({\u2_Display/lt131_c7 ,open_n2190}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_7  (
    .a(\u2_Display/n4128 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c7 ),
    .o({\u2_Display/lt131_c8 ,open_n2191}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_8  (
    .a(\u2_Display/n4127 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c8 ),
    .o({\u2_Display/lt131_c9 ,open_n2192}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_9  (
    .a(\u2_Display/n4126 ),
    .b(1'b0),
    .c(\u2_Display/lt131_c9 ),
    .o({\u2_Display/lt131_c10 ,open_n2193}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt131_cin  (
    .a(1'b0),
    .o({\u2_Display/lt131_c0 ,open_n2196}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt131_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt131_c32 ),
    .o({open_n2197,\u2_Display/n4136 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_0  (
    .a(\u2_Display/n4170 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c0 ),
    .o({\u2_Display/lt132_c1 ,open_n2198}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_1  (
    .a(\u2_Display/n4169 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c1 ),
    .o({\u2_Display/lt132_c2 ,open_n2199}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_10  (
    .a(\u2_Display/n4160 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c10 ),
    .o({\u2_Display/lt132_c11 ,open_n2200}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_11  (
    .a(\u2_Display/n4159 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c11 ),
    .o({\u2_Display/lt132_c12 ,open_n2201}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_12  (
    .a(\u2_Display/n4158 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c12 ),
    .o({\u2_Display/lt132_c13 ,open_n2202}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_13  (
    .a(\u2_Display/n4157 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c13 ),
    .o({\u2_Display/lt132_c14 ,open_n2203}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_14  (
    .a(\u2_Display/n4156 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c14 ),
    .o({\u2_Display/lt132_c15 ,open_n2204}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_15  (
    .a(\u2_Display/n4155 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c15 ),
    .o({\u2_Display/lt132_c16 ,open_n2205}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_16  (
    .a(\u2_Display/n4154 ),
    .b(1'b1),
    .c(\u2_Display/lt132_c16 ),
    .o({\u2_Display/lt132_c17 ,open_n2206}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_17  (
    .a(\u2_Display/n4153 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c17 ),
    .o({\u2_Display/lt132_c18 ,open_n2207}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_18  (
    .a(\u2_Display/n4152 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c18 ),
    .o({\u2_Display/lt132_c19 ,open_n2208}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_19  (
    .a(\u2_Display/n4151 ),
    .b(1'b1),
    .c(\u2_Display/lt132_c19 ),
    .o({\u2_Display/lt132_c20 ,open_n2209}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_2  (
    .a(\u2_Display/n4168 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c2 ),
    .o({\u2_Display/lt132_c3 ,open_n2210}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_20  (
    .a(\u2_Display/n4150 ),
    .b(1'b1),
    .c(\u2_Display/lt132_c20 ),
    .o({\u2_Display/lt132_c21 ,open_n2211}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_21  (
    .a(\u2_Display/n4149 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c21 ),
    .o({\u2_Display/lt132_c22 ,open_n2212}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_22  (
    .a(\u2_Display/n4148 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c22 ),
    .o({\u2_Display/lt132_c23 ,open_n2213}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_23  (
    .a(\u2_Display/n4147 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c23 ),
    .o({\u2_Display/lt132_c24 ,open_n2214}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_24  (
    .a(\u2_Display/n4146 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c24 ),
    .o({\u2_Display/lt132_c25 ,open_n2215}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_25  (
    .a(\u2_Display/n4145 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c25 ),
    .o({\u2_Display/lt132_c26 ,open_n2216}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_26  (
    .a(\u2_Display/n4144 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c26 ),
    .o({\u2_Display/lt132_c27 ,open_n2217}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_27  (
    .a(\u2_Display/n4143 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c27 ),
    .o({\u2_Display/lt132_c28 ,open_n2218}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_28  (
    .a(\u2_Display/n4142 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c28 ),
    .o({\u2_Display/lt132_c29 ,open_n2219}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_29  (
    .a(\u2_Display/n4141 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c29 ),
    .o({\u2_Display/lt132_c30 ,open_n2220}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_3  (
    .a(\u2_Display/n4167 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c3 ),
    .o({\u2_Display/lt132_c4 ,open_n2221}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_30  (
    .a(\u2_Display/n4140 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c30 ),
    .o({\u2_Display/lt132_c31 ,open_n2222}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_31  (
    .a(\u2_Display/n4139 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c31 ),
    .o({\u2_Display/lt132_c32 ,open_n2223}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_4  (
    .a(\u2_Display/n4166 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c4 ),
    .o({\u2_Display/lt132_c5 ,open_n2224}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_5  (
    .a(\u2_Display/n4165 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c5 ),
    .o({\u2_Display/lt132_c6 ,open_n2225}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_6  (
    .a(\u2_Display/n4164 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c6 ),
    .o({\u2_Display/lt132_c7 ,open_n2226}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_7  (
    .a(\u2_Display/n4163 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c7 ),
    .o({\u2_Display/lt132_c8 ,open_n2227}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_8  (
    .a(\u2_Display/n4162 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c8 ),
    .o({\u2_Display/lt132_c9 ,open_n2228}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_9  (
    .a(\u2_Display/n4161 ),
    .b(1'b0),
    .c(\u2_Display/lt132_c9 ),
    .o({\u2_Display/lt132_c10 ,open_n2229}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt132_cin  (
    .a(1'b0),
    .o({\u2_Display/lt132_c0 ,open_n2232}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt132_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt132_c32 ),
    .o({open_n2233,\u2_Display/n4171 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_0  (
    .a(\u2_Display/n4205 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c0 ),
    .o({\u2_Display/lt133_c1 ,open_n2234}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_1  (
    .a(\u2_Display/n4204 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c1 ),
    .o({\u2_Display/lt133_c2 ,open_n2235}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_10  (
    .a(\u2_Display/n4195 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c10 ),
    .o({\u2_Display/lt133_c11 ,open_n2236}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_11  (
    .a(\u2_Display/n4194 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c11 ),
    .o({\u2_Display/lt133_c12 ,open_n2237}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_12  (
    .a(\u2_Display/n4193 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c12 ),
    .o({\u2_Display/lt133_c13 ,open_n2238}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_13  (
    .a(\u2_Display/n4192 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c13 ),
    .o({\u2_Display/lt133_c14 ,open_n2239}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_14  (
    .a(\u2_Display/n4191 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c14 ),
    .o({\u2_Display/lt133_c15 ,open_n2240}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_15  (
    .a(\u2_Display/n4190 ),
    .b(1'b1),
    .c(\u2_Display/lt133_c15 ),
    .o({\u2_Display/lt133_c16 ,open_n2241}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_16  (
    .a(\u2_Display/n4189 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c16 ),
    .o({\u2_Display/lt133_c17 ,open_n2242}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_17  (
    .a(\u2_Display/n4188 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c17 ),
    .o({\u2_Display/lt133_c18 ,open_n2243}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_18  (
    .a(\u2_Display/n4187 ),
    .b(1'b1),
    .c(\u2_Display/lt133_c18 ),
    .o({\u2_Display/lt133_c19 ,open_n2244}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_19  (
    .a(\u2_Display/n4186 ),
    .b(1'b1),
    .c(\u2_Display/lt133_c19 ),
    .o({\u2_Display/lt133_c20 ,open_n2245}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_2  (
    .a(\u2_Display/n4203 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c2 ),
    .o({\u2_Display/lt133_c3 ,open_n2246}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_20  (
    .a(\u2_Display/n4185 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c20 ),
    .o({\u2_Display/lt133_c21 ,open_n2247}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_21  (
    .a(\u2_Display/n4184 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c21 ),
    .o({\u2_Display/lt133_c22 ,open_n2248}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_22  (
    .a(\u2_Display/n4183 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c22 ),
    .o({\u2_Display/lt133_c23 ,open_n2249}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_23  (
    .a(\u2_Display/n4182 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c23 ),
    .o({\u2_Display/lt133_c24 ,open_n2250}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_24  (
    .a(\u2_Display/n4181 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c24 ),
    .o({\u2_Display/lt133_c25 ,open_n2251}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_25  (
    .a(\u2_Display/n4180 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c25 ),
    .o({\u2_Display/lt133_c26 ,open_n2252}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_26  (
    .a(\u2_Display/n4179 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c26 ),
    .o({\u2_Display/lt133_c27 ,open_n2253}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_27  (
    .a(\u2_Display/n4178 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c27 ),
    .o({\u2_Display/lt133_c28 ,open_n2254}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_28  (
    .a(\u2_Display/n4177 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c28 ),
    .o({\u2_Display/lt133_c29 ,open_n2255}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_29  (
    .a(\u2_Display/n4176 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c29 ),
    .o({\u2_Display/lt133_c30 ,open_n2256}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_3  (
    .a(\u2_Display/n4202 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c3 ),
    .o({\u2_Display/lt133_c4 ,open_n2257}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_30  (
    .a(\u2_Display/n4175 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c30 ),
    .o({\u2_Display/lt133_c31 ,open_n2258}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_31  (
    .a(\u2_Display/n4174 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c31 ),
    .o({\u2_Display/lt133_c32 ,open_n2259}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_4  (
    .a(\u2_Display/n4201 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c4 ),
    .o({\u2_Display/lt133_c5 ,open_n2260}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_5  (
    .a(\u2_Display/n4200 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c5 ),
    .o({\u2_Display/lt133_c6 ,open_n2261}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_6  (
    .a(\u2_Display/n4199 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c6 ),
    .o({\u2_Display/lt133_c7 ,open_n2262}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_7  (
    .a(\u2_Display/n4198 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c7 ),
    .o({\u2_Display/lt133_c8 ,open_n2263}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_8  (
    .a(\u2_Display/n4197 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c8 ),
    .o({\u2_Display/lt133_c9 ,open_n2264}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_9  (
    .a(\u2_Display/n4196 ),
    .b(1'b0),
    .c(\u2_Display/lt133_c9 ),
    .o({\u2_Display/lt133_c10 ,open_n2265}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt133_cin  (
    .a(1'b0),
    .o({\u2_Display/lt133_c0 ,open_n2268}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt133_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt133_c32 ),
    .o({open_n2269,\u2_Display/n4206 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_0  (
    .a(\u2_Display/n4240 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c0 ),
    .o({\u2_Display/lt134_c1 ,open_n2270}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_1  (
    .a(\u2_Display/n4239 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c1 ),
    .o({\u2_Display/lt134_c2 ,open_n2271}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_10  (
    .a(\u2_Display/n4230 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c10 ),
    .o({\u2_Display/lt134_c11 ,open_n2272}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_11  (
    .a(\u2_Display/n4229 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c11 ),
    .o({\u2_Display/lt134_c12 ,open_n2273}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_12  (
    .a(\u2_Display/n4228 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c12 ),
    .o({\u2_Display/lt134_c13 ,open_n2274}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_13  (
    .a(\u2_Display/n4227 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c13 ),
    .o({\u2_Display/lt134_c14 ,open_n2275}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_14  (
    .a(\u2_Display/n4226 ),
    .b(1'b1),
    .c(\u2_Display/lt134_c14 ),
    .o({\u2_Display/lt134_c15 ,open_n2276}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_15  (
    .a(\u2_Display/n4225 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c15 ),
    .o({\u2_Display/lt134_c16 ,open_n2277}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_16  (
    .a(\u2_Display/n4224 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c16 ),
    .o({\u2_Display/lt134_c17 ,open_n2278}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_17  (
    .a(\u2_Display/n4223 ),
    .b(1'b1),
    .c(\u2_Display/lt134_c17 ),
    .o({\u2_Display/lt134_c18 ,open_n2279}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_18  (
    .a(\u2_Display/n4222 ),
    .b(1'b1),
    .c(\u2_Display/lt134_c18 ),
    .o({\u2_Display/lt134_c19 ,open_n2280}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_19  (
    .a(\u2_Display/n4221 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c19 ),
    .o({\u2_Display/lt134_c20 ,open_n2281}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_2  (
    .a(\u2_Display/n4238 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c2 ),
    .o({\u2_Display/lt134_c3 ,open_n2282}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_20  (
    .a(\u2_Display/n4220 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c20 ),
    .o({\u2_Display/lt134_c21 ,open_n2283}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_21  (
    .a(\u2_Display/n4219 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c21 ),
    .o({\u2_Display/lt134_c22 ,open_n2284}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_22  (
    .a(\u2_Display/n4218 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c22 ),
    .o({\u2_Display/lt134_c23 ,open_n2285}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_23  (
    .a(\u2_Display/n4217 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c23 ),
    .o({\u2_Display/lt134_c24 ,open_n2286}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_24  (
    .a(\u2_Display/n4216 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c24 ),
    .o({\u2_Display/lt134_c25 ,open_n2287}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_25  (
    .a(\u2_Display/n4215 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c25 ),
    .o({\u2_Display/lt134_c26 ,open_n2288}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_26  (
    .a(\u2_Display/n4214 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c26 ),
    .o({\u2_Display/lt134_c27 ,open_n2289}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_27  (
    .a(\u2_Display/n4213 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c27 ),
    .o({\u2_Display/lt134_c28 ,open_n2290}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_28  (
    .a(\u2_Display/n4212 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c28 ),
    .o({\u2_Display/lt134_c29 ,open_n2291}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_29  (
    .a(\u2_Display/n4211 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c29 ),
    .o({\u2_Display/lt134_c30 ,open_n2292}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_3  (
    .a(\u2_Display/n4237 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c3 ),
    .o({\u2_Display/lt134_c4 ,open_n2293}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_30  (
    .a(\u2_Display/n4210 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c30 ),
    .o({\u2_Display/lt134_c31 ,open_n2294}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_31  (
    .a(\u2_Display/n4209 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c31 ),
    .o({\u2_Display/lt134_c32 ,open_n2295}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_4  (
    .a(\u2_Display/n4236 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c4 ),
    .o({\u2_Display/lt134_c5 ,open_n2296}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_5  (
    .a(\u2_Display/n4235 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c5 ),
    .o({\u2_Display/lt134_c6 ,open_n2297}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_6  (
    .a(\u2_Display/n4234 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c6 ),
    .o({\u2_Display/lt134_c7 ,open_n2298}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_7  (
    .a(\u2_Display/n4233 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c7 ),
    .o({\u2_Display/lt134_c8 ,open_n2299}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_8  (
    .a(\u2_Display/n4232 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c8 ),
    .o({\u2_Display/lt134_c9 ,open_n2300}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_9  (
    .a(\u2_Display/n4231 ),
    .b(1'b0),
    .c(\u2_Display/lt134_c9 ),
    .o({\u2_Display/lt134_c10 ,open_n2301}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt134_cin  (
    .a(1'b0),
    .o({\u2_Display/lt134_c0 ,open_n2304}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt134_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt134_c32 ),
    .o({open_n2305,\u2_Display/n4241 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_0  (
    .a(\u2_Display/n4275 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c0 ),
    .o({\u2_Display/lt135_c1 ,open_n2306}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_1  (
    .a(\u2_Display/n4274 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c1 ),
    .o({\u2_Display/lt135_c2 ,open_n2307}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_10  (
    .a(\u2_Display/n4265 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c10 ),
    .o({\u2_Display/lt135_c11 ,open_n2308}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_11  (
    .a(\u2_Display/n4264 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c11 ),
    .o({\u2_Display/lt135_c12 ,open_n2309}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_12  (
    .a(\u2_Display/n4263 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c12 ),
    .o({\u2_Display/lt135_c13 ,open_n2310}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_13  (
    .a(\u2_Display/n4262 ),
    .b(1'b1),
    .c(\u2_Display/lt135_c13 ),
    .o({\u2_Display/lt135_c14 ,open_n2311}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_14  (
    .a(\u2_Display/n4261 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c14 ),
    .o({\u2_Display/lt135_c15 ,open_n2312}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_15  (
    .a(\u2_Display/n4260 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c15 ),
    .o({\u2_Display/lt135_c16 ,open_n2313}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_16  (
    .a(\u2_Display/n4259 ),
    .b(1'b1),
    .c(\u2_Display/lt135_c16 ),
    .o({\u2_Display/lt135_c17 ,open_n2314}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_17  (
    .a(\u2_Display/n4258 ),
    .b(1'b1),
    .c(\u2_Display/lt135_c17 ),
    .o({\u2_Display/lt135_c18 ,open_n2315}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_18  (
    .a(\u2_Display/n4257 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c18 ),
    .o({\u2_Display/lt135_c19 ,open_n2316}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_19  (
    .a(\u2_Display/n4256 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c19 ),
    .o({\u2_Display/lt135_c20 ,open_n2317}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_2  (
    .a(\u2_Display/n4273 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c2 ),
    .o({\u2_Display/lt135_c3 ,open_n2318}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_20  (
    .a(\u2_Display/n4255 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c20 ),
    .o({\u2_Display/lt135_c21 ,open_n2319}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_21  (
    .a(\u2_Display/n4254 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c21 ),
    .o({\u2_Display/lt135_c22 ,open_n2320}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_22  (
    .a(\u2_Display/n4253 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c22 ),
    .o({\u2_Display/lt135_c23 ,open_n2321}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_23  (
    .a(\u2_Display/n4252 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c23 ),
    .o({\u2_Display/lt135_c24 ,open_n2322}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_24  (
    .a(\u2_Display/n4251 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c24 ),
    .o({\u2_Display/lt135_c25 ,open_n2323}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_25  (
    .a(\u2_Display/n4250 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c25 ),
    .o({\u2_Display/lt135_c26 ,open_n2324}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_26  (
    .a(\u2_Display/n4249 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c26 ),
    .o({\u2_Display/lt135_c27 ,open_n2325}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_27  (
    .a(\u2_Display/n4248 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c27 ),
    .o({\u2_Display/lt135_c28 ,open_n2326}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_28  (
    .a(\u2_Display/n4247 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c28 ),
    .o({\u2_Display/lt135_c29 ,open_n2327}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_29  (
    .a(\u2_Display/n4246 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c29 ),
    .o({\u2_Display/lt135_c30 ,open_n2328}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_3  (
    .a(\u2_Display/n4272 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c3 ),
    .o({\u2_Display/lt135_c4 ,open_n2329}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_30  (
    .a(\u2_Display/n4245 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c30 ),
    .o({\u2_Display/lt135_c31 ,open_n2330}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_31  (
    .a(\u2_Display/n4244 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c31 ),
    .o({\u2_Display/lt135_c32 ,open_n2331}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_4  (
    .a(\u2_Display/n4271 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c4 ),
    .o({\u2_Display/lt135_c5 ,open_n2332}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_5  (
    .a(\u2_Display/n4270 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c5 ),
    .o({\u2_Display/lt135_c6 ,open_n2333}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_6  (
    .a(\u2_Display/n4269 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c6 ),
    .o({\u2_Display/lt135_c7 ,open_n2334}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_7  (
    .a(\u2_Display/n4268 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c7 ),
    .o({\u2_Display/lt135_c8 ,open_n2335}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_8  (
    .a(\u2_Display/n4267 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c8 ),
    .o({\u2_Display/lt135_c9 ,open_n2336}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_9  (
    .a(\u2_Display/n4266 ),
    .b(1'b0),
    .c(\u2_Display/lt135_c9 ),
    .o({\u2_Display/lt135_c10 ,open_n2337}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt135_cin  (
    .a(1'b0),
    .o({\u2_Display/lt135_c0 ,open_n2340}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt135_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt135_c32 ),
    .o({open_n2341,\u2_Display/n4276 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_0  (
    .a(\u2_Display/n4310 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c0 ),
    .o({\u2_Display/lt136_c1 ,open_n2342}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_1  (
    .a(\u2_Display/n4309 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c1 ),
    .o({\u2_Display/lt136_c2 ,open_n2343}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_10  (
    .a(\u2_Display/n4300 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c10 ),
    .o({\u2_Display/lt136_c11 ,open_n2344}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_11  (
    .a(\u2_Display/n4299 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c11 ),
    .o({\u2_Display/lt136_c12 ,open_n2345}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_12  (
    .a(\u2_Display/n4298 ),
    .b(1'b1),
    .c(\u2_Display/lt136_c12 ),
    .o({\u2_Display/lt136_c13 ,open_n2346}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_13  (
    .a(\u2_Display/n4297 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c13 ),
    .o({\u2_Display/lt136_c14 ,open_n2347}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_14  (
    .a(\u2_Display/n4296 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c14 ),
    .o({\u2_Display/lt136_c15 ,open_n2348}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_15  (
    .a(\u2_Display/n4295 ),
    .b(1'b1),
    .c(\u2_Display/lt136_c15 ),
    .o({\u2_Display/lt136_c16 ,open_n2349}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_16  (
    .a(\u2_Display/n4294 ),
    .b(1'b1),
    .c(\u2_Display/lt136_c16 ),
    .o({\u2_Display/lt136_c17 ,open_n2350}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_17  (
    .a(\u2_Display/n4293 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c17 ),
    .o({\u2_Display/lt136_c18 ,open_n2351}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_18  (
    .a(\u2_Display/n4292 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c18 ),
    .o({\u2_Display/lt136_c19 ,open_n2352}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_19  (
    .a(\u2_Display/n4291 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c19 ),
    .o({\u2_Display/lt136_c20 ,open_n2353}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_2  (
    .a(\u2_Display/n4308 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c2 ),
    .o({\u2_Display/lt136_c3 ,open_n2354}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_20  (
    .a(\u2_Display/n4290 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c20 ),
    .o({\u2_Display/lt136_c21 ,open_n2355}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_21  (
    .a(\u2_Display/n4289 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c21 ),
    .o({\u2_Display/lt136_c22 ,open_n2356}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_22  (
    .a(\u2_Display/n4288 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c22 ),
    .o({\u2_Display/lt136_c23 ,open_n2357}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_23  (
    .a(\u2_Display/n4287 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c23 ),
    .o({\u2_Display/lt136_c24 ,open_n2358}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_24  (
    .a(\u2_Display/n4286 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c24 ),
    .o({\u2_Display/lt136_c25 ,open_n2359}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_25  (
    .a(\u2_Display/n4285 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c25 ),
    .o({\u2_Display/lt136_c26 ,open_n2360}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_26  (
    .a(\u2_Display/n4284 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c26 ),
    .o({\u2_Display/lt136_c27 ,open_n2361}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_27  (
    .a(\u2_Display/n4283 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c27 ),
    .o({\u2_Display/lt136_c28 ,open_n2362}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_28  (
    .a(\u2_Display/n4282 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c28 ),
    .o({\u2_Display/lt136_c29 ,open_n2363}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_29  (
    .a(\u2_Display/n4281 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c29 ),
    .o({\u2_Display/lt136_c30 ,open_n2364}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_3  (
    .a(\u2_Display/n4307 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c3 ),
    .o({\u2_Display/lt136_c4 ,open_n2365}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_30  (
    .a(\u2_Display/n4280 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c30 ),
    .o({\u2_Display/lt136_c31 ,open_n2366}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_31  (
    .a(\u2_Display/n4279 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c31 ),
    .o({\u2_Display/lt136_c32 ,open_n2367}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_4  (
    .a(\u2_Display/n4306 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c4 ),
    .o({\u2_Display/lt136_c5 ,open_n2368}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_5  (
    .a(\u2_Display/n4305 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c5 ),
    .o({\u2_Display/lt136_c6 ,open_n2369}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_6  (
    .a(\u2_Display/n4304 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c6 ),
    .o({\u2_Display/lt136_c7 ,open_n2370}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_7  (
    .a(\u2_Display/n4303 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c7 ),
    .o({\u2_Display/lt136_c8 ,open_n2371}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_8  (
    .a(\u2_Display/n4302 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c8 ),
    .o({\u2_Display/lt136_c9 ,open_n2372}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_9  (
    .a(\u2_Display/n4301 ),
    .b(1'b0),
    .c(\u2_Display/lt136_c9 ),
    .o({\u2_Display/lt136_c10 ,open_n2373}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt136_cin  (
    .a(1'b0),
    .o({\u2_Display/lt136_c0 ,open_n2376}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt136_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt136_c32 ),
    .o({open_n2377,\u2_Display/n4311 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_0  (
    .a(\u2_Display/n4345 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c0 ),
    .o({\u2_Display/lt137_c1 ,open_n2378}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_1  (
    .a(\u2_Display/n4344 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c1 ),
    .o({\u2_Display/lt137_c2 ,open_n2379}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_10  (
    .a(\u2_Display/n4335 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c10 ),
    .o({\u2_Display/lt137_c11 ,open_n2380}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_11  (
    .a(\u2_Display/n4334 ),
    .b(1'b1),
    .c(\u2_Display/lt137_c11 ),
    .o({\u2_Display/lt137_c12 ,open_n2381}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_12  (
    .a(\u2_Display/n4333 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c12 ),
    .o({\u2_Display/lt137_c13 ,open_n2382}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_13  (
    .a(\u2_Display/n4332 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c13 ),
    .o({\u2_Display/lt137_c14 ,open_n2383}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_14  (
    .a(\u2_Display/n4331 ),
    .b(1'b1),
    .c(\u2_Display/lt137_c14 ),
    .o({\u2_Display/lt137_c15 ,open_n2384}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_15  (
    .a(\u2_Display/n4330 ),
    .b(1'b1),
    .c(\u2_Display/lt137_c15 ),
    .o({\u2_Display/lt137_c16 ,open_n2385}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_16  (
    .a(\u2_Display/n4329 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c16 ),
    .o({\u2_Display/lt137_c17 ,open_n2386}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_17  (
    .a(\u2_Display/n4328 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c17 ),
    .o({\u2_Display/lt137_c18 ,open_n2387}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_18  (
    .a(\u2_Display/n4327 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c18 ),
    .o({\u2_Display/lt137_c19 ,open_n2388}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_19  (
    .a(\u2_Display/n4326 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c19 ),
    .o({\u2_Display/lt137_c20 ,open_n2389}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_2  (
    .a(\u2_Display/n4343 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c2 ),
    .o({\u2_Display/lt137_c3 ,open_n2390}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_20  (
    .a(\u2_Display/n4325 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c20 ),
    .o({\u2_Display/lt137_c21 ,open_n2391}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_21  (
    .a(\u2_Display/n4324 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c21 ),
    .o({\u2_Display/lt137_c22 ,open_n2392}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_22  (
    .a(\u2_Display/n4323 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c22 ),
    .o({\u2_Display/lt137_c23 ,open_n2393}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_23  (
    .a(\u2_Display/n4322 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c23 ),
    .o({\u2_Display/lt137_c24 ,open_n2394}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_24  (
    .a(\u2_Display/n4321 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c24 ),
    .o({\u2_Display/lt137_c25 ,open_n2395}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_25  (
    .a(\u2_Display/n4320 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c25 ),
    .o({\u2_Display/lt137_c26 ,open_n2396}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_26  (
    .a(\u2_Display/n4319 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c26 ),
    .o({\u2_Display/lt137_c27 ,open_n2397}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_27  (
    .a(\u2_Display/n4318 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c27 ),
    .o({\u2_Display/lt137_c28 ,open_n2398}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_28  (
    .a(\u2_Display/n4317 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c28 ),
    .o({\u2_Display/lt137_c29 ,open_n2399}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_29  (
    .a(\u2_Display/n4316 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c29 ),
    .o({\u2_Display/lt137_c30 ,open_n2400}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_3  (
    .a(\u2_Display/n4342 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c3 ),
    .o({\u2_Display/lt137_c4 ,open_n2401}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_30  (
    .a(\u2_Display/n4315 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c30 ),
    .o({\u2_Display/lt137_c31 ,open_n2402}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_31  (
    .a(\u2_Display/n4314 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c31 ),
    .o({\u2_Display/lt137_c32 ,open_n2403}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_4  (
    .a(\u2_Display/n4341 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c4 ),
    .o({\u2_Display/lt137_c5 ,open_n2404}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_5  (
    .a(\u2_Display/n4340 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c5 ),
    .o({\u2_Display/lt137_c6 ,open_n2405}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_6  (
    .a(\u2_Display/n4339 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c6 ),
    .o({\u2_Display/lt137_c7 ,open_n2406}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_7  (
    .a(\u2_Display/n4338 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c7 ),
    .o({\u2_Display/lt137_c8 ,open_n2407}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_8  (
    .a(\u2_Display/n4337 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c8 ),
    .o({\u2_Display/lt137_c9 ,open_n2408}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_9  (
    .a(\u2_Display/n4336 ),
    .b(1'b0),
    .c(\u2_Display/lt137_c9 ),
    .o({\u2_Display/lt137_c10 ,open_n2409}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt137_cin  (
    .a(1'b0),
    .o({\u2_Display/lt137_c0 ,open_n2412}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt137_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt137_c32 ),
    .o({open_n2413,\u2_Display/n4346 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_0  (
    .a(\u2_Display/n4380 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c0 ),
    .o({\u2_Display/lt138_c1 ,open_n2414}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_1  (
    .a(\u2_Display/n4379 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c1 ),
    .o({\u2_Display/lt138_c2 ,open_n2415}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_10  (
    .a(\u2_Display/n4370 ),
    .b(1'b1),
    .c(\u2_Display/lt138_c10 ),
    .o({\u2_Display/lt138_c11 ,open_n2416}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_11  (
    .a(\u2_Display/n4369 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c11 ),
    .o({\u2_Display/lt138_c12 ,open_n2417}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_12  (
    .a(\u2_Display/n4368 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c12 ),
    .o({\u2_Display/lt138_c13 ,open_n2418}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_13  (
    .a(\u2_Display/n4367 ),
    .b(1'b1),
    .c(\u2_Display/lt138_c13 ),
    .o({\u2_Display/lt138_c14 ,open_n2419}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_14  (
    .a(\u2_Display/n4366 ),
    .b(1'b1),
    .c(\u2_Display/lt138_c14 ),
    .o({\u2_Display/lt138_c15 ,open_n2420}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_15  (
    .a(\u2_Display/n4365 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c15 ),
    .o({\u2_Display/lt138_c16 ,open_n2421}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_16  (
    .a(\u2_Display/n4364 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c16 ),
    .o({\u2_Display/lt138_c17 ,open_n2422}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_17  (
    .a(\u2_Display/n4363 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c17 ),
    .o({\u2_Display/lt138_c18 ,open_n2423}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_18  (
    .a(\u2_Display/n4362 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c18 ),
    .o({\u2_Display/lt138_c19 ,open_n2424}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_19  (
    .a(\u2_Display/n4361 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c19 ),
    .o({\u2_Display/lt138_c20 ,open_n2425}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_2  (
    .a(\u2_Display/n4378 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c2 ),
    .o({\u2_Display/lt138_c3 ,open_n2426}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_20  (
    .a(\u2_Display/n4360 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c20 ),
    .o({\u2_Display/lt138_c21 ,open_n2427}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_21  (
    .a(\u2_Display/n4359 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c21 ),
    .o({\u2_Display/lt138_c22 ,open_n2428}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_22  (
    .a(\u2_Display/n4358 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c22 ),
    .o({\u2_Display/lt138_c23 ,open_n2429}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_23  (
    .a(\u2_Display/n4357 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c23 ),
    .o({\u2_Display/lt138_c24 ,open_n2430}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_24  (
    .a(\u2_Display/n4356 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c24 ),
    .o({\u2_Display/lt138_c25 ,open_n2431}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_25  (
    .a(\u2_Display/n4355 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c25 ),
    .o({\u2_Display/lt138_c26 ,open_n2432}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_26  (
    .a(\u2_Display/n4354 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c26 ),
    .o({\u2_Display/lt138_c27 ,open_n2433}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_27  (
    .a(\u2_Display/n4353 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c27 ),
    .o({\u2_Display/lt138_c28 ,open_n2434}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_28  (
    .a(\u2_Display/n4352 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c28 ),
    .o({\u2_Display/lt138_c29 ,open_n2435}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_29  (
    .a(\u2_Display/n4351 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c29 ),
    .o({\u2_Display/lt138_c30 ,open_n2436}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_3  (
    .a(\u2_Display/n4377 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c3 ),
    .o({\u2_Display/lt138_c4 ,open_n2437}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_30  (
    .a(\u2_Display/n4350 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c30 ),
    .o({\u2_Display/lt138_c31 ,open_n2438}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_31  (
    .a(\u2_Display/n4349 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c31 ),
    .o({\u2_Display/lt138_c32 ,open_n2439}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_4  (
    .a(\u2_Display/n4376 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c4 ),
    .o({\u2_Display/lt138_c5 ,open_n2440}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_5  (
    .a(\u2_Display/n4375 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c5 ),
    .o({\u2_Display/lt138_c6 ,open_n2441}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_6  (
    .a(\u2_Display/n4374 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c6 ),
    .o({\u2_Display/lt138_c7 ,open_n2442}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_7  (
    .a(\u2_Display/n4373 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c7 ),
    .o({\u2_Display/lt138_c8 ,open_n2443}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_8  (
    .a(\u2_Display/n4372 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c8 ),
    .o({\u2_Display/lt138_c9 ,open_n2444}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_9  (
    .a(\u2_Display/n4371 ),
    .b(1'b0),
    .c(\u2_Display/lt138_c9 ),
    .o({\u2_Display/lt138_c10 ,open_n2445}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt138_cin  (
    .a(1'b0),
    .o({\u2_Display/lt138_c0 ,open_n2448}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt138_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt138_c32 ),
    .o({open_n2449,\u2_Display/n4381 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_0  (
    .a(\u2_Display/n4415 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c0 ),
    .o({\u2_Display/lt139_c1 ,open_n2450}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_1  (
    .a(\u2_Display/n4414 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c1 ),
    .o({\u2_Display/lt139_c2 ,open_n2451}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_10  (
    .a(\u2_Display/n4405 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c10 ),
    .o({\u2_Display/lt139_c11 ,open_n2452}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_11  (
    .a(\u2_Display/n4404 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c11 ),
    .o({\u2_Display/lt139_c12 ,open_n2453}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_12  (
    .a(\u2_Display/n4403 ),
    .b(1'b1),
    .c(\u2_Display/lt139_c12 ),
    .o({\u2_Display/lt139_c13 ,open_n2454}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_13  (
    .a(\u2_Display/n4402 ),
    .b(1'b1),
    .c(\u2_Display/lt139_c13 ),
    .o({\u2_Display/lt139_c14 ,open_n2455}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_14  (
    .a(\u2_Display/n4401 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c14 ),
    .o({\u2_Display/lt139_c15 ,open_n2456}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_15  (
    .a(\u2_Display/n4400 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c15 ),
    .o({\u2_Display/lt139_c16 ,open_n2457}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_16  (
    .a(\u2_Display/n4399 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c16 ),
    .o({\u2_Display/lt139_c17 ,open_n2458}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_17  (
    .a(\u2_Display/n4398 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c17 ),
    .o({\u2_Display/lt139_c18 ,open_n2459}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_18  (
    .a(\u2_Display/n4397 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c18 ),
    .o({\u2_Display/lt139_c19 ,open_n2460}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_19  (
    .a(\u2_Display/n4396 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c19 ),
    .o({\u2_Display/lt139_c20 ,open_n2461}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_2  (
    .a(\u2_Display/n4413 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c2 ),
    .o({\u2_Display/lt139_c3 ,open_n2462}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_20  (
    .a(\u2_Display/n4395 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c20 ),
    .o({\u2_Display/lt139_c21 ,open_n2463}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_21  (
    .a(\u2_Display/n4394 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c21 ),
    .o({\u2_Display/lt139_c22 ,open_n2464}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_22  (
    .a(\u2_Display/n4393 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c22 ),
    .o({\u2_Display/lt139_c23 ,open_n2465}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_23  (
    .a(\u2_Display/n4392 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c23 ),
    .o({\u2_Display/lt139_c24 ,open_n2466}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_24  (
    .a(\u2_Display/n4391 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c24 ),
    .o({\u2_Display/lt139_c25 ,open_n2467}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_25  (
    .a(\u2_Display/n4390 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c25 ),
    .o({\u2_Display/lt139_c26 ,open_n2468}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_26  (
    .a(\u2_Display/n4389 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c26 ),
    .o({\u2_Display/lt139_c27 ,open_n2469}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_27  (
    .a(\u2_Display/n4388 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c27 ),
    .o({\u2_Display/lt139_c28 ,open_n2470}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_28  (
    .a(\u2_Display/n4387 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c28 ),
    .o({\u2_Display/lt139_c29 ,open_n2471}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_29  (
    .a(\u2_Display/n4386 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c29 ),
    .o({\u2_Display/lt139_c30 ,open_n2472}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_3  (
    .a(\u2_Display/n4412 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c3 ),
    .o({\u2_Display/lt139_c4 ,open_n2473}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_30  (
    .a(\u2_Display/n4385 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c30 ),
    .o({\u2_Display/lt139_c31 ,open_n2474}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_31  (
    .a(\u2_Display/n4384 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c31 ),
    .o({\u2_Display/lt139_c32 ,open_n2475}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_4  (
    .a(\u2_Display/n4411 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c4 ),
    .o({\u2_Display/lt139_c5 ,open_n2476}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_5  (
    .a(\u2_Display/n4410 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c5 ),
    .o({\u2_Display/lt139_c6 ,open_n2477}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_6  (
    .a(\u2_Display/n4409 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c6 ),
    .o({\u2_Display/lt139_c7 ,open_n2478}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_7  (
    .a(\u2_Display/n4408 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c7 ),
    .o({\u2_Display/lt139_c8 ,open_n2479}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_8  (
    .a(\u2_Display/n4407 ),
    .b(1'b0),
    .c(\u2_Display/lt139_c8 ),
    .o({\u2_Display/lt139_c9 ,open_n2480}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_9  (
    .a(\u2_Display/n4406 ),
    .b(1'b1),
    .c(\u2_Display/lt139_c9 ),
    .o({\u2_Display/lt139_c10 ,open_n2481}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt139_cin  (
    .a(1'b0),
    .o({\u2_Display/lt139_c0 ,open_n2484}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt139_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt139_c32 ),
    .o({open_n2485,\u2_Display/n4416 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_0  (
    .a(\u2_Display/n4450 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c0 ),
    .o({\u2_Display/lt140_c1 ,open_n2486}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_1  (
    .a(\u2_Display/n4449 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c1 ),
    .o({\u2_Display/lt140_c2 ,open_n2487}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_10  (
    .a(\u2_Display/n4440 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c10 ),
    .o({\u2_Display/lt140_c11 ,open_n2488}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_11  (
    .a(\u2_Display/n4439 ),
    .b(1'b1),
    .c(\u2_Display/lt140_c11 ),
    .o({\u2_Display/lt140_c12 ,open_n2489}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_12  (
    .a(\u2_Display/n4438 ),
    .b(1'b1),
    .c(\u2_Display/lt140_c12 ),
    .o({\u2_Display/lt140_c13 ,open_n2490}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_13  (
    .a(\u2_Display/n4437 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c13 ),
    .o({\u2_Display/lt140_c14 ,open_n2491}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_14  (
    .a(\u2_Display/n4436 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c14 ),
    .o({\u2_Display/lt140_c15 ,open_n2492}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_15  (
    .a(\u2_Display/n4435 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c15 ),
    .o({\u2_Display/lt140_c16 ,open_n2493}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_16  (
    .a(\u2_Display/n4434 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c16 ),
    .o({\u2_Display/lt140_c17 ,open_n2494}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_17  (
    .a(\u2_Display/n4433 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c17 ),
    .o({\u2_Display/lt140_c18 ,open_n2495}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_18  (
    .a(\u2_Display/n4432 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c18 ),
    .o({\u2_Display/lt140_c19 ,open_n2496}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_19  (
    .a(\u2_Display/n4431 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c19 ),
    .o({\u2_Display/lt140_c20 ,open_n2497}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_2  (
    .a(\u2_Display/n4448 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c2 ),
    .o({\u2_Display/lt140_c3 ,open_n2498}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_20  (
    .a(\u2_Display/n4430 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c20 ),
    .o({\u2_Display/lt140_c21 ,open_n2499}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_21  (
    .a(\u2_Display/n4429 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c21 ),
    .o({\u2_Display/lt140_c22 ,open_n2500}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_22  (
    .a(\u2_Display/n4428 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c22 ),
    .o({\u2_Display/lt140_c23 ,open_n2501}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_23  (
    .a(\u2_Display/n4427 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c23 ),
    .o({\u2_Display/lt140_c24 ,open_n2502}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_24  (
    .a(\u2_Display/n4426 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c24 ),
    .o({\u2_Display/lt140_c25 ,open_n2503}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_25  (
    .a(\u2_Display/n4425 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c25 ),
    .o({\u2_Display/lt140_c26 ,open_n2504}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_26  (
    .a(\u2_Display/n4424 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c26 ),
    .o({\u2_Display/lt140_c27 ,open_n2505}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_27  (
    .a(\u2_Display/n4423 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c27 ),
    .o({\u2_Display/lt140_c28 ,open_n2506}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_28  (
    .a(\u2_Display/n4422 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c28 ),
    .o({\u2_Display/lt140_c29 ,open_n2507}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_29  (
    .a(\u2_Display/n4421 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c29 ),
    .o({\u2_Display/lt140_c30 ,open_n2508}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_3  (
    .a(\u2_Display/n4447 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c3 ),
    .o({\u2_Display/lt140_c4 ,open_n2509}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_30  (
    .a(\u2_Display/n4420 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c30 ),
    .o({\u2_Display/lt140_c31 ,open_n2510}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_31  (
    .a(\u2_Display/n4419 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c31 ),
    .o({\u2_Display/lt140_c32 ,open_n2511}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_4  (
    .a(\u2_Display/n4446 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c4 ),
    .o({\u2_Display/lt140_c5 ,open_n2512}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_5  (
    .a(\u2_Display/n4445 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c5 ),
    .o({\u2_Display/lt140_c6 ,open_n2513}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_6  (
    .a(\u2_Display/n4444 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c6 ),
    .o({\u2_Display/lt140_c7 ,open_n2514}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_7  (
    .a(\u2_Display/n4443 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c7 ),
    .o({\u2_Display/lt140_c8 ,open_n2515}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_8  (
    .a(\u2_Display/n4442 ),
    .b(1'b1),
    .c(\u2_Display/lt140_c8 ),
    .o({\u2_Display/lt140_c9 ,open_n2516}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_9  (
    .a(\u2_Display/n4441 ),
    .b(1'b0),
    .c(\u2_Display/lt140_c9 ),
    .o({\u2_Display/lt140_c10 ,open_n2517}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt140_cin  (
    .a(1'b0),
    .o({\u2_Display/lt140_c0 ,open_n2520}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt140_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt140_c32 ),
    .o({open_n2521,\u2_Display/n4451 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_0  (
    .a(\u2_Display/n4485 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c0 ),
    .o({\u2_Display/lt141_c1 ,open_n2522}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_1  (
    .a(\u2_Display/n4484 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c1 ),
    .o({\u2_Display/lt141_c2 ,open_n2523}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_10  (
    .a(\u2_Display/n4475 ),
    .b(1'b1),
    .c(\u2_Display/lt141_c10 ),
    .o({\u2_Display/lt141_c11 ,open_n2524}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_11  (
    .a(\u2_Display/n4474 ),
    .b(1'b1),
    .c(\u2_Display/lt141_c11 ),
    .o({\u2_Display/lt141_c12 ,open_n2525}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_12  (
    .a(\u2_Display/n4473 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c12 ),
    .o({\u2_Display/lt141_c13 ,open_n2526}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_13  (
    .a(\u2_Display/n4472 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c13 ),
    .o({\u2_Display/lt141_c14 ,open_n2527}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_14  (
    .a(\u2_Display/n4471 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c14 ),
    .o({\u2_Display/lt141_c15 ,open_n2528}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_15  (
    .a(\u2_Display/n4470 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c15 ),
    .o({\u2_Display/lt141_c16 ,open_n2529}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_16  (
    .a(\u2_Display/n4469 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c16 ),
    .o({\u2_Display/lt141_c17 ,open_n2530}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_17  (
    .a(\u2_Display/n4468 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c17 ),
    .o({\u2_Display/lt141_c18 ,open_n2531}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_18  (
    .a(\u2_Display/n4467 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c18 ),
    .o({\u2_Display/lt141_c19 ,open_n2532}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_19  (
    .a(\u2_Display/n4466 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c19 ),
    .o({\u2_Display/lt141_c20 ,open_n2533}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_2  (
    .a(\u2_Display/n4483 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c2 ),
    .o({\u2_Display/lt141_c3 ,open_n2534}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_20  (
    .a(\u2_Display/n4465 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c20 ),
    .o({\u2_Display/lt141_c21 ,open_n2535}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_21  (
    .a(\u2_Display/n4464 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c21 ),
    .o({\u2_Display/lt141_c22 ,open_n2536}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_22  (
    .a(\u2_Display/n4463 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c22 ),
    .o({\u2_Display/lt141_c23 ,open_n2537}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_23  (
    .a(\u2_Display/n4462 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c23 ),
    .o({\u2_Display/lt141_c24 ,open_n2538}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_24  (
    .a(\u2_Display/n4461 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c24 ),
    .o({\u2_Display/lt141_c25 ,open_n2539}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_25  (
    .a(\u2_Display/n4460 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c25 ),
    .o({\u2_Display/lt141_c26 ,open_n2540}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_26  (
    .a(\u2_Display/n4459 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c26 ),
    .o({\u2_Display/lt141_c27 ,open_n2541}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_27  (
    .a(\u2_Display/n4458 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c27 ),
    .o({\u2_Display/lt141_c28 ,open_n2542}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_28  (
    .a(\u2_Display/n4457 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c28 ),
    .o({\u2_Display/lt141_c29 ,open_n2543}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_29  (
    .a(\u2_Display/n4456 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c29 ),
    .o({\u2_Display/lt141_c30 ,open_n2544}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_3  (
    .a(\u2_Display/n4482 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c3 ),
    .o({\u2_Display/lt141_c4 ,open_n2545}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_30  (
    .a(\u2_Display/n4455 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c30 ),
    .o({\u2_Display/lt141_c31 ,open_n2546}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_31  (
    .a(\u2_Display/n4454 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c31 ),
    .o({\u2_Display/lt141_c32 ,open_n2547}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_4  (
    .a(\u2_Display/n4481 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c4 ),
    .o({\u2_Display/lt141_c5 ,open_n2548}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_5  (
    .a(\u2_Display/n4480 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c5 ),
    .o({\u2_Display/lt141_c6 ,open_n2549}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_6  (
    .a(\u2_Display/n4479 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c6 ),
    .o({\u2_Display/lt141_c7 ,open_n2550}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_7  (
    .a(\u2_Display/n4478 ),
    .b(1'b1),
    .c(\u2_Display/lt141_c7 ),
    .o({\u2_Display/lt141_c8 ,open_n2551}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_8  (
    .a(\u2_Display/n4477 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c8 ),
    .o({\u2_Display/lt141_c9 ,open_n2552}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_9  (
    .a(\u2_Display/n4476 ),
    .b(1'b0),
    .c(\u2_Display/lt141_c9 ),
    .o({\u2_Display/lt141_c10 ,open_n2553}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt141_cin  (
    .a(1'b0),
    .o({\u2_Display/lt141_c0 ,open_n2556}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt141_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt141_c32 ),
    .o({open_n2557,\u2_Display/n4486 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_0  (
    .a(\u2_Display/n4520 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c0 ),
    .o({\u2_Display/lt142_c1 ,open_n2558}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_1  (
    .a(\u2_Display/n4519 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c1 ),
    .o({\u2_Display/lt142_c2 ,open_n2559}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_10  (
    .a(\u2_Display/n4510 ),
    .b(1'b1),
    .c(\u2_Display/lt142_c10 ),
    .o({\u2_Display/lt142_c11 ,open_n2560}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_11  (
    .a(\u2_Display/n4509 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c11 ),
    .o({\u2_Display/lt142_c12 ,open_n2561}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_12  (
    .a(\u2_Display/n4508 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c12 ),
    .o({\u2_Display/lt142_c13 ,open_n2562}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_13  (
    .a(\u2_Display/n4507 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c13 ),
    .o({\u2_Display/lt142_c14 ,open_n2563}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_14  (
    .a(\u2_Display/n4506 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c14 ),
    .o({\u2_Display/lt142_c15 ,open_n2564}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_15  (
    .a(\u2_Display/n4505 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c15 ),
    .o({\u2_Display/lt142_c16 ,open_n2565}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_16  (
    .a(\u2_Display/n4504 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c16 ),
    .o({\u2_Display/lt142_c17 ,open_n2566}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_17  (
    .a(\u2_Display/n4503 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c17 ),
    .o({\u2_Display/lt142_c18 ,open_n2567}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_18  (
    .a(\u2_Display/n4502 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c18 ),
    .o({\u2_Display/lt142_c19 ,open_n2568}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_19  (
    .a(\u2_Display/n4501 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c19 ),
    .o({\u2_Display/lt142_c20 ,open_n2569}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_2  (
    .a(\u2_Display/n4518 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c2 ),
    .o({\u2_Display/lt142_c3 ,open_n2570}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_20  (
    .a(\u2_Display/n4500 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c20 ),
    .o({\u2_Display/lt142_c21 ,open_n2571}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_21  (
    .a(\u2_Display/n4499 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c21 ),
    .o({\u2_Display/lt142_c22 ,open_n2572}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_22  (
    .a(\u2_Display/n4498 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c22 ),
    .o({\u2_Display/lt142_c23 ,open_n2573}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_23  (
    .a(\u2_Display/n4497 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c23 ),
    .o({\u2_Display/lt142_c24 ,open_n2574}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_24  (
    .a(\u2_Display/n4496 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c24 ),
    .o({\u2_Display/lt142_c25 ,open_n2575}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_25  (
    .a(\u2_Display/n4495 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c25 ),
    .o({\u2_Display/lt142_c26 ,open_n2576}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_26  (
    .a(\u2_Display/n4494 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c26 ),
    .o({\u2_Display/lt142_c27 ,open_n2577}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_27  (
    .a(\u2_Display/n4493 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c27 ),
    .o({\u2_Display/lt142_c28 ,open_n2578}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_28  (
    .a(\u2_Display/n4492 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c28 ),
    .o({\u2_Display/lt142_c29 ,open_n2579}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_29  (
    .a(\u2_Display/n4491 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c29 ),
    .o({\u2_Display/lt142_c30 ,open_n2580}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_3  (
    .a(\u2_Display/n4517 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c3 ),
    .o({\u2_Display/lt142_c4 ,open_n2581}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_30  (
    .a(\u2_Display/n4490 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c30 ),
    .o({\u2_Display/lt142_c31 ,open_n2582}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_31  (
    .a(\u2_Display/n4489 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c31 ),
    .o({\u2_Display/lt142_c32 ,open_n2583}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_4  (
    .a(\u2_Display/n4516 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c4 ),
    .o({\u2_Display/lt142_c5 ,open_n2584}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_5  (
    .a(\u2_Display/n4515 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c5 ),
    .o({\u2_Display/lt142_c6 ,open_n2585}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_6  (
    .a(\u2_Display/n4514 ),
    .b(1'b1),
    .c(\u2_Display/lt142_c6 ),
    .o({\u2_Display/lt142_c7 ,open_n2586}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_7  (
    .a(\u2_Display/n4513 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c7 ),
    .o({\u2_Display/lt142_c8 ,open_n2587}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_8  (
    .a(\u2_Display/n4512 ),
    .b(1'b0),
    .c(\u2_Display/lt142_c8 ),
    .o({\u2_Display/lt142_c9 ,open_n2588}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_9  (
    .a(\u2_Display/n4511 ),
    .b(1'b1),
    .c(\u2_Display/lt142_c9 ),
    .o({\u2_Display/lt142_c10 ,open_n2589}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt142_cin  (
    .a(1'b0),
    .o({\u2_Display/lt142_c0 ,open_n2592}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt142_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt142_c32 ),
    .o({open_n2593,\u2_Display/n4521 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_0  (
    .a(\u2_Display/n4555 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c0 ),
    .o({\u2_Display/lt143_c1 ,open_n2594}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_1  (
    .a(\u2_Display/n4554 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c1 ),
    .o({\u2_Display/lt143_c2 ,open_n2595}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_10  (
    .a(\u2_Display/n4545 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c10 ),
    .o({\u2_Display/lt143_c11 ,open_n2596}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_11  (
    .a(\u2_Display/n4544 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c11 ),
    .o({\u2_Display/lt143_c12 ,open_n2597}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_12  (
    .a(\u2_Display/n4543 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c12 ),
    .o({\u2_Display/lt143_c13 ,open_n2598}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_13  (
    .a(\u2_Display/n4542 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c13 ),
    .o({\u2_Display/lt143_c14 ,open_n2599}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_14  (
    .a(\u2_Display/n4541 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c14 ),
    .o({\u2_Display/lt143_c15 ,open_n2600}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_15  (
    .a(\u2_Display/n4540 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c15 ),
    .o({\u2_Display/lt143_c16 ,open_n2601}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_16  (
    .a(\u2_Display/n4539 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c16 ),
    .o({\u2_Display/lt143_c17 ,open_n2602}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_17  (
    .a(\u2_Display/n4538 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c17 ),
    .o({\u2_Display/lt143_c18 ,open_n2603}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_18  (
    .a(\u2_Display/n4537 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c18 ),
    .o({\u2_Display/lt143_c19 ,open_n2604}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_19  (
    .a(\u2_Display/n4536 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c19 ),
    .o({\u2_Display/lt143_c20 ,open_n2605}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_2  (
    .a(\u2_Display/n4553 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c2 ),
    .o({\u2_Display/lt143_c3 ,open_n2606}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_20  (
    .a(\u2_Display/n4535 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c20 ),
    .o({\u2_Display/lt143_c21 ,open_n2607}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_21  (
    .a(\u2_Display/n4534 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c21 ),
    .o({\u2_Display/lt143_c22 ,open_n2608}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_22  (
    .a(\u2_Display/n4533 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c22 ),
    .o({\u2_Display/lt143_c23 ,open_n2609}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_23  (
    .a(\u2_Display/n4532 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c23 ),
    .o({\u2_Display/lt143_c24 ,open_n2610}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_24  (
    .a(\u2_Display/n4531 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c24 ),
    .o({\u2_Display/lt143_c25 ,open_n2611}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_25  (
    .a(\u2_Display/n4530 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c25 ),
    .o({\u2_Display/lt143_c26 ,open_n2612}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_26  (
    .a(\u2_Display/n4529 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c26 ),
    .o({\u2_Display/lt143_c27 ,open_n2613}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_27  (
    .a(\u2_Display/n4528 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c27 ),
    .o({\u2_Display/lt143_c28 ,open_n2614}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_28  (
    .a(\u2_Display/n4527 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c28 ),
    .o({\u2_Display/lt143_c29 ,open_n2615}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_29  (
    .a(\u2_Display/n4526 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c29 ),
    .o({\u2_Display/lt143_c30 ,open_n2616}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_3  (
    .a(\u2_Display/n4552 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c3 ),
    .o({\u2_Display/lt143_c4 ,open_n2617}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_30  (
    .a(\u2_Display/n4525 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c30 ),
    .o({\u2_Display/lt143_c31 ,open_n2618}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_31  (
    .a(\u2_Display/n4524 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c31 ),
    .o({\u2_Display/lt143_c32 ,open_n2619}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_4  (
    .a(\u2_Display/n4551 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c4 ),
    .o({\u2_Display/lt143_c5 ,open_n2620}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_5  (
    .a(\u2_Display/n4550 ),
    .b(1'b1),
    .c(\u2_Display/lt143_c5 ),
    .o({\u2_Display/lt143_c6 ,open_n2621}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_6  (
    .a(\u2_Display/n4549 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c6 ),
    .o({\u2_Display/lt143_c7 ,open_n2622}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_7  (
    .a(\u2_Display/n4548 ),
    .b(1'b0),
    .c(\u2_Display/lt143_c7 ),
    .o({\u2_Display/lt143_c8 ,open_n2623}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_8  (
    .a(\u2_Display/n4547 ),
    .b(1'b1),
    .c(\u2_Display/lt143_c8 ),
    .o({\u2_Display/lt143_c9 ,open_n2624}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_9  (
    .a(\u2_Display/n4546 ),
    .b(1'b1),
    .c(\u2_Display/lt143_c9 ),
    .o({\u2_Display/lt143_c10 ,open_n2625}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt143_cin  (
    .a(1'b0),
    .o({\u2_Display/lt143_c0 ,open_n2628}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt143_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt143_c32 ),
    .o({open_n2629,\u2_Display/n4556 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_0  (
    .a(\u2_Display/counta [0]),
    .b(1'b0),
    .c(\u2_Display/lt154_c0 ),
    .o({\u2_Display/lt154_c1 ,open_n2630}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_1  (
    .a(\u2_Display/counta [1]),
    .b(1'b0),
    .c(\u2_Display/lt154_c1 ),
    .o({\u2_Display/lt154_c2 ,open_n2631}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_10  (
    .a(\u2_Display/counta [10]),
    .b(1'b0),
    .c(\u2_Display/lt154_c10 ),
    .o({\u2_Display/lt154_c11 ,open_n2632}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_11  (
    .a(\u2_Display/counta [11]),
    .b(1'b0),
    .c(\u2_Display/lt154_c11 ),
    .o({\u2_Display/lt154_c12 ,open_n2633}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_12  (
    .a(\u2_Display/counta [12]),
    .b(1'b0),
    .c(\u2_Display/lt154_c12 ),
    .o({\u2_Display/lt154_c13 ,open_n2634}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_13  (
    .a(\u2_Display/counta [13]),
    .b(1'b0),
    .c(\u2_Display/lt154_c13 ),
    .o({\u2_Display/lt154_c14 ,open_n2635}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_14  (
    .a(\u2_Display/counta [14]),
    .b(1'b0),
    .c(\u2_Display/lt154_c14 ),
    .o({\u2_Display/lt154_c15 ,open_n2636}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_15  (
    .a(\u2_Display/counta [15]),
    .b(1'b0),
    .c(\u2_Display/lt154_c15 ),
    .o({\u2_Display/lt154_c16 ,open_n2637}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_16  (
    .a(\u2_Display/counta [16]),
    .b(1'b0),
    .c(\u2_Display/lt154_c16 ),
    .o({\u2_Display/lt154_c17 ,open_n2638}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_17  (
    .a(\u2_Display/counta [17]),
    .b(1'b0),
    .c(\u2_Display/lt154_c17 ),
    .o({\u2_Display/lt154_c18 ,open_n2639}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_18  (
    .a(\u2_Display/counta [18]),
    .b(1'b0),
    .c(\u2_Display/lt154_c18 ),
    .o({\u2_Display/lt154_c19 ,open_n2640}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_19  (
    .a(\u2_Display/counta [19]),
    .b(1'b0),
    .c(\u2_Display/lt154_c19 ),
    .o({\u2_Display/lt154_c20 ,open_n2641}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_2  (
    .a(\u2_Display/counta [2]),
    .b(1'b0),
    .c(\u2_Display/lt154_c2 ),
    .o({\u2_Display/lt154_c3 ,open_n2642}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_20  (
    .a(\u2_Display/counta [20]),
    .b(1'b0),
    .c(\u2_Display/lt154_c20 ),
    .o({\u2_Display/lt154_c21 ,open_n2643}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_21  (
    .a(\u2_Display/counta [21]),
    .b(1'b0),
    .c(\u2_Display/lt154_c21 ),
    .o({\u2_Display/lt154_c22 ,open_n2644}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_22  (
    .a(\u2_Display/counta [22]),
    .b(1'b0),
    .c(\u2_Display/lt154_c22 ),
    .o({\u2_Display/lt154_c23 ,open_n2645}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_23  (
    .a(\u2_Display/counta [23]),
    .b(1'b0),
    .c(\u2_Display/lt154_c23 ),
    .o({\u2_Display/lt154_c24 ,open_n2646}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_24  (
    .a(\u2_Display/counta [24]),
    .b(1'b0),
    .c(\u2_Display/lt154_c24 ),
    .o({\u2_Display/lt154_c25 ,open_n2647}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_25  (
    .a(\u2_Display/counta [25]),
    .b(1'b0),
    .c(\u2_Display/lt154_c25 ),
    .o({\u2_Display/lt154_c26 ,open_n2648}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_26  (
    .a(\u2_Display/counta [26]),
    .b(1'b0),
    .c(\u2_Display/lt154_c26 ),
    .o({\u2_Display/lt154_c27 ,open_n2649}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_27  (
    .a(\u2_Display/counta [27]),
    .b(1'b0),
    .c(\u2_Display/lt154_c27 ),
    .o({\u2_Display/lt154_c28 ,open_n2650}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_28  (
    .a(\u2_Display/counta [28]),
    .b(1'b0),
    .c(\u2_Display/lt154_c28 ),
    .o({\u2_Display/lt154_c29 ,open_n2651}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_29  (
    .a(\u2_Display/counta [29]),
    .b(1'b1),
    .c(\u2_Display/lt154_c29 ),
    .o({\u2_Display/lt154_c30 ,open_n2652}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_3  (
    .a(\u2_Display/counta [3]),
    .b(1'b0),
    .c(\u2_Display/lt154_c3 ),
    .o({\u2_Display/lt154_c4 ,open_n2653}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_30  (
    .a(\u2_Display/counta [30]),
    .b(1'b0),
    .c(\u2_Display/lt154_c30 ),
    .o({\u2_Display/lt154_c31 ,open_n2654}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_31  (
    .a(\u2_Display/counta [31]),
    .b(1'b1),
    .c(\u2_Display/lt154_c31 ),
    .o({\u2_Display/lt154_c32 ,open_n2655}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_4  (
    .a(\u2_Display/counta [4]),
    .b(1'b0),
    .c(\u2_Display/lt154_c4 ),
    .o({\u2_Display/lt154_c5 ,open_n2656}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_5  (
    .a(\u2_Display/counta [5]),
    .b(1'b0),
    .c(\u2_Display/lt154_c5 ),
    .o({\u2_Display/lt154_c6 ,open_n2657}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_6  (
    .a(\u2_Display/counta [6]),
    .b(1'b0),
    .c(\u2_Display/lt154_c6 ),
    .o({\u2_Display/lt154_c7 ,open_n2658}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_7  (
    .a(\u2_Display/counta [7]),
    .b(1'b0),
    .c(\u2_Display/lt154_c7 ),
    .o({\u2_Display/lt154_c8 ,open_n2659}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_8  (
    .a(\u2_Display/counta [8]),
    .b(1'b0),
    .c(\u2_Display/lt154_c8 ),
    .o({\u2_Display/lt154_c9 ,open_n2660}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_9  (
    .a(\u2_Display/counta [9]),
    .b(1'b0),
    .c(\u2_Display/lt154_c9 ),
    .o({\u2_Display/lt154_c10 ,open_n2661}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt154_cin  (
    .a(1'b0),
    .o({\u2_Display/lt154_c0 ,open_n2664}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt154_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt154_c32 ),
    .o({open_n2665,\u2_Display/n4909 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_0  (
    .a(\u2_Display/n6101 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c0 ),
    .o({\u2_Display/lt155_c1 ,open_n2666}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_1  (
    .a(\u2_Display/n6100 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c1 ),
    .o({\u2_Display/lt155_c2 ,open_n2667}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_10  (
    .a(\u2_Display/n6091 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c10 ),
    .o({\u2_Display/lt155_c11 ,open_n2668}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_11  (
    .a(\u2_Display/n6090 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c11 ),
    .o({\u2_Display/lt155_c12 ,open_n2669}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_12  (
    .a(\u2_Display/n6089 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c12 ),
    .o({\u2_Display/lt155_c13 ,open_n2670}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_13  (
    .a(\u2_Display/n6088 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c13 ),
    .o({\u2_Display/lt155_c14 ,open_n2671}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_14  (
    .a(\u2_Display/n6087 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c14 ),
    .o({\u2_Display/lt155_c15 ,open_n2672}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_15  (
    .a(\u2_Display/n6086 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c15 ),
    .o({\u2_Display/lt155_c16 ,open_n2673}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_16  (
    .a(\u2_Display/n6085 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c16 ),
    .o({\u2_Display/lt155_c17 ,open_n2674}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_17  (
    .a(\u2_Display/n6084 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c17 ),
    .o({\u2_Display/lt155_c18 ,open_n2675}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_18  (
    .a(\u2_Display/n6083 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c18 ),
    .o({\u2_Display/lt155_c19 ,open_n2676}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_19  (
    .a(\u2_Display/n6082 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c19 ),
    .o({\u2_Display/lt155_c20 ,open_n2677}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_2  (
    .a(\u2_Display/n6099 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c2 ),
    .o({\u2_Display/lt155_c3 ,open_n2678}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_20  (
    .a(\u2_Display/n6081 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c20 ),
    .o({\u2_Display/lt155_c21 ,open_n2679}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_21  (
    .a(\u2_Display/n6080 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c21 ),
    .o({\u2_Display/lt155_c22 ,open_n2680}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_22  (
    .a(\u2_Display/n6079 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c22 ),
    .o({\u2_Display/lt155_c23 ,open_n2681}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_23  (
    .a(\u2_Display/n6078 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c23 ),
    .o({\u2_Display/lt155_c24 ,open_n2682}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_24  (
    .a(\u2_Display/n6077 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c24 ),
    .o({\u2_Display/lt155_c25 ,open_n2683}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_25  (
    .a(\u2_Display/n6076 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c25 ),
    .o({\u2_Display/lt155_c26 ,open_n2684}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_26  (
    .a(\u2_Display/n6075 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c26 ),
    .o({\u2_Display/lt155_c27 ,open_n2685}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_27  (
    .a(\u2_Display/n6074 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c27 ),
    .o({\u2_Display/lt155_c28 ,open_n2686}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_28  (
    .a(\u2_Display/n6073 ),
    .b(1'b1),
    .c(\u2_Display/lt155_c28 ),
    .o({\u2_Display/lt155_c29 ,open_n2687}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_29  (
    .a(\u2_Display/n6072 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c29 ),
    .o({\u2_Display/lt155_c30 ,open_n2688}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_3  (
    .a(\u2_Display/n6098 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c3 ),
    .o({\u2_Display/lt155_c4 ,open_n2689}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_30  (
    .a(\u2_Display/n6071 ),
    .b(1'b1),
    .c(\u2_Display/lt155_c30 ),
    .o({\u2_Display/lt155_c31 ,open_n2690}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_31  (
    .a(\u2_Display/n6070 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c31 ),
    .o({\u2_Display/lt155_c32 ,open_n2691}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_4  (
    .a(\u2_Display/n6097 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c4 ),
    .o({\u2_Display/lt155_c5 ,open_n2692}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_5  (
    .a(\u2_Display/n6096 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c5 ),
    .o({\u2_Display/lt155_c6 ,open_n2693}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_6  (
    .a(\u2_Display/n6095 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c6 ),
    .o({\u2_Display/lt155_c7 ,open_n2694}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_7  (
    .a(\u2_Display/n6094 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c7 ),
    .o({\u2_Display/lt155_c8 ,open_n2695}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_8  (
    .a(\u2_Display/n6093 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c8 ),
    .o({\u2_Display/lt155_c9 ,open_n2696}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_9  (
    .a(\u2_Display/n6092 ),
    .b(1'b0),
    .c(\u2_Display/lt155_c9 ),
    .o({\u2_Display/lt155_c10 ,open_n2697}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt155_cin  (
    .a(1'b0),
    .o({\u2_Display/lt155_c0 ,open_n2700}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt155_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt155_c32 ),
    .o({open_n2701,\u2_Display/n4944 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_0  (
    .a(\u2_Display/n6136 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c0 ),
    .o({\u2_Display/lt156_c1 ,open_n2702}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_1  (
    .a(\u2_Display/n6135 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c1 ),
    .o({\u2_Display/lt156_c2 ,open_n2703}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_10  (
    .a(\u2_Display/n6126 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c10 ),
    .o({\u2_Display/lt156_c11 ,open_n2704}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_11  (
    .a(\u2_Display/n6125 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c11 ),
    .o({\u2_Display/lt156_c12 ,open_n2705}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_12  (
    .a(\u2_Display/n6124 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c12 ),
    .o({\u2_Display/lt156_c13 ,open_n2706}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_13  (
    .a(\u2_Display/n6123 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c13 ),
    .o({\u2_Display/lt156_c14 ,open_n2707}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_14  (
    .a(\u2_Display/n6122 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c14 ),
    .o({\u2_Display/lt156_c15 ,open_n2708}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_15  (
    .a(\u2_Display/n6121 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c15 ),
    .o({\u2_Display/lt156_c16 ,open_n2709}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_16  (
    .a(\u2_Display/n6120 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c16 ),
    .o({\u2_Display/lt156_c17 ,open_n2710}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_17  (
    .a(\u2_Display/n6119 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c17 ),
    .o({\u2_Display/lt156_c18 ,open_n2711}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_18  (
    .a(\u2_Display/n6118 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c18 ),
    .o({\u2_Display/lt156_c19 ,open_n2712}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_19  (
    .a(\u2_Display/n6117 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c19 ),
    .o({\u2_Display/lt156_c20 ,open_n2713}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_2  (
    .a(\u2_Display/n6134 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c2 ),
    .o({\u2_Display/lt156_c3 ,open_n2714}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_20  (
    .a(\u2_Display/n6116 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c20 ),
    .o({\u2_Display/lt156_c21 ,open_n2715}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_21  (
    .a(\u2_Display/n6115 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c21 ),
    .o({\u2_Display/lt156_c22 ,open_n2716}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_22  (
    .a(\u2_Display/n6114 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c22 ),
    .o({\u2_Display/lt156_c23 ,open_n2717}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_23  (
    .a(\u2_Display/n6113 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c23 ),
    .o({\u2_Display/lt156_c24 ,open_n2718}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_24  (
    .a(\u2_Display/n6112 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c24 ),
    .o({\u2_Display/lt156_c25 ,open_n2719}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_25  (
    .a(\u2_Display/n6111 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c25 ),
    .o({\u2_Display/lt156_c26 ,open_n2720}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_26  (
    .a(\u2_Display/n6110 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c26 ),
    .o({\u2_Display/lt156_c27 ,open_n2721}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_27  (
    .a(\u2_Display/n6109 ),
    .b(1'b1),
    .c(\u2_Display/lt156_c27 ),
    .o({\u2_Display/lt156_c28 ,open_n2722}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_28  (
    .a(\u2_Display/n6108 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c28 ),
    .o({\u2_Display/lt156_c29 ,open_n2723}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_29  (
    .a(\u2_Display/n6107 ),
    .b(1'b1),
    .c(\u2_Display/lt156_c29 ),
    .o({\u2_Display/lt156_c30 ,open_n2724}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_3  (
    .a(\u2_Display/n6133 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c3 ),
    .o({\u2_Display/lt156_c4 ,open_n2725}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_30  (
    .a(\u2_Display/n6106 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c30 ),
    .o({\u2_Display/lt156_c31 ,open_n2726}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_31  (
    .a(\u2_Display/n6105 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c31 ),
    .o({\u2_Display/lt156_c32 ,open_n2727}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_4  (
    .a(\u2_Display/n6132 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c4 ),
    .o({\u2_Display/lt156_c5 ,open_n2728}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_5  (
    .a(\u2_Display/n6131 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c5 ),
    .o({\u2_Display/lt156_c6 ,open_n2729}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_6  (
    .a(\u2_Display/n6130 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c6 ),
    .o({\u2_Display/lt156_c7 ,open_n2730}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_7  (
    .a(\u2_Display/n6129 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c7 ),
    .o({\u2_Display/lt156_c8 ,open_n2731}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_8  (
    .a(\u2_Display/n6128 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c8 ),
    .o({\u2_Display/lt156_c9 ,open_n2732}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_9  (
    .a(\u2_Display/n6127 ),
    .b(1'b0),
    .c(\u2_Display/lt156_c9 ),
    .o({\u2_Display/lt156_c10 ,open_n2733}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt156_cin  (
    .a(1'b0),
    .o({\u2_Display/lt156_c0 ,open_n2736}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt156_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt156_c32 ),
    .o({open_n2737,\u2_Display/n4979 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_0  (
    .a(\u2_Display/n6171 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c0 ),
    .o({\u2_Display/lt157_c1 ,open_n2738}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_1  (
    .a(\u2_Display/n6170 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c1 ),
    .o({\u2_Display/lt157_c2 ,open_n2739}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_10  (
    .a(\u2_Display/n6161 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c10 ),
    .o({\u2_Display/lt157_c11 ,open_n2740}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_11  (
    .a(\u2_Display/n6160 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c11 ),
    .o({\u2_Display/lt157_c12 ,open_n2741}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_12  (
    .a(\u2_Display/n6159 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c12 ),
    .o({\u2_Display/lt157_c13 ,open_n2742}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_13  (
    .a(\u2_Display/n6158 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c13 ),
    .o({\u2_Display/lt157_c14 ,open_n2743}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_14  (
    .a(\u2_Display/n6157 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c14 ),
    .o({\u2_Display/lt157_c15 ,open_n2744}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_15  (
    .a(\u2_Display/n6156 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c15 ),
    .o({\u2_Display/lt157_c16 ,open_n2745}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_16  (
    .a(\u2_Display/n6155 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c16 ),
    .o({\u2_Display/lt157_c17 ,open_n2746}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_17  (
    .a(\u2_Display/n6154 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c17 ),
    .o({\u2_Display/lt157_c18 ,open_n2747}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_18  (
    .a(\u2_Display/n6153 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c18 ),
    .o({\u2_Display/lt157_c19 ,open_n2748}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_19  (
    .a(\u2_Display/n6152 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c19 ),
    .o({\u2_Display/lt157_c20 ,open_n2749}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_2  (
    .a(\u2_Display/n6169 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c2 ),
    .o({\u2_Display/lt157_c3 ,open_n2750}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_20  (
    .a(\u2_Display/n6151 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c20 ),
    .o({\u2_Display/lt157_c21 ,open_n2751}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_21  (
    .a(\u2_Display/n6150 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c21 ),
    .o({\u2_Display/lt157_c22 ,open_n2752}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_22  (
    .a(\u2_Display/n6149 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c22 ),
    .o({\u2_Display/lt157_c23 ,open_n2753}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_23  (
    .a(\u2_Display/n6148 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c23 ),
    .o({\u2_Display/lt157_c24 ,open_n2754}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_24  (
    .a(\u2_Display/n6147 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c24 ),
    .o({\u2_Display/lt157_c25 ,open_n2755}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_25  (
    .a(\u2_Display/n6146 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c25 ),
    .o({\u2_Display/lt157_c26 ,open_n2756}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_26  (
    .a(\u2_Display/n6145 ),
    .b(1'b1),
    .c(\u2_Display/lt157_c26 ),
    .o({\u2_Display/lt157_c27 ,open_n2757}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_27  (
    .a(\u2_Display/n6144 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c27 ),
    .o({\u2_Display/lt157_c28 ,open_n2758}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_28  (
    .a(\u2_Display/n6143 ),
    .b(1'b1),
    .c(\u2_Display/lt157_c28 ),
    .o({\u2_Display/lt157_c29 ,open_n2759}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_29  (
    .a(\u2_Display/n6142 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c29 ),
    .o({\u2_Display/lt157_c30 ,open_n2760}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_3  (
    .a(\u2_Display/n6168 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c3 ),
    .o({\u2_Display/lt157_c4 ,open_n2761}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_30  (
    .a(\u2_Display/n6141 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c30 ),
    .o({\u2_Display/lt157_c31 ,open_n2762}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_31  (
    .a(\u2_Display/n6140 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c31 ),
    .o({\u2_Display/lt157_c32 ,open_n2763}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_4  (
    .a(\u2_Display/n6167 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c4 ),
    .o({\u2_Display/lt157_c5 ,open_n2764}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_5  (
    .a(\u2_Display/n6166 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c5 ),
    .o({\u2_Display/lt157_c6 ,open_n2765}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_6  (
    .a(\u2_Display/n6165 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c6 ),
    .o({\u2_Display/lt157_c7 ,open_n2766}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_7  (
    .a(\u2_Display/n6164 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c7 ),
    .o({\u2_Display/lt157_c8 ,open_n2767}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_8  (
    .a(\u2_Display/n6163 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c8 ),
    .o({\u2_Display/lt157_c9 ,open_n2768}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_9  (
    .a(\u2_Display/n6162 ),
    .b(1'b0),
    .c(\u2_Display/lt157_c9 ),
    .o({\u2_Display/lt157_c10 ,open_n2769}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt157_cin  (
    .a(1'b0),
    .o({\u2_Display/lt157_c0 ,open_n2772}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt157_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt157_c32 ),
    .o({open_n2773,\u2_Display/n5014 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_0  (
    .a(\u2_Display/n6206 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c0 ),
    .o({\u2_Display/lt158_c1 ,open_n2774}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_1  (
    .a(\u2_Display/n6205 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c1 ),
    .o({\u2_Display/lt158_c2 ,open_n2775}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_10  (
    .a(\u2_Display/n6196 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c10 ),
    .o({\u2_Display/lt158_c11 ,open_n2776}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_11  (
    .a(\u2_Display/n6195 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c11 ),
    .o({\u2_Display/lt158_c12 ,open_n2777}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_12  (
    .a(\u2_Display/n6194 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c12 ),
    .o({\u2_Display/lt158_c13 ,open_n2778}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_13  (
    .a(\u2_Display/n6193 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c13 ),
    .o({\u2_Display/lt158_c14 ,open_n2779}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_14  (
    .a(\u2_Display/n6192 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c14 ),
    .o({\u2_Display/lt158_c15 ,open_n2780}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_15  (
    .a(\u2_Display/n6191 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c15 ),
    .o({\u2_Display/lt158_c16 ,open_n2781}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_16  (
    .a(\u2_Display/n6190 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c16 ),
    .o({\u2_Display/lt158_c17 ,open_n2782}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_17  (
    .a(\u2_Display/n6189 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c17 ),
    .o({\u2_Display/lt158_c18 ,open_n2783}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_18  (
    .a(\u2_Display/n6188 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c18 ),
    .o({\u2_Display/lt158_c19 ,open_n2784}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_19  (
    .a(\u2_Display/n6187 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c19 ),
    .o({\u2_Display/lt158_c20 ,open_n2785}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_2  (
    .a(\u2_Display/n6204 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c2 ),
    .o({\u2_Display/lt158_c3 ,open_n2786}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_20  (
    .a(\u2_Display/n6186 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c20 ),
    .o({\u2_Display/lt158_c21 ,open_n2787}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_21  (
    .a(\u2_Display/n6185 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c21 ),
    .o({\u2_Display/lt158_c22 ,open_n2788}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_22  (
    .a(\u2_Display/n6184 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c22 ),
    .o({\u2_Display/lt158_c23 ,open_n2789}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_23  (
    .a(\u2_Display/n6183 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c23 ),
    .o({\u2_Display/lt158_c24 ,open_n2790}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_24  (
    .a(\u2_Display/n6182 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c24 ),
    .o({\u2_Display/lt158_c25 ,open_n2791}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_25  (
    .a(\u2_Display/n6181 ),
    .b(1'b1),
    .c(\u2_Display/lt158_c25 ),
    .o({\u2_Display/lt158_c26 ,open_n2792}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_26  (
    .a(\u2_Display/n6180 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c26 ),
    .o({\u2_Display/lt158_c27 ,open_n2793}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_27  (
    .a(\u2_Display/n6179 ),
    .b(1'b1),
    .c(\u2_Display/lt158_c27 ),
    .o({\u2_Display/lt158_c28 ,open_n2794}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_28  (
    .a(\u2_Display/n6178 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c28 ),
    .o({\u2_Display/lt158_c29 ,open_n2795}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_29  (
    .a(\u2_Display/n6177 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c29 ),
    .o({\u2_Display/lt158_c30 ,open_n2796}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_3  (
    .a(\u2_Display/n6203 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c3 ),
    .o({\u2_Display/lt158_c4 ,open_n2797}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_30  (
    .a(\u2_Display/n6176 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c30 ),
    .o({\u2_Display/lt158_c31 ,open_n2798}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_31  (
    .a(\u2_Display/n6175 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c31 ),
    .o({\u2_Display/lt158_c32 ,open_n2799}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_4  (
    .a(\u2_Display/n6202 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c4 ),
    .o({\u2_Display/lt158_c5 ,open_n2800}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_5  (
    .a(\u2_Display/n6201 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c5 ),
    .o({\u2_Display/lt158_c6 ,open_n2801}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_6  (
    .a(\u2_Display/n6200 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c6 ),
    .o({\u2_Display/lt158_c7 ,open_n2802}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_7  (
    .a(\u2_Display/n6199 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c7 ),
    .o({\u2_Display/lt158_c8 ,open_n2803}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_8  (
    .a(\u2_Display/n6198 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c8 ),
    .o({\u2_Display/lt158_c9 ,open_n2804}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_9  (
    .a(\u2_Display/n6197 ),
    .b(1'b0),
    .c(\u2_Display/lt158_c9 ),
    .o({\u2_Display/lt158_c10 ,open_n2805}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt158_cin  (
    .a(1'b0),
    .o({\u2_Display/lt158_c0 ,open_n2808}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt158_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt158_c32 ),
    .o({open_n2809,\u2_Display/n5049 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_0  (
    .a(\u2_Display/n6241 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c0 ),
    .o({\u2_Display/lt159_c1 ,open_n2810}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_1  (
    .a(\u2_Display/n6240 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c1 ),
    .o({\u2_Display/lt159_c2 ,open_n2811}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_10  (
    .a(\u2_Display/n6231 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c10 ),
    .o({\u2_Display/lt159_c11 ,open_n2812}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_11  (
    .a(\u2_Display/n6230 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c11 ),
    .o({\u2_Display/lt159_c12 ,open_n2813}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_12  (
    .a(\u2_Display/n6229 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c12 ),
    .o({\u2_Display/lt159_c13 ,open_n2814}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_13  (
    .a(\u2_Display/n6228 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c13 ),
    .o({\u2_Display/lt159_c14 ,open_n2815}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_14  (
    .a(\u2_Display/n6227 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c14 ),
    .o({\u2_Display/lt159_c15 ,open_n2816}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_15  (
    .a(\u2_Display/n6226 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c15 ),
    .o({\u2_Display/lt159_c16 ,open_n2817}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_16  (
    .a(\u2_Display/n6225 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c16 ),
    .o({\u2_Display/lt159_c17 ,open_n2818}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_17  (
    .a(\u2_Display/n6224 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c17 ),
    .o({\u2_Display/lt159_c18 ,open_n2819}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_18  (
    .a(\u2_Display/n6223 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c18 ),
    .o({\u2_Display/lt159_c19 ,open_n2820}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_19  (
    .a(\u2_Display/n6222 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c19 ),
    .o({\u2_Display/lt159_c20 ,open_n2821}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_2  (
    .a(\u2_Display/n6239 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c2 ),
    .o({\u2_Display/lt159_c3 ,open_n2822}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_20  (
    .a(\u2_Display/n6221 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c20 ),
    .o({\u2_Display/lt159_c21 ,open_n2823}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_21  (
    .a(\u2_Display/n6220 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c21 ),
    .o({\u2_Display/lt159_c22 ,open_n2824}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_22  (
    .a(\u2_Display/n6219 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c22 ),
    .o({\u2_Display/lt159_c23 ,open_n2825}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_23  (
    .a(\u2_Display/n6218 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c23 ),
    .o({\u2_Display/lt159_c24 ,open_n2826}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_24  (
    .a(\u2_Display/n6217 ),
    .b(1'b1),
    .c(\u2_Display/lt159_c24 ),
    .o({\u2_Display/lt159_c25 ,open_n2827}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_25  (
    .a(\u2_Display/n6216 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c25 ),
    .o({\u2_Display/lt159_c26 ,open_n2828}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_26  (
    .a(\u2_Display/n6215 ),
    .b(1'b1),
    .c(\u2_Display/lt159_c26 ),
    .o({\u2_Display/lt159_c27 ,open_n2829}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_27  (
    .a(\u2_Display/n6214 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c27 ),
    .o({\u2_Display/lt159_c28 ,open_n2830}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_28  (
    .a(\u2_Display/n6213 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c28 ),
    .o({\u2_Display/lt159_c29 ,open_n2831}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_29  (
    .a(\u2_Display/n6212 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c29 ),
    .o({\u2_Display/lt159_c30 ,open_n2832}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_3  (
    .a(\u2_Display/n6238 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c3 ),
    .o({\u2_Display/lt159_c4 ,open_n2833}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_30  (
    .a(\u2_Display/n6211 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c30 ),
    .o({\u2_Display/lt159_c31 ,open_n2834}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_31  (
    .a(\u2_Display/n6210 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c31 ),
    .o({\u2_Display/lt159_c32 ,open_n2835}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_4  (
    .a(\u2_Display/n6237 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c4 ),
    .o({\u2_Display/lt159_c5 ,open_n2836}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_5  (
    .a(\u2_Display/n6236 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c5 ),
    .o({\u2_Display/lt159_c6 ,open_n2837}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_6  (
    .a(\u2_Display/n6235 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c6 ),
    .o({\u2_Display/lt159_c7 ,open_n2838}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_7  (
    .a(\u2_Display/n6234 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c7 ),
    .o({\u2_Display/lt159_c8 ,open_n2839}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_8  (
    .a(\u2_Display/n6233 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c8 ),
    .o({\u2_Display/lt159_c9 ,open_n2840}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_9  (
    .a(\u2_Display/n6232 ),
    .b(1'b0),
    .c(\u2_Display/lt159_c9 ),
    .o({\u2_Display/lt159_c10 ,open_n2841}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt159_cin  (
    .a(1'b0),
    .o({\u2_Display/lt159_c0 ,open_n2844}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt159_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt159_c32 ),
    .o({open_n2845,\u2_Display/n5084 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_0  (
    .a(\u2_Display/n6276 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c0 ),
    .o({\u2_Display/lt160_c1 ,open_n2846}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_1  (
    .a(\u2_Display/n6275 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c1 ),
    .o({\u2_Display/lt160_c2 ,open_n2847}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_10  (
    .a(\u2_Display/n6266 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c10 ),
    .o({\u2_Display/lt160_c11 ,open_n2848}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_11  (
    .a(\u2_Display/n6265 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c11 ),
    .o({\u2_Display/lt160_c12 ,open_n2849}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_12  (
    .a(\u2_Display/n6264 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c12 ),
    .o({\u2_Display/lt160_c13 ,open_n2850}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_13  (
    .a(\u2_Display/n6263 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c13 ),
    .o({\u2_Display/lt160_c14 ,open_n2851}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_14  (
    .a(\u2_Display/n6262 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c14 ),
    .o({\u2_Display/lt160_c15 ,open_n2852}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_15  (
    .a(\u2_Display/n6261 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c15 ),
    .o({\u2_Display/lt160_c16 ,open_n2853}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_16  (
    .a(\u2_Display/n6260 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c16 ),
    .o({\u2_Display/lt160_c17 ,open_n2854}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_17  (
    .a(\u2_Display/n6259 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c17 ),
    .o({\u2_Display/lt160_c18 ,open_n2855}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_18  (
    .a(\u2_Display/n6258 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c18 ),
    .o({\u2_Display/lt160_c19 ,open_n2856}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_19  (
    .a(\u2_Display/n6257 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c19 ),
    .o({\u2_Display/lt160_c20 ,open_n2857}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_2  (
    .a(\u2_Display/n6274 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c2 ),
    .o({\u2_Display/lt160_c3 ,open_n2858}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_20  (
    .a(\u2_Display/n6256 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c20 ),
    .o({\u2_Display/lt160_c21 ,open_n2859}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_21  (
    .a(\u2_Display/n6255 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c21 ),
    .o({\u2_Display/lt160_c22 ,open_n2860}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_22  (
    .a(\u2_Display/n6254 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c22 ),
    .o({\u2_Display/lt160_c23 ,open_n2861}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_23  (
    .a(\u2_Display/n6253 ),
    .b(1'b1),
    .c(\u2_Display/lt160_c23 ),
    .o({\u2_Display/lt160_c24 ,open_n2862}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_24  (
    .a(\u2_Display/n6252 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c24 ),
    .o({\u2_Display/lt160_c25 ,open_n2863}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_25  (
    .a(\u2_Display/n6251 ),
    .b(1'b1),
    .c(\u2_Display/lt160_c25 ),
    .o({\u2_Display/lt160_c26 ,open_n2864}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_26  (
    .a(\u2_Display/n6250 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c26 ),
    .o({\u2_Display/lt160_c27 ,open_n2865}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_27  (
    .a(\u2_Display/n6249 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c27 ),
    .o({\u2_Display/lt160_c28 ,open_n2866}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_28  (
    .a(\u2_Display/n6248 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c28 ),
    .o({\u2_Display/lt160_c29 ,open_n2867}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_29  (
    .a(\u2_Display/n6247 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c29 ),
    .o({\u2_Display/lt160_c30 ,open_n2868}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_3  (
    .a(\u2_Display/n6273 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c3 ),
    .o({\u2_Display/lt160_c4 ,open_n2869}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_30  (
    .a(\u2_Display/n6246 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c30 ),
    .o({\u2_Display/lt160_c31 ,open_n2870}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_31  (
    .a(\u2_Display/n6245 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c31 ),
    .o({\u2_Display/lt160_c32 ,open_n2871}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_4  (
    .a(\u2_Display/n6272 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c4 ),
    .o({\u2_Display/lt160_c5 ,open_n2872}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_5  (
    .a(\u2_Display/n6271 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c5 ),
    .o({\u2_Display/lt160_c6 ,open_n2873}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_6  (
    .a(\u2_Display/n6270 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c6 ),
    .o({\u2_Display/lt160_c7 ,open_n2874}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_7  (
    .a(\u2_Display/n6269 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c7 ),
    .o({\u2_Display/lt160_c8 ,open_n2875}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_8  (
    .a(\u2_Display/n6268 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c8 ),
    .o({\u2_Display/lt160_c9 ,open_n2876}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_9  (
    .a(\u2_Display/n6267 ),
    .b(1'b0),
    .c(\u2_Display/lt160_c9 ),
    .o({\u2_Display/lt160_c10 ,open_n2877}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt160_cin  (
    .a(1'b0),
    .o({\u2_Display/lt160_c0 ,open_n2880}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt160_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt160_c32 ),
    .o({open_n2881,\u2_Display/n5119 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_0  (
    .a(\u2_Display/n6311 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c0 ),
    .o({\u2_Display/lt161_c1 ,open_n2882}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_1  (
    .a(\u2_Display/n6310 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c1 ),
    .o({\u2_Display/lt161_c2 ,open_n2883}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_10  (
    .a(\u2_Display/n6301 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c10 ),
    .o({\u2_Display/lt161_c11 ,open_n2884}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_11  (
    .a(\u2_Display/n6300 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c11 ),
    .o({\u2_Display/lt161_c12 ,open_n2885}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_12  (
    .a(\u2_Display/n6299 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c12 ),
    .o({\u2_Display/lt161_c13 ,open_n2886}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_13  (
    .a(\u2_Display/n6298 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c13 ),
    .o({\u2_Display/lt161_c14 ,open_n2887}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_14  (
    .a(\u2_Display/n6297 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c14 ),
    .o({\u2_Display/lt161_c15 ,open_n2888}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_15  (
    .a(\u2_Display/n6296 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c15 ),
    .o({\u2_Display/lt161_c16 ,open_n2889}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_16  (
    .a(\u2_Display/n6295 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c16 ),
    .o({\u2_Display/lt161_c17 ,open_n2890}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_17  (
    .a(\u2_Display/n6294 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c17 ),
    .o({\u2_Display/lt161_c18 ,open_n2891}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_18  (
    .a(\u2_Display/n6293 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c18 ),
    .o({\u2_Display/lt161_c19 ,open_n2892}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_19  (
    .a(\u2_Display/n6292 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c19 ),
    .o({\u2_Display/lt161_c20 ,open_n2893}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_2  (
    .a(\u2_Display/n6309 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c2 ),
    .o({\u2_Display/lt161_c3 ,open_n2894}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_20  (
    .a(\u2_Display/n6291 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c20 ),
    .o({\u2_Display/lt161_c21 ,open_n2895}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_21  (
    .a(\u2_Display/n6290 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c21 ),
    .o({\u2_Display/lt161_c22 ,open_n2896}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_22  (
    .a(\u2_Display/n6289 ),
    .b(1'b1),
    .c(\u2_Display/lt161_c22 ),
    .o({\u2_Display/lt161_c23 ,open_n2897}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_23  (
    .a(\u2_Display/n6288 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c23 ),
    .o({\u2_Display/lt161_c24 ,open_n2898}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_24  (
    .a(\u2_Display/n6287 ),
    .b(1'b1),
    .c(\u2_Display/lt161_c24 ),
    .o({\u2_Display/lt161_c25 ,open_n2899}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_25  (
    .a(\u2_Display/n6286 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c25 ),
    .o({\u2_Display/lt161_c26 ,open_n2900}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_26  (
    .a(\u2_Display/n6285 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c26 ),
    .o({\u2_Display/lt161_c27 ,open_n2901}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_27  (
    .a(\u2_Display/n6284 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c27 ),
    .o({\u2_Display/lt161_c28 ,open_n2902}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_28  (
    .a(\u2_Display/n6283 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c28 ),
    .o({\u2_Display/lt161_c29 ,open_n2903}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_29  (
    .a(\u2_Display/n6282 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c29 ),
    .o({\u2_Display/lt161_c30 ,open_n2904}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_3  (
    .a(\u2_Display/n6308 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c3 ),
    .o({\u2_Display/lt161_c4 ,open_n2905}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_30  (
    .a(\u2_Display/n6281 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c30 ),
    .o({\u2_Display/lt161_c31 ,open_n2906}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_31  (
    .a(\u2_Display/n6280 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c31 ),
    .o({\u2_Display/lt161_c32 ,open_n2907}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_4  (
    .a(\u2_Display/n6307 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c4 ),
    .o({\u2_Display/lt161_c5 ,open_n2908}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_5  (
    .a(\u2_Display/n6306 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c5 ),
    .o({\u2_Display/lt161_c6 ,open_n2909}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_6  (
    .a(\u2_Display/n6305 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c6 ),
    .o({\u2_Display/lt161_c7 ,open_n2910}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_7  (
    .a(\u2_Display/n6304 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c7 ),
    .o({\u2_Display/lt161_c8 ,open_n2911}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_8  (
    .a(\u2_Display/n6303 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c8 ),
    .o({\u2_Display/lt161_c9 ,open_n2912}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_9  (
    .a(\u2_Display/n6302 ),
    .b(1'b0),
    .c(\u2_Display/lt161_c9 ),
    .o({\u2_Display/lt161_c10 ,open_n2913}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt161_cin  (
    .a(1'b0),
    .o({\u2_Display/lt161_c0 ,open_n2916}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt161_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt161_c32 ),
    .o({open_n2917,\u2_Display/n5154 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_0  (
    .a(\u2_Display/n6346 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c0 ),
    .o({\u2_Display/lt162_c1 ,open_n2918}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_1  (
    .a(\u2_Display/n6345 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c1 ),
    .o({\u2_Display/lt162_c2 ,open_n2919}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_10  (
    .a(\u2_Display/n6336 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c10 ),
    .o({\u2_Display/lt162_c11 ,open_n2920}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_11  (
    .a(\u2_Display/n6335 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c11 ),
    .o({\u2_Display/lt162_c12 ,open_n2921}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_12  (
    .a(\u2_Display/n6334 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c12 ),
    .o({\u2_Display/lt162_c13 ,open_n2922}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_13  (
    .a(\u2_Display/n6333 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c13 ),
    .o({\u2_Display/lt162_c14 ,open_n2923}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_14  (
    .a(\u2_Display/n6332 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c14 ),
    .o({\u2_Display/lt162_c15 ,open_n2924}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_15  (
    .a(\u2_Display/n6331 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c15 ),
    .o({\u2_Display/lt162_c16 ,open_n2925}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_16  (
    .a(\u2_Display/n6330 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c16 ),
    .o({\u2_Display/lt162_c17 ,open_n2926}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_17  (
    .a(\u2_Display/n6329 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c17 ),
    .o({\u2_Display/lt162_c18 ,open_n2927}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_18  (
    .a(\u2_Display/n6328 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c18 ),
    .o({\u2_Display/lt162_c19 ,open_n2928}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_19  (
    .a(\u2_Display/n6327 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c19 ),
    .o({\u2_Display/lt162_c20 ,open_n2929}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_2  (
    .a(\u2_Display/n6344 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c2 ),
    .o({\u2_Display/lt162_c3 ,open_n2930}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_20  (
    .a(\u2_Display/n6326 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c20 ),
    .o({\u2_Display/lt162_c21 ,open_n2931}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_21  (
    .a(\u2_Display/n6325 ),
    .b(1'b1),
    .c(\u2_Display/lt162_c21 ),
    .o({\u2_Display/lt162_c22 ,open_n2932}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_22  (
    .a(\u2_Display/n6324 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c22 ),
    .o({\u2_Display/lt162_c23 ,open_n2933}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_23  (
    .a(\u2_Display/n6323 ),
    .b(1'b1),
    .c(\u2_Display/lt162_c23 ),
    .o({\u2_Display/lt162_c24 ,open_n2934}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_24  (
    .a(\u2_Display/n6322 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c24 ),
    .o({\u2_Display/lt162_c25 ,open_n2935}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_25  (
    .a(\u2_Display/n6321 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c25 ),
    .o({\u2_Display/lt162_c26 ,open_n2936}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_26  (
    .a(\u2_Display/n6320 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c26 ),
    .o({\u2_Display/lt162_c27 ,open_n2937}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_27  (
    .a(\u2_Display/n6319 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c27 ),
    .o({\u2_Display/lt162_c28 ,open_n2938}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_28  (
    .a(\u2_Display/n6318 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c28 ),
    .o({\u2_Display/lt162_c29 ,open_n2939}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_29  (
    .a(\u2_Display/n6317 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c29 ),
    .o({\u2_Display/lt162_c30 ,open_n2940}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_3  (
    .a(\u2_Display/n6343 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c3 ),
    .o({\u2_Display/lt162_c4 ,open_n2941}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_30  (
    .a(\u2_Display/n6316 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c30 ),
    .o({\u2_Display/lt162_c31 ,open_n2942}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_31  (
    .a(\u2_Display/n6315 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c31 ),
    .o({\u2_Display/lt162_c32 ,open_n2943}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_4  (
    .a(\u2_Display/n6342 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c4 ),
    .o({\u2_Display/lt162_c5 ,open_n2944}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_5  (
    .a(\u2_Display/n6341 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c5 ),
    .o({\u2_Display/lt162_c6 ,open_n2945}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_6  (
    .a(\u2_Display/n6340 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c6 ),
    .o({\u2_Display/lt162_c7 ,open_n2946}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_7  (
    .a(\u2_Display/n6339 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c7 ),
    .o({\u2_Display/lt162_c8 ,open_n2947}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_8  (
    .a(\u2_Display/n6338 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c8 ),
    .o({\u2_Display/lt162_c9 ,open_n2948}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_9  (
    .a(\u2_Display/n6337 ),
    .b(1'b0),
    .c(\u2_Display/lt162_c9 ),
    .o({\u2_Display/lt162_c10 ,open_n2949}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt162_cin  (
    .a(1'b0),
    .o({\u2_Display/lt162_c0 ,open_n2952}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt162_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt162_c32 ),
    .o({open_n2953,\u2_Display/n5189 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_0  (
    .a(\u2_Display/n5223 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c0 ),
    .o({\u2_Display/lt163_c1 ,open_n2954}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_1  (
    .a(\u2_Display/n5222 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c1 ),
    .o({\u2_Display/lt163_c2 ,open_n2955}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_10  (
    .a(\u2_Display/n5213 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c10 ),
    .o({\u2_Display/lt163_c11 ,open_n2956}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_11  (
    .a(\u2_Display/n5212 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c11 ),
    .o({\u2_Display/lt163_c12 ,open_n2957}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_12  (
    .a(\u2_Display/n5211 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c12 ),
    .o({\u2_Display/lt163_c13 ,open_n2958}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_13  (
    .a(\u2_Display/n5210 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c13 ),
    .o({\u2_Display/lt163_c14 ,open_n2959}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_14  (
    .a(\u2_Display/n5209 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c14 ),
    .o({\u2_Display/lt163_c15 ,open_n2960}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_15  (
    .a(\u2_Display/n5208 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c15 ),
    .o({\u2_Display/lt163_c16 ,open_n2961}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_16  (
    .a(\u2_Display/n5207 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c16 ),
    .o({\u2_Display/lt163_c17 ,open_n2962}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_17  (
    .a(\u2_Display/n5206 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c17 ),
    .o({\u2_Display/lt163_c18 ,open_n2963}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_18  (
    .a(\u2_Display/n5205 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c18 ),
    .o({\u2_Display/lt163_c19 ,open_n2964}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_19  (
    .a(\u2_Display/n5204 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c19 ),
    .o({\u2_Display/lt163_c20 ,open_n2965}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_2  (
    .a(\u2_Display/n5221 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c2 ),
    .o({\u2_Display/lt163_c3 ,open_n2966}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_20  (
    .a(\u2_Display/n5203 ),
    .b(1'b1),
    .c(\u2_Display/lt163_c20 ),
    .o({\u2_Display/lt163_c21 ,open_n2967}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_21  (
    .a(\u2_Display/n5202 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c21 ),
    .o({\u2_Display/lt163_c22 ,open_n2968}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_22  (
    .a(\u2_Display/n5201 ),
    .b(1'b1),
    .c(\u2_Display/lt163_c22 ),
    .o({\u2_Display/lt163_c23 ,open_n2969}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_23  (
    .a(\u2_Display/n5200 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c23 ),
    .o({\u2_Display/lt163_c24 ,open_n2970}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_24  (
    .a(\u2_Display/n5199 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c24 ),
    .o({\u2_Display/lt163_c25 ,open_n2971}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_25  (
    .a(\u2_Display/n5198 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c25 ),
    .o({\u2_Display/lt163_c26 ,open_n2972}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_26  (
    .a(\u2_Display/n5197 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c26 ),
    .o({\u2_Display/lt163_c27 ,open_n2973}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_27  (
    .a(\u2_Display/n5196 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c27 ),
    .o({\u2_Display/lt163_c28 ,open_n2974}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_28  (
    .a(\u2_Display/n6353 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c28 ),
    .o({\u2_Display/lt163_c29 ,open_n2975}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_29  (
    .a(\u2_Display/n6352 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c29 ),
    .o({\u2_Display/lt163_c30 ,open_n2976}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_3  (
    .a(\u2_Display/n5220 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c3 ),
    .o({\u2_Display/lt163_c4 ,open_n2977}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_30  (
    .a(\u2_Display/n6351 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c30 ),
    .o({\u2_Display/lt163_c31 ,open_n2978}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_31  (
    .a(\u2_Display/n6350 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c31 ),
    .o({\u2_Display/lt163_c32 ,open_n2979}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_4  (
    .a(\u2_Display/n5219 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c4 ),
    .o({\u2_Display/lt163_c5 ,open_n2980}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_5  (
    .a(\u2_Display/n5218 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c5 ),
    .o({\u2_Display/lt163_c6 ,open_n2981}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_6  (
    .a(\u2_Display/n5217 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c6 ),
    .o({\u2_Display/lt163_c7 ,open_n2982}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_7  (
    .a(\u2_Display/n5216 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c7 ),
    .o({\u2_Display/lt163_c8 ,open_n2983}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_8  (
    .a(\u2_Display/n5215 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c8 ),
    .o({\u2_Display/lt163_c9 ,open_n2984}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_9  (
    .a(\u2_Display/n5214 ),
    .b(1'b0),
    .c(\u2_Display/lt163_c9 ),
    .o({\u2_Display/lt163_c10 ,open_n2985}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt163_cin  (
    .a(1'b0),
    .o({\u2_Display/lt163_c0 ,open_n2988}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt163_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt163_c32 ),
    .o({open_n2989,\u2_Display/n5224 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_0  (
    .a(\u2_Display/n5258 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c0 ),
    .o({\u2_Display/lt164_c1 ,open_n2990}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_1  (
    .a(\u2_Display/n5257 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c1 ),
    .o({\u2_Display/lt164_c2 ,open_n2991}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_10  (
    .a(\u2_Display/n5248 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c10 ),
    .o({\u2_Display/lt164_c11 ,open_n2992}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_11  (
    .a(\u2_Display/n5247 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c11 ),
    .o({\u2_Display/lt164_c12 ,open_n2993}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_12  (
    .a(\u2_Display/n5246 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c12 ),
    .o({\u2_Display/lt164_c13 ,open_n2994}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_13  (
    .a(\u2_Display/n5245 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c13 ),
    .o({\u2_Display/lt164_c14 ,open_n2995}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_14  (
    .a(\u2_Display/n5244 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c14 ),
    .o({\u2_Display/lt164_c15 ,open_n2996}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_15  (
    .a(\u2_Display/n5243 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c15 ),
    .o({\u2_Display/lt164_c16 ,open_n2997}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_16  (
    .a(\u2_Display/n5242 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c16 ),
    .o({\u2_Display/lt164_c17 ,open_n2998}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_17  (
    .a(\u2_Display/n5241 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c17 ),
    .o({\u2_Display/lt164_c18 ,open_n2999}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_18  (
    .a(\u2_Display/n5240 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c18 ),
    .o({\u2_Display/lt164_c19 ,open_n3000}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_19  (
    .a(\u2_Display/n5239 ),
    .b(1'b1),
    .c(\u2_Display/lt164_c19 ),
    .o({\u2_Display/lt164_c20 ,open_n3001}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_2  (
    .a(\u2_Display/n5256 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c2 ),
    .o({\u2_Display/lt164_c3 ,open_n3002}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_20  (
    .a(\u2_Display/n5238 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c20 ),
    .o({\u2_Display/lt164_c21 ,open_n3003}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_21  (
    .a(\u2_Display/n5237 ),
    .b(1'b1),
    .c(\u2_Display/lt164_c21 ),
    .o({\u2_Display/lt164_c22 ,open_n3004}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_22  (
    .a(\u2_Display/n5236 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c22 ),
    .o({\u2_Display/lt164_c23 ,open_n3005}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_23  (
    .a(\u2_Display/n5235 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c23 ),
    .o({\u2_Display/lt164_c24 ,open_n3006}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_24  (
    .a(\u2_Display/n5234 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c24 ),
    .o({\u2_Display/lt164_c25 ,open_n3007}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_25  (
    .a(\u2_Display/n5233 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c25 ),
    .o({\u2_Display/lt164_c26 ,open_n3008}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_26  (
    .a(\u2_Display/n5232 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c26 ),
    .o({\u2_Display/lt164_c27 ,open_n3009}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_27  (
    .a(\u2_Display/n5231 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c27 ),
    .o({\u2_Display/lt164_c28 ,open_n3010}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_28  (
    .a(\u2_Display/n5230 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c28 ),
    .o({\u2_Display/lt164_c29 ,open_n3011}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_29  (
    .a(\u2_Display/n5229 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c29 ),
    .o({\u2_Display/lt164_c30 ,open_n3012}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_3  (
    .a(\u2_Display/n5255 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c3 ),
    .o({\u2_Display/lt164_c4 ,open_n3013}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_30  (
    .a(\u2_Display/n5228 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c30 ),
    .o({\u2_Display/lt164_c31 ,open_n3014}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_31  (
    .a(\u2_Display/n5227 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c31 ),
    .o({\u2_Display/lt164_c32 ,open_n3015}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_4  (
    .a(\u2_Display/n5254 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c4 ),
    .o({\u2_Display/lt164_c5 ,open_n3016}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_5  (
    .a(\u2_Display/n5253 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c5 ),
    .o({\u2_Display/lt164_c6 ,open_n3017}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_6  (
    .a(\u2_Display/n5252 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c6 ),
    .o({\u2_Display/lt164_c7 ,open_n3018}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_7  (
    .a(\u2_Display/n5251 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c7 ),
    .o({\u2_Display/lt164_c8 ,open_n3019}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_8  (
    .a(\u2_Display/n5250 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c8 ),
    .o({\u2_Display/lt164_c9 ,open_n3020}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_9  (
    .a(\u2_Display/n5249 ),
    .b(1'b0),
    .c(\u2_Display/lt164_c9 ),
    .o({\u2_Display/lt164_c10 ,open_n3021}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt164_cin  (
    .a(1'b0),
    .o({\u2_Display/lt164_c0 ,open_n3024}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt164_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt164_c32 ),
    .o({open_n3025,\u2_Display/n5259 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_0  (
    .a(\u2_Display/n5293 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c0 ),
    .o({\u2_Display/lt165_c1 ,open_n3026}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_1  (
    .a(\u2_Display/n5292 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c1 ),
    .o({\u2_Display/lt165_c2 ,open_n3027}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_10  (
    .a(\u2_Display/n5283 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c10 ),
    .o({\u2_Display/lt165_c11 ,open_n3028}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_11  (
    .a(\u2_Display/n5282 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c11 ),
    .o({\u2_Display/lt165_c12 ,open_n3029}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_12  (
    .a(\u2_Display/n5281 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c12 ),
    .o({\u2_Display/lt165_c13 ,open_n3030}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_13  (
    .a(\u2_Display/n5280 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c13 ),
    .o({\u2_Display/lt165_c14 ,open_n3031}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_14  (
    .a(\u2_Display/n5279 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c14 ),
    .o({\u2_Display/lt165_c15 ,open_n3032}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_15  (
    .a(\u2_Display/n5278 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c15 ),
    .o({\u2_Display/lt165_c16 ,open_n3033}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_16  (
    .a(\u2_Display/n5277 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c16 ),
    .o({\u2_Display/lt165_c17 ,open_n3034}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_17  (
    .a(\u2_Display/n5276 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c17 ),
    .o({\u2_Display/lt165_c18 ,open_n3035}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_18  (
    .a(\u2_Display/n5275 ),
    .b(1'b1),
    .c(\u2_Display/lt165_c18 ),
    .o({\u2_Display/lt165_c19 ,open_n3036}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_19  (
    .a(\u2_Display/n5274 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c19 ),
    .o({\u2_Display/lt165_c20 ,open_n3037}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_2  (
    .a(\u2_Display/n5291 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c2 ),
    .o({\u2_Display/lt165_c3 ,open_n3038}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_20  (
    .a(\u2_Display/n5273 ),
    .b(1'b1),
    .c(\u2_Display/lt165_c20 ),
    .o({\u2_Display/lt165_c21 ,open_n3039}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_21  (
    .a(\u2_Display/n5272 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c21 ),
    .o({\u2_Display/lt165_c22 ,open_n3040}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_22  (
    .a(\u2_Display/n5271 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c22 ),
    .o({\u2_Display/lt165_c23 ,open_n3041}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_23  (
    .a(\u2_Display/n5270 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c23 ),
    .o({\u2_Display/lt165_c24 ,open_n3042}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_24  (
    .a(\u2_Display/n5269 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c24 ),
    .o({\u2_Display/lt165_c25 ,open_n3043}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_25  (
    .a(\u2_Display/n5268 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c25 ),
    .o({\u2_Display/lt165_c26 ,open_n3044}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_26  (
    .a(\u2_Display/n5267 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c26 ),
    .o({\u2_Display/lt165_c27 ,open_n3045}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_27  (
    .a(\u2_Display/n5266 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c27 ),
    .o({\u2_Display/lt165_c28 ,open_n3046}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_28  (
    .a(\u2_Display/n5265 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c28 ),
    .o({\u2_Display/lt165_c29 ,open_n3047}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_29  (
    .a(\u2_Display/n5264 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c29 ),
    .o({\u2_Display/lt165_c30 ,open_n3048}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_3  (
    .a(\u2_Display/n5290 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c3 ),
    .o({\u2_Display/lt165_c4 ,open_n3049}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_30  (
    .a(\u2_Display/n5263 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c30 ),
    .o({\u2_Display/lt165_c31 ,open_n3050}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_31  (
    .a(\u2_Display/n5262 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c31 ),
    .o({\u2_Display/lt165_c32 ,open_n3051}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_4  (
    .a(\u2_Display/n5289 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c4 ),
    .o({\u2_Display/lt165_c5 ,open_n3052}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_5  (
    .a(\u2_Display/n5288 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c5 ),
    .o({\u2_Display/lt165_c6 ,open_n3053}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_6  (
    .a(\u2_Display/n5287 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c6 ),
    .o({\u2_Display/lt165_c7 ,open_n3054}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_7  (
    .a(\u2_Display/n5286 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c7 ),
    .o({\u2_Display/lt165_c8 ,open_n3055}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_8  (
    .a(\u2_Display/n5285 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c8 ),
    .o({\u2_Display/lt165_c9 ,open_n3056}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_9  (
    .a(\u2_Display/n5284 ),
    .b(1'b0),
    .c(\u2_Display/lt165_c9 ),
    .o({\u2_Display/lt165_c10 ,open_n3057}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt165_cin  (
    .a(1'b0),
    .o({\u2_Display/lt165_c0 ,open_n3060}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt165_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt165_c32 ),
    .o({open_n3061,\u2_Display/n5294 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_0  (
    .a(\u2_Display/n5328 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c0 ),
    .o({\u2_Display/lt166_c1 ,open_n3062}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_1  (
    .a(\u2_Display/n5327 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c1 ),
    .o({\u2_Display/lt166_c2 ,open_n3063}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_10  (
    .a(\u2_Display/n5318 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c10 ),
    .o({\u2_Display/lt166_c11 ,open_n3064}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_11  (
    .a(\u2_Display/n5317 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c11 ),
    .o({\u2_Display/lt166_c12 ,open_n3065}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_12  (
    .a(\u2_Display/n5316 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c12 ),
    .o({\u2_Display/lt166_c13 ,open_n3066}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_13  (
    .a(\u2_Display/n5315 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c13 ),
    .o({\u2_Display/lt166_c14 ,open_n3067}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_14  (
    .a(\u2_Display/n5314 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c14 ),
    .o({\u2_Display/lt166_c15 ,open_n3068}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_15  (
    .a(\u2_Display/n5313 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c15 ),
    .o({\u2_Display/lt166_c16 ,open_n3069}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_16  (
    .a(\u2_Display/n5312 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c16 ),
    .o({\u2_Display/lt166_c17 ,open_n3070}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_17  (
    .a(\u2_Display/n5311 ),
    .b(1'b1),
    .c(\u2_Display/lt166_c17 ),
    .o({\u2_Display/lt166_c18 ,open_n3071}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_18  (
    .a(\u2_Display/n5310 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c18 ),
    .o({\u2_Display/lt166_c19 ,open_n3072}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_19  (
    .a(\u2_Display/n5309 ),
    .b(1'b1),
    .c(\u2_Display/lt166_c19 ),
    .o({\u2_Display/lt166_c20 ,open_n3073}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_2  (
    .a(\u2_Display/n5326 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c2 ),
    .o({\u2_Display/lt166_c3 ,open_n3074}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_20  (
    .a(\u2_Display/n5308 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c20 ),
    .o({\u2_Display/lt166_c21 ,open_n3075}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_21  (
    .a(\u2_Display/n5307 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c21 ),
    .o({\u2_Display/lt166_c22 ,open_n3076}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_22  (
    .a(\u2_Display/n5306 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c22 ),
    .o({\u2_Display/lt166_c23 ,open_n3077}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_23  (
    .a(\u2_Display/n5305 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c23 ),
    .o({\u2_Display/lt166_c24 ,open_n3078}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_24  (
    .a(\u2_Display/n5304 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c24 ),
    .o({\u2_Display/lt166_c25 ,open_n3079}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_25  (
    .a(\u2_Display/n5303 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c25 ),
    .o({\u2_Display/lt166_c26 ,open_n3080}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_26  (
    .a(\u2_Display/n5302 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c26 ),
    .o({\u2_Display/lt166_c27 ,open_n3081}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_27  (
    .a(\u2_Display/n5301 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c27 ),
    .o({\u2_Display/lt166_c28 ,open_n3082}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_28  (
    .a(\u2_Display/n5300 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c28 ),
    .o({\u2_Display/lt166_c29 ,open_n3083}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_29  (
    .a(\u2_Display/n5299 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c29 ),
    .o({\u2_Display/lt166_c30 ,open_n3084}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_3  (
    .a(\u2_Display/n5325 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c3 ),
    .o({\u2_Display/lt166_c4 ,open_n3085}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_30  (
    .a(\u2_Display/n5298 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c30 ),
    .o({\u2_Display/lt166_c31 ,open_n3086}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_31  (
    .a(\u2_Display/n5297 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c31 ),
    .o({\u2_Display/lt166_c32 ,open_n3087}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_4  (
    .a(\u2_Display/n5324 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c4 ),
    .o({\u2_Display/lt166_c5 ,open_n3088}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_5  (
    .a(\u2_Display/n5323 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c5 ),
    .o({\u2_Display/lt166_c6 ,open_n3089}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_6  (
    .a(\u2_Display/n5322 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c6 ),
    .o({\u2_Display/lt166_c7 ,open_n3090}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_7  (
    .a(\u2_Display/n5321 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c7 ),
    .o({\u2_Display/lt166_c8 ,open_n3091}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_8  (
    .a(\u2_Display/n5320 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c8 ),
    .o({\u2_Display/lt166_c9 ,open_n3092}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_9  (
    .a(\u2_Display/n5319 ),
    .b(1'b0),
    .c(\u2_Display/lt166_c9 ),
    .o({\u2_Display/lt166_c10 ,open_n3093}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt166_cin  (
    .a(1'b0),
    .o({\u2_Display/lt166_c0 ,open_n3096}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt166_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt166_c32 ),
    .o({open_n3097,\u2_Display/n5329 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_0  (
    .a(\u2_Display/n5363 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c0 ),
    .o({\u2_Display/lt167_c1 ,open_n3098}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_1  (
    .a(\u2_Display/n5362 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c1 ),
    .o({\u2_Display/lt167_c2 ,open_n3099}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_10  (
    .a(\u2_Display/n5353 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c10 ),
    .o({\u2_Display/lt167_c11 ,open_n3100}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_11  (
    .a(\u2_Display/n5352 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c11 ),
    .o({\u2_Display/lt167_c12 ,open_n3101}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_12  (
    .a(\u2_Display/n5351 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c12 ),
    .o({\u2_Display/lt167_c13 ,open_n3102}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_13  (
    .a(\u2_Display/n5350 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c13 ),
    .o({\u2_Display/lt167_c14 ,open_n3103}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_14  (
    .a(\u2_Display/n5349 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c14 ),
    .o({\u2_Display/lt167_c15 ,open_n3104}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_15  (
    .a(\u2_Display/n5348 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c15 ),
    .o({\u2_Display/lt167_c16 ,open_n3105}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_16  (
    .a(\u2_Display/n5347 ),
    .b(1'b1),
    .c(\u2_Display/lt167_c16 ),
    .o({\u2_Display/lt167_c17 ,open_n3106}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_17  (
    .a(\u2_Display/n5346 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c17 ),
    .o({\u2_Display/lt167_c18 ,open_n3107}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_18  (
    .a(\u2_Display/n5345 ),
    .b(1'b1),
    .c(\u2_Display/lt167_c18 ),
    .o({\u2_Display/lt167_c19 ,open_n3108}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_19  (
    .a(\u2_Display/n5344 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c19 ),
    .o({\u2_Display/lt167_c20 ,open_n3109}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_2  (
    .a(\u2_Display/n5361 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c2 ),
    .o({\u2_Display/lt167_c3 ,open_n3110}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_20  (
    .a(\u2_Display/n5343 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c20 ),
    .o({\u2_Display/lt167_c21 ,open_n3111}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_21  (
    .a(\u2_Display/n5342 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c21 ),
    .o({\u2_Display/lt167_c22 ,open_n3112}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_22  (
    .a(\u2_Display/n5341 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c22 ),
    .o({\u2_Display/lt167_c23 ,open_n3113}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_23  (
    .a(\u2_Display/n5340 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c23 ),
    .o({\u2_Display/lt167_c24 ,open_n3114}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_24  (
    .a(\u2_Display/n5339 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c24 ),
    .o({\u2_Display/lt167_c25 ,open_n3115}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_25  (
    .a(\u2_Display/n5338 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c25 ),
    .o({\u2_Display/lt167_c26 ,open_n3116}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_26  (
    .a(\u2_Display/n5337 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c26 ),
    .o({\u2_Display/lt167_c27 ,open_n3117}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_27  (
    .a(\u2_Display/n5336 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c27 ),
    .o({\u2_Display/lt167_c28 ,open_n3118}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_28  (
    .a(\u2_Display/n5335 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c28 ),
    .o({\u2_Display/lt167_c29 ,open_n3119}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_29  (
    .a(\u2_Display/n5334 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c29 ),
    .o({\u2_Display/lt167_c30 ,open_n3120}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_3  (
    .a(\u2_Display/n5360 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c3 ),
    .o({\u2_Display/lt167_c4 ,open_n3121}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_30  (
    .a(\u2_Display/n5333 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c30 ),
    .o({\u2_Display/lt167_c31 ,open_n3122}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_31  (
    .a(\u2_Display/n5332 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c31 ),
    .o({\u2_Display/lt167_c32 ,open_n3123}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_4  (
    .a(\u2_Display/n5359 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c4 ),
    .o({\u2_Display/lt167_c5 ,open_n3124}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_5  (
    .a(\u2_Display/n5358 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c5 ),
    .o({\u2_Display/lt167_c6 ,open_n3125}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_6  (
    .a(\u2_Display/n5357 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c6 ),
    .o({\u2_Display/lt167_c7 ,open_n3126}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_7  (
    .a(\u2_Display/n5356 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c7 ),
    .o({\u2_Display/lt167_c8 ,open_n3127}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_8  (
    .a(\u2_Display/n5355 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c8 ),
    .o({\u2_Display/lt167_c9 ,open_n3128}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_9  (
    .a(\u2_Display/n5354 ),
    .b(1'b0),
    .c(\u2_Display/lt167_c9 ),
    .o({\u2_Display/lt167_c10 ,open_n3129}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt167_cin  (
    .a(1'b0),
    .o({\u2_Display/lt167_c0 ,open_n3132}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt167_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt167_c32 ),
    .o({open_n3133,\u2_Display/n5364 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_0  (
    .a(\u2_Display/n5398 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c0 ),
    .o({\u2_Display/lt168_c1 ,open_n3134}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_1  (
    .a(\u2_Display/n5397 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c1 ),
    .o({\u2_Display/lt168_c2 ,open_n3135}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_10  (
    .a(\u2_Display/n5388 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c10 ),
    .o({\u2_Display/lt168_c11 ,open_n3136}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_11  (
    .a(\u2_Display/n5387 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c11 ),
    .o({\u2_Display/lt168_c12 ,open_n3137}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_12  (
    .a(\u2_Display/n5386 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c12 ),
    .o({\u2_Display/lt168_c13 ,open_n3138}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_13  (
    .a(\u2_Display/n5385 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c13 ),
    .o({\u2_Display/lt168_c14 ,open_n3139}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_14  (
    .a(\u2_Display/n5384 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c14 ),
    .o({\u2_Display/lt168_c15 ,open_n3140}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_15  (
    .a(\u2_Display/n5383 ),
    .b(1'b1),
    .c(\u2_Display/lt168_c15 ),
    .o({\u2_Display/lt168_c16 ,open_n3141}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_16  (
    .a(\u2_Display/n5382 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c16 ),
    .o({\u2_Display/lt168_c17 ,open_n3142}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_17  (
    .a(\u2_Display/n5381 ),
    .b(1'b1),
    .c(\u2_Display/lt168_c17 ),
    .o({\u2_Display/lt168_c18 ,open_n3143}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_18  (
    .a(\u2_Display/n5380 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c18 ),
    .o({\u2_Display/lt168_c19 ,open_n3144}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_19  (
    .a(\u2_Display/n5379 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c19 ),
    .o({\u2_Display/lt168_c20 ,open_n3145}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_2  (
    .a(\u2_Display/n5396 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c2 ),
    .o({\u2_Display/lt168_c3 ,open_n3146}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_20  (
    .a(\u2_Display/n5378 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c20 ),
    .o({\u2_Display/lt168_c21 ,open_n3147}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_21  (
    .a(\u2_Display/n5377 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c21 ),
    .o({\u2_Display/lt168_c22 ,open_n3148}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_22  (
    .a(\u2_Display/n5376 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c22 ),
    .o({\u2_Display/lt168_c23 ,open_n3149}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_23  (
    .a(\u2_Display/n5375 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c23 ),
    .o({\u2_Display/lt168_c24 ,open_n3150}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_24  (
    .a(\u2_Display/n5374 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c24 ),
    .o({\u2_Display/lt168_c25 ,open_n3151}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_25  (
    .a(\u2_Display/n5373 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c25 ),
    .o({\u2_Display/lt168_c26 ,open_n3152}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_26  (
    .a(\u2_Display/n5372 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c26 ),
    .o({\u2_Display/lt168_c27 ,open_n3153}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_27  (
    .a(\u2_Display/n5371 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c27 ),
    .o({\u2_Display/lt168_c28 ,open_n3154}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_28  (
    .a(\u2_Display/n5370 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c28 ),
    .o({\u2_Display/lt168_c29 ,open_n3155}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_29  (
    .a(\u2_Display/n5369 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c29 ),
    .o({\u2_Display/lt168_c30 ,open_n3156}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_3  (
    .a(\u2_Display/n5395 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c3 ),
    .o({\u2_Display/lt168_c4 ,open_n3157}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_30  (
    .a(\u2_Display/n5368 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c30 ),
    .o({\u2_Display/lt168_c31 ,open_n3158}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_31  (
    .a(\u2_Display/n5367 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c31 ),
    .o({\u2_Display/lt168_c32 ,open_n3159}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_4  (
    .a(\u2_Display/n5394 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c4 ),
    .o({\u2_Display/lt168_c5 ,open_n3160}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_5  (
    .a(\u2_Display/n5393 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c5 ),
    .o({\u2_Display/lt168_c6 ,open_n3161}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_6  (
    .a(\u2_Display/n5392 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c6 ),
    .o({\u2_Display/lt168_c7 ,open_n3162}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_7  (
    .a(\u2_Display/n5391 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c7 ),
    .o({\u2_Display/lt168_c8 ,open_n3163}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_8  (
    .a(\u2_Display/n5390 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c8 ),
    .o({\u2_Display/lt168_c9 ,open_n3164}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_9  (
    .a(\u2_Display/n5389 ),
    .b(1'b0),
    .c(\u2_Display/lt168_c9 ),
    .o({\u2_Display/lt168_c10 ,open_n3165}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt168_cin  (
    .a(1'b0),
    .o({\u2_Display/lt168_c0 ,open_n3168}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt168_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt168_c32 ),
    .o({open_n3169,\u2_Display/n5399 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_0  (
    .a(\u2_Display/n5433 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c0 ),
    .o({\u2_Display/lt169_c1 ,open_n3170}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_1  (
    .a(\u2_Display/n5432 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c1 ),
    .o({\u2_Display/lt169_c2 ,open_n3171}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_10  (
    .a(\u2_Display/n5423 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c10 ),
    .o({\u2_Display/lt169_c11 ,open_n3172}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_11  (
    .a(\u2_Display/n5422 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c11 ),
    .o({\u2_Display/lt169_c12 ,open_n3173}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_12  (
    .a(\u2_Display/n5421 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c12 ),
    .o({\u2_Display/lt169_c13 ,open_n3174}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_13  (
    .a(\u2_Display/n5420 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c13 ),
    .o({\u2_Display/lt169_c14 ,open_n3175}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_14  (
    .a(\u2_Display/n5419 ),
    .b(1'b1),
    .c(\u2_Display/lt169_c14 ),
    .o({\u2_Display/lt169_c15 ,open_n3176}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_15  (
    .a(\u2_Display/n5418 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c15 ),
    .o({\u2_Display/lt169_c16 ,open_n3177}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_16  (
    .a(\u2_Display/n5417 ),
    .b(1'b1),
    .c(\u2_Display/lt169_c16 ),
    .o({\u2_Display/lt169_c17 ,open_n3178}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_17  (
    .a(\u2_Display/n5416 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c17 ),
    .o({\u2_Display/lt169_c18 ,open_n3179}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_18  (
    .a(\u2_Display/n5415 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c18 ),
    .o({\u2_Display/lt169_c19 ,open_n3180}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_19  (
    .a(\u2_Display/n5414 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c19 ),
    .o({\u2_Display/lt169_c20 ,open_n3181}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_2  (
    .a(\u2_Display/n5431 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c2 ),
    .o({\u2_Display/lt169_c3 ,open_n3182}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_20  (
    .a(\u2_Display/n5413 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c20 ),
    .o({\u2_Display/lt169_c21 ,open_n3183}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_21  (
    .a(\u2_Display/n5412 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c21 ),
    .o({\u2_Display/lt169_c22 ,open_n3184}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_22  (
    .a(\u2_Display/n5411 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c22 ),
    .o({\u2_Display/lt169_c23 ,open_n3185}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_23  (
    .a(\u2_Display/n5410 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c23 ),
    .o({\u2_Display/lt169_c24 ,open_n3186}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_24  (
    .a(\u2_Display/n5409 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c24 ),
    .o({\u2_Display/lt169_c25 ,open_n3187}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_25  (
    .a(\u2_Display/n5408 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c25 ),
    .o({\u2_Display/lt169_c26 ,open_n3188}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_26  (
    .a(\u2_Display/n5407 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c26 ),
    .o({\u2_Display/lt169_c27 ,open_n3189}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_27  (
    .a(\u2_Display/n5406 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c27 ),
    .o({\u2_Display/lt169_c28 ,open_n3190}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_28  (
    .a(\u2_Display/n5405 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c28 ),
    .o({\u2_Display/lt169_c29 ,open_n3191}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_29  (
    .a(\u2_Display/n5404 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c29 ),
    .o({\u2_Display/lt169_c30 ,open_n3192}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_3  (
    .a(\u2_Display/n5430 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c3 ),
    .o({\u2_Display/lt169_c4 ,open_n3193}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_30  (
    .a(\u2_Display/n5403 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c30 ),
    .o({\u2_Display/lt169_c31 ,open_n3194}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_31  (
    .a(\u2_Display/n5402 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c31 ),
    .o({\u2_Display/lt169_c32 ,open_n3195}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_4  (
    .a(\u2_Display/n5429 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c4 ),
    .o({\u2_Display/lt169_c5 ,open_n3196}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_5  (
    .a(\u2_Display/n5428 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c5 ),
    .o({\u2_Display/lt169_c6 ,open_n3197}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_6  (
    .a(\u2_Display/n5427 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c6 ),
    .o({\u2_Display/lt169_c7 ,open_n3198}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_7  (
    .a(\u2_Display/n5426 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c7 ),
    .o({\u2_Display/lt169_c8 ,open_n3199}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_8  (
    .a(\u2_Display/n5425 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c8 ),
    .o({\u2_Display/lt169_c9 ,open_n3200}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_9  (
    .a(\u2_Display/n5424 ),
    .b(1'b0),
    .c(\u2_Display/lt169_c9 ),
    .o({\u2_Display/lt169_c10 ,open_n3201}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt169_cin  (
    .a(1'b0),
    .o({\u2_Display/lt169_c0 ,open_n3204}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt169_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt169_c32 ),
    .o({open_n3205,\u2_Display/n5434 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_0  (
    .a(\u2_Display/n5468 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c0 ),
    .o({\u2_Display/lt170_c1 ,open_n3206}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_1  (
    .a(\u2_Display/n5467 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c1 ),
    .o({\u2_Display/lt170_c2 ,open_n3207}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_10  (
    .a(\u2_Display/n5458 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c10 ),
    .o({\u2_Display/lt170_c11 ,open_n3208}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_11  (
    .a(\u2_Display/n5457 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c11 ),
    .o({\u2_Display/lt170_c12 ,open_n3209}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_12  (
    .a(\u2_Display/n5456 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c12 ),
    .o({\u2_Display/lt170_c13 ,open_n3210}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_13  (
    .a(\u2_Display/n5455 ),
    .b(1'b1),
    .c(\u2_Display/lt170_c13 ),
    .o({\u2_Display/lt170_c14 ,open_n3211}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_14  (
    .a(\u2_Display/n5454 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c14 ),
    .o({\u2_Display/lt170_c15 ,open_n3212}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_15  (
    .a(\u2_Display/n5453 ),
    .b(1'b1),
    .c(\u2_Display/lt170_c15 ),
    .o({\u2_Display/lt170_c16 ,open_n3213}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_16  (
    .a(\u2_Display/n5452 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c16 ),
    .o({\u2_Display/lt170_c17 ,open_n3214}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_17  (
    .a(\u2_Display/n5451 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c17 ),
    .o({\u2_Display/lt170_c18 ,open_n3215}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_18  (
    .a(\u2_Display/n5450 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c18 ),
    .o({\u2_Display/lt170_c19 ,open_n3216}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_19  (
    .a(\u2_Display/n5449 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c19 ),
    .o({\u2_Display/lt170_c20 ,open_n3217}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_2  (
    .a(\u2_Display/n5466 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c2 ),
    .o({\u2_Display/lt170_c3 ,open_n3218}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_20  (
    .a(\u2_Display/n5448 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c20 ),
    .o({\u2_Display/lt170_c21 ,open_n3219}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_21  (
    .a(\u2_Display/n5447 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c21 ),
    .o({\u2_Display/lt170_c22 ,open_n3220}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_22  (
    .a(\u2_Display/n5446 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c22 ),
    .o({\u2_Display/lt170_c23 ,open_n3221}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_23  (
    .a(\u2_Display/n5445 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c23 ),
    .o({\u2_Display/lt170_c24 ,open_n3222}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_24  (
    .a(\u2_Display/n5444 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c24 ),
    .o({\u2_Display/lt170_c25 ,open_n3223}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_25  (
    .a(\u2_Display/n5443 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c25 ),
    .o({\u2_Display/lt170_c26 ,open_n3224}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_26  (
    .a(\u2_Display/n5442 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c26 ),
    .o({\u2_Display/lt170_c27 ,open_n3225}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_27  (
    .a(\u2_Display/n5441 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c27 ),
    .o({\u2_Display/lt170_c28 ,open_n3226}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_28  (
    .a(\u2_Display/n5440 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c28 ),
    .o({\u2_Display/lt170_c29 ,open_n3227}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_29  (
    .a(\u2_Display/n5439 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c29 ),
    .o({\u2_Display/lt170_c30 ,open_n3228}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_3  (
    .a(\u2_Display/n5465 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c3 ),
    .o({\u2_Display/lt170_c4 ,open_n3229}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_30  (
    .a(\u2_Display/n5438 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c30 ),
    .o({\u2_Display/lt170_c31 ,open_n3230}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_31  (
    .a(\u2_Display/n5437 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c31 ),
    .o({\u2_Display/lt170_c32 ,open_n3231}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_4  (
    .a(\u2_Display/n5464 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c4 ),
    .o({\u2_Display/lt170_c5 ,open_n3232}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_5  (
    .a(\u2_Display/n5463 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c5 ),
    .o({\u2_Display/lt170_c6 ,open_n3233}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_6  (
    .a(\u2_Display/n5462 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c6 ),
    .o({\u2_Display/lt170_c7 ,open_n3234}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_7  (
    .a(\u2_Display/n5461 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c7 ),
    .o({\u2_Display/lt170_c8 ,open_n3235}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_8  (
    .a(\u2_Display/n5460 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c8 ),
    .o({\u2_Display/lt170_c9 ,open_n3236}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_9  (
    .a(\u2_Display/n5459 ),
    .b(1'b0),
    .c(\u2_Display/lt170_c9 ),
    .o({\u2_Display/lt170_c10 ,open_n3237}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt170_cin  (
    .a(1'b0),
    .o({\u2_Display/lt170_c0 ,open_n3240}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt170_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt170_c32 ),
    .o({open_n3241,\u2_Display/n5469 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_0  (
    .a(\u2_Display/n5503 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c0 ),
    .o({\u2_Display/lt171_c1 ,open_n3242}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_1  (
    .a(\u2_Display/n5502 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c1 ),
    .o({\u2_Display/lt171_c2 ,open_n3243}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_10  (
    .a(\u2_Display/n5493 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c10 ),
    .o({\u2_Display/lt171_c11 ,open_n3244}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_11  (
    .a(\u2_Display/n5492 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c11 ),
    .o({\u2_Display/lt171_c12 ,open_n3245}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_12  (
    .a(\u2_Display/n5491 ),
    .b(1'b1),
    .c(\u2_Display/lt171_c12 ),
    .o({\u2_Display/lt171_c13 ,open_n3246}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_13  (
    .a(\u2_Display/n5490 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c13 ),
    .o({\u2_Display/lt171_c14 ,open_n3247}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_14  (
    .a(\u2_Display/n5489 ),
    .b(1'b1),
    .c(\u2_Display/lt171_c14 ),
    .o({\u2_Display/lt171_c15 ,open_n3248}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_15  (
    .a(\u2_Display/n5488 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c15 ),
    .o({\u2_Display/lt171_c16 ,open_n3249}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_16  (
    .a(\u2_Display/n5487 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c16 ),
    .o({\u2_Display/lt171_c17 ,open_n3250}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_17  (
    .a(\u2_Display/n5486 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c17 ),
    .o({\u2_Display/lt171_c18 ,open_n3251}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_18  (
    .a(\u2_Display/n5485 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c18 ),
    .o({\u2_Display/lt171_c19 ,open_n3252}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_19  (
    .a(\u2_Display/n5484 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c19 ),
    .o({\u2_Display/lt171_c20 ,open_n3253}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_2  (
    .a(\u2_Display/n5501 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c2 ),
    .o({\u2_Display/lt171_c3 ,open_n3254}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_20  (
    .a(\u2_Display/n5483 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c20 ),
    .o({\u2_Display/lt171_c21 ,open_n3255}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_21  (
    .a(\u2_Display/n5482 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c21 ),
    .o({\u2_Display/lt171_c22 ,open_n3256}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_22  (
    .a(\u2_Display/n5481 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c22 ),
    .o({\u2_Display/lt171_c23 ,open_n3257}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_23  (
    .a(\u2_Display/n5480 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c23 ),
    .o({\u2_Display/lt171_c24 ,open_n3258}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_24  (
    .a(\u2_Display/n5479 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c24 ),
    .o({\u2_Display/lt171_c25 ,open_n3259}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_25  (
    .a(\u2_Display/n5478 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c25 ),
    .o({\u2_Display/lt171_c26 ,open_n3260}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_26  (
    .a(\u2_Display/n5477 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c26 ),
    .o({\u2_Display/lt171_c27 ,open_n3261}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_27  (
    .a(\u2_Display/n5476 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c27 ),
    .o({\u2_Display/lt171_c28 ,open_n3262}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_28  (
    .a(\u2_Display/n5475 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c28 ),
    .o({\u2_Display/lt171_c29 ,open_n3263}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_29  (
    .a(\u2_Display/n5474 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c29 ),
    .o({\u2_Display/lt171_c30 ,open_n3264}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_3  (
    .a(\u2_Display/n5500 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c3 ),
    .o({\u2_Display/lt171_c4 ,open_n3265}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_30  (
    .a(\u2_Display/n5473 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c30 ),
    .o({\u2_Display/lt171_c31 ,open_n3266}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_31  (
    .a(\u2_Display/n5472 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c31 ),
    .o({\u2_Display/lt171_c32 ,open_n3267}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_4  (
    .a(\u2_Display/n5499 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c4 ),
    .o({\u2_Display/lt171_c5 ,open_n3268}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_5  (
    .a(\u2_Display/n5498 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c5 ),
    .o({\u2_Display/lt171_c6 ,open_n3269}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_6  (
    .a(\u2_Display/n5497 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c6 ),
    .o({\u2_Display/lt171_c7 ,open_n3270}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_7  (
    .a(\u2_Display/n5496 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c7 ),
    .o({\u2_Display/lt171_c8 ,open_n3271}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_8  (
    .a(\u2_Display/n5495 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c8 ),
    .o({\u2_Display/lt171_c9 ,open_n3272}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_9  (
    .a(\u2_Display/n5494 ),
    .b(1'b0),
    .c(\u2_Display/lt171_c9 ),
    .o({\u2_Display/lt171_c10 ,open_n3273}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt171_cin  (
    .a(1'b0),
    .o({\u2_Display/lt171_c0 ,open_n3276}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt171_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt171_c32 ),
    .o({open_n3277,\u2_Display/n5504 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_0  (
    .a(\u2_Display/n5538 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c0 ),
    .o({\u2_Display/lt172_c1 ,open_n3278}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_1  (
    .a(\u2_Display/n5537 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c1 ),
    .o({\u2_Display/lt172_c2 ,open_n3279}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_10  (
    .a(\u2_Display/n5528 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c10 ),
    .o({\u2_Display/lt172_c11 ,open_n3280}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_11  (
    .a(\u2_Display/n5527 ),
    .b(1'b1),
    .c(\u2_Display/lt172_c11 ),
    .o({\u2_Display/lt172_c12 ,open_n3281}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_12  (
    .a(\u2_Display/n5526 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c12 ),
    .o({\u2_Display/lt172_c13 ,open_n3282}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_13  (
    .a(\u2_Display/n5525 ),
    .b(1'b1),
    .c(\u2_Display/lt172_c13 ),
    .o({\u2_Display/lt172_c14 ,open_n3283}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_14  (
    .a(\u2_Display/n5524 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c14 ),
    .o({\u2_Display/lt172_c15 ,open_n3284}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_15  (
    .a(\u2_Display/n5523 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c15 ),
    .o({\u2_Display/lt172_c16 ,open_n3285}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_16  (
    .a(\u2_Display/n5522 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c16 ),
    .o({\u2_Display/lt172_c17 ,open_n3286}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_17  (
    .a(\u2_Display/n5521 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c17 ),
    .o({\u2_Display/lt172_c18 ,open_n3287}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_18  (
    .a(\u2_Display/n5520 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c18 ),
    .o({\u2_Display/lt172_c19 ,open_n3288}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_19  (
    .a(\u2_Display/n5519 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c19 ),
    .o({\u2_Display/lt172_c20 ,open_n3289}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_2  (
    .a(\u2_Display/n5536 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c2 ),
    .o({\u2_Display/lt172_c3 ,open_n3290}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_20  (
    .a(\u2_Display/n5518 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c20 ),
    .o({\u2_Display/lt172_c21 ,open_n3291}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_21  (
    .a(\u2_Display/n5517 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c21 ),
    .o({\u2_Display/lt172_c22 ,open_n3292}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_22  (
    .a(\u2_Display/n5516 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c22 ),
    .o({\u2_Display/lt172_c23 ,open_n3293}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_23  (
    .a(\u2_Display/n5515 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c23 ),
    .o({\u2_Display/lt172_c24 ,open_n3294}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_24  (
    .a(\u2_Display/n5514 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c24 ),
    .o({\u2_Display/lt172_c25 ,open_n3295}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_25  (
    .a(\u2_Display/n5513 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c25 ),
    .o({\u2_Display/lt172_c26 ,open_n3296}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_26  (
    .a(\u2_Display/n5512 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c26 ),
    .o({\u2_Display/lt172_c27 ,open_n3297}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_27  (
    .a(\u2_Display/n5511 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c27 ),
    .o({\u2_Display/lt172_c28 ,open_n3298}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_28  (
    .a(\u2_Display/n5510 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c28 ),
    .o({\u2_Display/lt172_c29 ,open_n3299}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_29  (
    .a(\u2_Display/n5509 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c29 ),
    .o({\u2_Display/lt172_c30 ,open_n3300}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_3  (
    .a(\u2_Display/n5535 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c3 ),
    .o({\u2_Display/lt172_c4 ,open_n3301}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_30  (
    .a(\u2_Display/n5508 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c30 ),
    .o({\u2_Display/lt172_c31 ,open_n3302}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_31  (
    .a(\u2_Display/n5507 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c31 ),
    .o({\u2_Display/lt172_c32 ,open_n3303}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_4  (
    .a(\u2_Display/n5534 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c4 ),
    .o({\u2_Display/lt172_c5 ,open_n3304}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_5  (
    .a(\u2_Display/n5533 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c5 ),
    .o({\u2_Display/lt172_c6 ,open_n3305}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_6  (
    .a(\u2_Display/n5532 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c6 ),
    .o({\u2_Display/lt172_c7 ,open_n3306}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_7  (
    .a(\u2_Display/n5531 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c7 ),
    .o({\u2_Display/lt172_c8 ,open_n3307}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_8  (
    .a(\u2_Display/n5530 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c8 ),
    .o({\u2_Display/lt172_c9 ,open_n3308}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_9  (
    .a(\u2_Display/n5529 ),
    .b(1'b0),
    .c(\u2_Display/lt172_c9 ),
    .o({\u2_Display/lt172_c10 ,open_n3309}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt172_cin  (
    .a(1'b0),
    .o({\u2_Display/lt172_c0 ,open_n3312}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt172_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt172_c32 ),
    .o({open_n3313,\u2_Display/n5539 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_0  (
    .a(\u2_Display/n5573 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c0 ),
    .o({\u2_Display/lt173_c1 ,open_n3314}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_1  (
    .a(\u2_Display/n5572 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c1 ),
    .o({\u2_Display/lt173_c2 ,open_n3315}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_10  (
    .a(\u2_Display/n5563 ),
    .b(1'b1),
    .c(\u2_Display/lt173_c10 ),
    .o({\u2_Display/lt173_c11 ,open_n3316}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_11  (
    .a(\u2_Display/n5562 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c11 ),
    .o({\u2_Display/lt173_c12 ,open_n3317}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_12  (
    .a(\u2_Display/n5561 ),
    .b(1'b1),
    .c(\u2_Display/lt173_c12 ),
    .o({\u2_Display/lt173_c13 ,open_n3318}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_13  (
    .a(\u2_Display/n5560 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c13 ),
    .o({\u2_Display/lt173_c14 ,open_n3319}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_14  (
    .a(\u2_Display/n5559 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c14 ),
    .o({\u2_Display/lt173_c15 ,open_n3320}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_15  (
    .a(\u2_Display/n5558 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c15 ),
    .o({\u2_Display/lt173_c16 ,open_n3321}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_16  (
    .a(\u2_Display/n5557 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c16 ),
    .o({\u2_Display/lt173_c17 ,open_n3322}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_17  (
    .a(\u2_Display/n5556 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c17 ),
    .o({\u2_Display/lt173_c18 ,open_n3323}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_18  (
    .a(\u2_Display/n5555 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c18 ),
    .o({\u2_Display/lt173_c19 ,open_n3324}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_19  (
    .a(\u2_Display/n5554 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c19 ),
    .o({\u2_Display/lt173_c20 ,open_n3325}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_2  (
    .a(\u2_Display/n5571 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c2 ),
    .o({\u2_Display/lt173_c3 ,open_n3326}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_20  (
    .a(\u2_Display/n5553 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c20 ),
    .o({\u2_Display/lt173_c21 ,open_n3327}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_21  (
    .a(\u2_Display/n5552 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c21 ),
    .o({\u2_Display/lt173_c22 ,open_n3328}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_22  (
    .a(\u2_Display/n5551 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c22 ),
    .o({\u2_Display/lt173_c23 ,open_n3329}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_23  (
    .a(\u2_Display/n5550 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c23 ),
    .o({\u2_Display/lt173_c24 ,open_n3330}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_24  (
    .a(\u2_Display/n5549 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c24 ),
    .o({\u2_Display/lt173_c25 ,open_n3331}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_25  (
    .a(\u2_Display/n5548 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c25 ),
    .o({\u2_Display/lt173_c26 ,open_n3332}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_26  (
    .a(\u2_Display/n5547 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c26 ),
    .o({\u2_Display/lt173_c27 ,open_n3333}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_27  (
    .a(\u2_Display/n5546 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c27 ),
    .o({\u2_Display/lt173_c28 ,open_n3334}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_28  (
    .a(\u2_Display/n5545 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c28 ),
    .o({\u2_Display/lt173_c29 ,open_n3335}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_29  (
    .a(\u2_Display/n5544 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c29 ),
    .o({\u2_Display/lt173_c30 ,open_n3336}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_3  (
    .a(\u2_Display/n5570 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c3 ),
    .o({\u2_Display/lt173_c4 ,open_n3337}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_30  (
    .a(\u2_Display/n5543 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c30 ),
    .o({\u2_Display/lt173_c31 ,open_n3338}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_31  (
    .a(\u2_Display/n5542 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c31 ),
    .o({\u2_Display/lt173_c32 ,open_n3339}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_4  (
    .a(\u2_Display/n5569 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c4 ),
    .o({\u2_Display/lt173_c5 ,open_n3340}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_5  (
    .a(\u2_Display/n5568 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c5 ),
    .o({\u2_Display/lt173_c6 ,open_n3341}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_6  (
    .a(\u2_Display/n5567 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c6 ),
    .o({\u2_Display/lt173_c7 ,open_n3342}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_7  (
    .a(\u2_Display/n5566 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c7 ),
    .o({\u2_Display/lt173_c8 ,open_n3343}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_8  (
    .a(\u2_Display/n5565 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c8 ),
    .o({\u2_Display/lt173_c9 ,open_n3344}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_9  (
    .a(\u2_Display/n5564 ),
    .b(1'b0),
    .c(\u2_Display/lt173_c9 ),
    .o({\u2_Display/lt173_c10 ,open_n3345}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt173_cin  (
    .a(1'b0),
    .o({\u2_Display/lt173_c0 ,open_n3348}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt173_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt173_c32 ),
    .o({open_n3349,\u2_Display/n5574 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_0  (
    .a(\u2_Display/n5608 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c0 ),
    .o({\u2_Display/lt174_c1 ,open_n3350}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_1  (
    .a(\u2_Display/n5607 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c1 ),
    .o({\u2_Display/lt174_c2 ,open_n3351}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_10  (
    .a(\u2_Display/n5598 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c10 ),
    .o({\u2_Display/lt174_c11 ,open_n3352}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_11  (
    .a(\u2_Display/n5597 ),
    .b(1'b1),
    .c(\u2_Display/lt174_c11 ),
    .o({\u2_Display/lt174_c12 ,open_n3353}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_12  (
    .a(\u2_Display/n5596 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c12 ),
    .o({\u2_Display/lt174_c13 ,open_n3354}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_13  (
    .a(\u2_Display/n5595 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c13 ),
    .o({\u2_Display/lt174_c14 ,open_n3355}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_14  (
    .a(\u2_Display/n5594 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c14 ),
    .o({\u2_Display/lt174_c15 ,open_n3356}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_15  (
    .a(\u2_Display/n5593 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c15 ),
    .o({\u2_Display/lt174_c16 ,open_n3357}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_16  (
    .a(\u2_Display/n5592 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c16 ),
    .o({\u2_Display/lt174_c17 ,open_n3358}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_17  (
    .a(\u2_Display/n5591 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c17 ),
    .o({\u2_Display/lt174_c18 ,open_n3359}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_18  (
    .a(\u2_Display/n5590 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c18 ),
    .o({\u2_Display/lt174_c19 ,open_n3360}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_19  (
    .a(\u2_Display/n5589 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c19 ),
    .o({\u2_Display/lt174_c20 ,open_n3361}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_2  (
    .a(\u2_Display/n5606 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c2 ),
    .o({\u2_Display/lt174_c3 ,open_n3362}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_20  (
    .a(\u2_Display/n5588 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c20 ),
    .o({\u2_Display/lt174_c21 ,open_n3363}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_21  (
    .a(\u2_Display/n5587 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c21 ),
    .o({\u2_Display/lt174_c22 ,open_n3364}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_22  (
    .a(\u2_Display/n5586 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c22 ),
    .o({\u2_Display/lt174_c23 ,open_n3365}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_23  (
    .a(\u2_Display/n5585 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c23 ),
    .o({\u2_Display/lt174_c24 ,open_n3366}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_24  (
    .a(\u2_Display/n5584 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c24 ),
    .o({\u2_Display/lt174_c25 ,open_n3367}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_25  (
    .a(\u2_Display/n5583 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c25 ),
    .o({\u2_Display/lt174_c26 ,open_n3368}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_26  (
    .a(\u2_Display/n5582 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c26 ),
    .o({\u2_Display/lt174_c27 ,open_n3369}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_27  (
    .a(\u2_Display/n5581 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c27 ),
    .o({\u2_Display/lt174_c28 ,open_n3370}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_28  (
    .a(\u2_Display/n5580 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c28 ),
    .o({\u2_Display/lt174_c29 ,open_n3371}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_29  (
    .a(\u2_Display/n5579 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c29 ),
    .o({\u2_Display/lt174_c30 ,open_n3372}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_3  (
    .a(\u2_Display/n5605 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c3 ),
    .o({\u2_Display/lt174_c4 ,open_n3373}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_30  (
    .a(\u2_Display/n5578 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c30 ),
    .o({\u2_Display/lt174_c31 ,open_n3374}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_31  (
    .a(\u2_Display/n5577 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c31 ),
    .o({\u2_Display/lt174_c32 ,open_n3375}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_4  (
    .a(\u2_Display/n5604 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c4 ),
    .o({\u2_Display/lt174_c5 ,open_n3376}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_5  (
    .a(\u2_Display/n5603 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c5 ),
    .o({\u2_Display/lt174_c6 ,open_n3377}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_6  (
    .a(\u2_Display/n5602 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c6 ),
    .o({\u2_Display/lt174_c7 ,open_n3378}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_7  (
    .a(\u2_Display/n5601 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c7 ),
    .o({\u2_Display/lt174_c8 ,open_n3379}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_8  (
    .a(\u2_Display/n5600 ),
    .b(1'b0),
    .c(\u2_Display/lt174_c8 ),
    .o({\u2_Display/lt174_c9 ,open_n3380}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_9  (
    .a(\u2_Display/n5599 ),
    .b(1'b1),
    .c(\u2_Display/lt174_c9 ),
    .o({\u2_Display/lt174_c10 ,open_n3381}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt174_cin  (
    .a(1'b0),
    .o({\u2_Display/lt174_c0 ,open_n3384}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt174_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt174_c32 ),
    .o({open_n3385,\u2_Display/n5609 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_0  (
    .a(\u2_Display/n5643 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c0 ),
    .o({\u2_Display/lt175_c1 ,open_n3386}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_1  (
    .a(\u2_Display/n5642 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c1 ),
    .o({\u2_Display/lt175_c2 ,open_n3387}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_10  (
    .a(\u2_Display/n5633 ),
    .b(1'b1),
    .c(\u2_Display/lt175_c10 ),
    .o({\u2_Display/lt175_c11 ,open_n3388}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_11  (
    .a(\u2_Display/n5632 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c11 ),
    .o({\u2_Display/lt175_c12 ,open_n3389}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_12  (
    .a(\u2_Display/n5631 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c12 ),
    .o({\u2_Display/lt175_c13 ,open_n3390}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_13  (
    .a(\u2_Display/n5630 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c13 ),
    .o({\u2_Display/lt175_c14 ,open_n3391}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_14  (
    .a(\u2_Display/n5629 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c14 ),
    .o({\u2_Display/lt175_c15 ,open_n3392}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_15  (
    .a(\u2_Display/n5628 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c15 ),
    .o({\u2_Display/lt175_c16 ,open_n3393}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_16  (
    .a(\u2_Display/n5627 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c16 ),
    .o({\u2_Display/lt175_c17 ,open_n3394}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_17  (
    .a(\u2_Display/n5626 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c17 ),
    .o({\u2_Display/lt175_c18 ,open_n3395}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_18  (
    .a(\u2_Display/n5625 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c18 ),
    .o({\u2_Display/lt175_c19 ,open_n3396}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_19  (
    .a(\u2_Display/n5624 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c19 ),
    .o({\u2_Display/lt175_c20 ,open_n3397}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_2  (
    .a(\u2_Display/n5641 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c2 ),
    .o({\u2_Display/lt175_c3 ,open_n3398}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_20  (
    .a(\u2_Display/n5623 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c20 ),
    .o({\u2_Display/lt175_c21 ,open_n3399}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_21  (
    .a(\u2_Display/n5622 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c21 ),
    .o({\u2_Display/lt175_c22 ,open_n3400}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_22  (
    .a(\u2_Display/n5621 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c22 ),
    .o({\u2_Display/lt175_c23 ,open_n3401}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_23  (
    .a(\u2_Display/n5620 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c23 ),
    .o({\u2_Display/lt175_c24 ,open_n3402}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_24  (
    .a(\u2_Display/n5619 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c24 ),
    .o({\u2_Display/lt175_c25 ,open_n3403}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_25  (
    .a(\u2_Display/n5618 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c25 ),
    .o({\u2_Display/lt175_c26 ,open_n3404}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_26  (
    .a(\u2_Display/n5617 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c26 ),
    .o({\u2_Display/lt175_c27 ,open_n3405}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_27  (
    .a(\u2_Display/n5616 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c27 ),
    .o({\u2_Display/lt175_c28 ,open_n3406}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_28  (
    .a(\u2_Display/n5615 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c28 ),
    .o({\u2_Display/lt175_c29 ,open_n3407}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_29  (
    .a(\u2_Display/n5614 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c29 ),
    .o({\u2_Display/lt175_c30 ,open_n3408}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_3  (
    .a(\u2_Display/n5640 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c3 ),
    .o({\u2_Display/lt175_c4 ,open_n3409}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_30  (
    .a(\u2_Display/n5613 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c30 ),
    .o({\u2_Display/lt175_c31 ,open_n3410}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_31  (
    .a(\u2_Display/n5612 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c31 ),
    .o({\u2_Display/lt175_c32 ,open_n3411}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_4  (
    .a(\u2_Display/n5639 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c4 ),
    .o({\u2_Display/lt175_c5 ,open_n3412}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_5  (
    .a(\u2_Display/n5638 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c5 ),
    .o({\u2_Display/lt175_c6 ,open_n3413}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_6  (
    .a(\u2_Display/n5637 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c6 ),
    .o({\u2_Display/lt175_c7 ,open_n3414}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_7  (
    .a(\u2_Display/n5636 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c7 ),
    .o({\u2_Display/lt175_c8 ,open_n3415}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_8  (
    .a(\u2_Display/n5635 ),
    .b(1'b1),
    .c(\u2_Display/lt175_c8 ),
    .o({\u2_Display/lt175_c9 ,open_n3416}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_9  (
    .a(\u2_Display/n5634 ),
    .b(1'b0),
    .c(\u2_Display/lt175_c9 ),
    .o({\u2_Display/lt175_c10 ,open_n3417}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt175_cin  (
    .a(1'b0),
    .o({\u2_Display/lt175_c0 ,open_n3420}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt175_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt175_c32 ),
    .o({open_n3421,\u2_Display/n5644 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_0  (
    .a(\u2_Display/n5678 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c0 ),
    .o({\u2_Display/lt176_c1 ,open_n3422}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_1  (
    .a(\u2_Display/n5677 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c1 ),
    .o({\u2_Display/lt176_c2 ,open_n3423}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_10  (
    .a(\u2_Display/n5668 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c10 ),
    .o({\u2_Display/lt176_c11 ,open_n3424}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_11  (
    .a(\u2_Display/n5667 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c11 ),
    .o({\u2_Display/lt176_c12 ,open_n3425}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_12  (
    .a(\u2_Display/n5666 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c12 ),
    .o({\u2_Display/lt176_c13 ,open_n3426}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_13  (
    .a(\u2_Display/n5665 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c13 ),
    .o({\u2_Display/lt176_c14 ,open_n3427}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_14  (
    .a(\u2_Display/n5664 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c14 ),
    .o({\u2_Display/lt176_c15 ,open_n3428}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_15  (
    .a(\u2_Display/n5663 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c15 ),
    .o({\u2_Display/lt176_c16 ,open_n3429}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_16  (
    .a(\u2_Display/n5662 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c16 ),
    .o({\u2_Display/lt176_c17 ,open_n3430}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_17  (
    .a(\u2_Display/n5661 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c17 ),
    .o({\u2_Display/lt176_c18 ,open_n3431}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_18  (
    .a(\u2_Display/n5660 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c18 ),
    .o({\u2_Display/lt176_c19 ,open_n3432}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_19  (
    .a(\u2_Display/n5659 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c19 ),
    .o({\u2_Display/lt176_c20 ,open_n3433}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_2  (
    .a(\u2_Display/n5676 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c2 ),
    .o({\u2_Display/lt176_c3 ,open_n3434}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_20  (
    .a(\u2_Display/n5658 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c20 ),
    .o({\u2_Display/lt176_c21 ,open_n3435}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_21  (
    .a(\u2_Display/n5657 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c21 ),
    .o({\u2_Display/lt176_c22 ,open_n3436}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_22  (
    .a(\u2_Display/n5656 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c22 ),
    .o({\u2_Display/lt176_c23 ,open_n3437}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_23  (
    .a(\u2_Display/n5655 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c23 ),
    .o({\u2_Display/lt176_c24 ,open_n3438}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_24  (
    .a(\u2_Display/n5654 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c24 ),
    .o({\u2_Display/lt176_c25 ,open_n3439}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_25  (
    .a(\u2_Display/n5653 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c25 ),
    .o({\u2_Display/lt176_c26 ,open_n3440}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_26  (
    .a(\u2_Display/n5652 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c26 ),
    .o({\u2_Display/lt176_c27 ,open_n3441}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_27  (
    .a(\u2_Display/n5651 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c27 ),
    .o({\u2_Display/lt176_c28 ,open_n3442}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_28  (
    .a(\u2_Display/n5650 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c28 ),
    .o({\u2_Display/lt176_c29 ,open_n3443}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_29  (
    .a(\u2_Display/n5649 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c29 ),
    .o({\u2_Display/lt176_c30 ,open_n3444}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_3  (
    .a(\u2_Display/n5675 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c3 ),
    .o({\u2_Display/lt176_c4 ,open_n3445}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_30  (
    .a(\u2_Display/n5648 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c30 ),
    .o({\u2_Display/lt176_c31 ,open_n3446}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_31  (
    .a(\u2_Display/n5647 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c31 ),
    .o({\u2_Display/lt176_c32 ,open_n3447}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_4  (
    .a(\u2_Display/n5674 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c4 ),
    .o({\u2_Display/lt176_c5 ,open_n3448}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_5  (
    .a(\u2_Display/n5673 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c5 ),
    .o({\u2_Display/lt176_c6 ,open_n3449}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_6  (
    .a(\u2_Display/n5672 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c6 ),
    .o({\u2_Display/lt176_c7 ,open_n3450}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_7  (
    .a(\u2_Display/n5671 ),
    .b(1'b1),
    .c(\u2_Display/lt176_c7 ),
    .o({\u2_Display/lt176_c8 ,open_n3451}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_8  (
    .a(\u2_Display/n5670 ),
    .b(1'b0),
    .c(\u2_Display/lt176_c8 ),
    .o({\u2_Display/lt176_c9 ,open_n3452}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_9  (
    .a(\u2_Display/n5669 ),
    .b(1'b1),
    .c(\u2_Display/lt176_c9 ),
    .o({\u2_Display/lt176_c10 ,open_n3453}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt176_cin  (
    .a(1'b0),
    .o({\u2_Display/lt176_c0 ,open_n3456}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt176_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt176_c32 ),
    .o({open_n3457,\u2_Display/n5679 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt1_0  (
    .a(\u2_Display/i [0]),
    .b(lcd_xpos[0]),
    .c(\u2_Display/lt1_c0 ),
    .o({\u2_Display/lt1_c1 ,open_n3458}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt1_1  (
    .a(\u2_Display/i [1]),
    .b(lcd_xpos[1]),
    .c(\u2_Display/lt1_c1 ),
    .o({\u2_Display/lt1_c2 ,open_n3459}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt1_10  (
    .a(\u2_Display/i [10]),
    .b(lcd_xpos[10]),
    .c(\u2_Display/lt1_c10 ),
    .o({\u2_Display/lt1_c11 ,open_n3460}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt1_11  (
    .a(1'b0),
    .b(lcd_xpos[11]),
    .c(\u2_Display/lt1_c11 ),
    .o({\u2_Display/lt1_c12 ,open_n3461}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt1_2  (
    .a(\u2_Display/i [2]),
    .b(lcd_xpos[2]),
    .c(\u2_Display/lt1_c2 ),
    .o({\u2_Display/lt1_c3 ,open_n3462}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt1_3  (
    .a(\u2_Display/i [3]),
    .b(lcd_xpos[3]),
    .c(\u2_Display/lt1_c3 ),
    .o({\u2_Display/lt1_c4 ,open_n3463}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt1_4  (
    .a(\u2_Display/i [4]),
    .b(lcd_xpos[4]),
    .c(\u2_Display/lt1_c4 ),
    .o({\u2_Display/lt1_c5 ,open_n3464}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt1_5  (
    .a(\u2_Display/i [5]),
    .b(lcd_xpos[5]),
    .c(\u2_Display/lt1_c5 ),
    .o({\u2_Display/lt1_c6 ,open_n3465}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt1_6  (
    .a(\u2_Display/i [6]),
    .b(lcd_xpos[6]),
    .c(\u2_Display/lt1_c6 ),
    .o({\u2_Display/lt1_c7 ,open_n3466}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt1_7  (
    .a(\u2_Display/i [7]),
    .b(lcd_xpos[7]),
    .c(\u2_Display/lt1_c7 ),
    .o({\u2_Display/lt1_c8 ,open_n3467}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt1_8  (
    .a(\u2_Display/i [8]),
    .b(lcd_xpos[8]),
    .c(\u2_Display/lt1_c8 ),
    .o({\u2_Display/lt1_c9 ,open_n3468}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt1_9  (
    .a(\u2_Display/i [9]),
    .b(lcd_xpos[9]),
    .c(\u2_Display/lt1_c9 ),
    .o({\u2_Display/lt1_c10 ,open_n3469}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt1_cin  (
    .a(1'b0),
    .o({\u2_Display/lt1_c0 ,open_n3472}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt1_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt1_c12 ),
    .o({open_n3473,\u2_Display/n45 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_0  (
    .a(\u2_Display/counta [0]),
    .b(1'b0),
    .c(\u2_Display/lt22_c0 ),
    .o({\u2_Display/lt22_c1 ,open_n3474}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_1  (
    .a(\u2_Display/counta [1]),
    .b(1'b0),
    .c(\u2_Display/lt22_c1 ),
    .o({\u2_Display/lt22_c2 ,open_n3475}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_10  (
    .a(\u2_Display/counta [10]),
    .b(1'b0),
    .c(\u2_Display/lt22_c10 ),
    .o({\u2_Display/lt22_c11 ,open_n3476}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_11  (
    .a(\u2_Display/counta [11]),
    .b(1'b0),
    .c(\u2_Display/lt22_c11 ),
    .o({\u2_Display/lt22_c12 ,open_n3477}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_12  (
    .a(\u2_Display/counta [12]),
    .b(1'b0),
    .c(\u2_Display/lt22_c12 ),
    .o({\u2_Display/lt22_c13 ,open_n3478}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_13  (
    .a(\u2_Display/counta [13]),
    .b(1'b0),
    .c(\u2_Display/lt22_c13 ),
    .o({\u2_Display/lt22_c14 ,open_n3479}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_14  (
    .a(\u2_Display/counta [14]),
    .b(1'b0),
    .c(\u2_Display/lt22_c14 ),
    .o({\u2_Display/lt22_c15 ,open_n3480}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_15  (
    .a(\u2_Display/counta [15]),
    .b(1'b0),
    .c(\u2_Display/lt22_c15 ),
    .o({\u2_Display/lt22_c16 ,open_n3481}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_16  (
    .a(\u2_Display/counta [16]),
    .b(1'b0),
    .c(\u2_Display/lt22_c16 ),
    .o({\u2_Display/lt22_c17 ,open_n3482}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_17  (
    .a(\u2_Display/counta [17]),
    .b(1'b0),
    .c(\u2_Display/lt22_c17 ),
    .o({\u2_Display/lt22_c18 ,open_n3483}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_18  (
    .a(\u2_Display/counta [18]),
    .b(1'b0),
    .c(\u2_Display/lt22_c18 ),
    .o({\u2_Display/lt22_c19 ,open_n3484}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_19  (
    .a(\u2_Display/counta [19]),
    .b(1'b0),
    .c(\u2_Display/lt22_c19 ),
    .o({\u2_Display/lt22_c20 ,open_n3485}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_2  (
    .a(\u2_Display/counta [2]),
    .b(1'b0),
    .c(\u2_Display/lt22_c2 ),
    .o({\u2_Display/lt22_c3 ,open_n3486}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_20  (
    .a(\u2_Display/counta [20]),
    .b(1'b0),
    .c(\u2_Display/lt22_c20 ),
    .o({\u2_Display/lt22_c21 ,open_n3487}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_21  (
    .a(\u2_Display/counta [21]),
    .b(1'b0),
    .c(\u2_Display/lt22_c21 ),
    .o({\u2_Display/lt22_c22 ,open_n3488}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_22  (
    .a(\u2_Display/counta [22]),
    .b(1'b0),
    .c(\u2_Display/lt22_c22 ),
    .o({\u2_Display/lt22_c23 ,open_n3489}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_23  (
    .a(\u2_Display/counta [23]),
    .b(1'b0),
    .c(\u2_Display/lt22_c23 ),
    .o({\u2_Display/lt22_c24 ,open_n3490}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_24  (
    .a(\u2_Display/counta [24]),
    .b(1'b0),
    .c(\u2_Display/lt22_c24 ),
    .o({\u2_Display/lt22_c25 ,open_n3491}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_25  (
    .a(\u2_Display/counta [25]),
    .b(1'b1),
    .c(\u2_Display/lt22_c25 ),
    .o({\u2_Display/lt22_c26 ,open_n3492}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_26  (
    .a(\u2_Display/counta [26]),
    .b(1'b0),
    .c(\u2_Display/lt22_c26 ),
    .o({\u2_Display/lt22_c27 ,open_n3493}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_27  (
    .a(\u2_Display/counta [27]),
    .b(1'b1),
    .c(\u2_Display/lt22_c27 ),
    .o({\u2_Display/lt22_c28 ,open_n3494}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_28  (
    .a(\u2_Display/counta [28]),
    .b(1'b1),
    .c(\u2_Display/lt22_c28 ),
    .o({\u2_Display/lt22_c29 ,open_n3495}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_29  (
    .a(\u2_Display/counta [29]),
    .b(1'b1),
    .c(\u2_Display/lt22_c29 ),
    .o({\u2_Display/lt22_c30 ,open_n3496}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_3  (
    .a(\u2_Display/counta [3]),
    .b(1'b0),
    .c(\u2_Display/lt22_c3 ),
    .o({\u2_Display/lt22_c4 ,open_n3497}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_30  (
    .a(\u2_Display/counta [30]),
    .b(1'b1),
    .c(\u2_Display/lt22_c30 ),
    .o({\u2_Display/lt22_c31 ,open_n3498}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_31  (
    .a(\u2_Display/counta [31]),
    .b(1'b1),
    .c(\u2_Display/lt22_c31 ),
    .o({\u2_Display/lt22_c32 ,open_n3499}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_4  (
    .a(\u2_Display/counta [4]),
    .b(1'b0),
    .c(\u2_Display/lt22_c4 ),
    .o({\u2_Display/lt22_c5 ,open_n3500}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_5  (
    .a(\u2_Display/counta [5]),
    .b(1'b0),
    .c(\u2_Display/lt22_c5 ),
    .o({\u2_Display/lt22_c6 ,open_n3501}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_6  (
    .a(\u2_Display/counta [6]),
    .b(1'b0),
    .c(\u2_Display/lt22_c6 ),
    .o({\u2_Display/lt22_c7 ,open_n3502}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_7  (
    .a(\u2_Display/counta [7]),
    .b(1'b0),
    .c(\u2_Display/lt22_c7 ),
    .o({\u2_Display/lt22_c8 ,open_n3503}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_8  (
    .a(\u2_Display/counta [8]),
    .b(1'b0),
    .c(\u2_Display/lt22_c8 ),
    .o({\u2_Display/lt22_c9 ,open_n3504}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_9  (
    .a(\u2_Display/counta [9]),
    .b(1'b0),
    .c(\u2_Display/lt22_c9 ),
    .o({\u2_Display/lt22_c10 ,open_n3505}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt22_cin  (
    .a(1'b0),
    .o({\u2_Display/lt22_c0 ,open_n3508}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt22_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt22_c32 ),
    .o({open_n3509,\u2_Display/n417 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_0  (
    .a(\u2_Display/n451 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c0 ),
    .o({\u2_Display/lt23_c1 ,open_n3510}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_1  (
    .a(\u2_Display/n450 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c1 ),
    .o({\u2_Display/lt23_c2 ,open_n3511}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_10  (
    .a(\u2_Display/n441 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c10 ),
    .o({\u2_Display/lt23_c11 ,open_n3512}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_11  (
    .a(\u2_Display/n440 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c11 ),
    .o({\u2_Display/lt23_c12 ,open_n3513}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_12  (
    .a(\u2_Display/n439 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c12 ),
    .o({\u2_Display/lt23_c13 ,open_n3514}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_13  (
    .a(\u2_Display/n438 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c13 ),
    .o({\u2_Display/lt23_c14 ,open_n3515}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_14  (
    .a(\u2_Display/n437 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c14 ),
    .o({\u2_Display/lt23_c15 ,open_n3516}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_15  (
    .a(\u2_Display/n436 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c15 ),
    .o({\u2_Display/lt23_c16 ,open_n3517}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_16  (
    .a(\u2_Display/n435 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c16 ),
    .o({\u2_Display/lt23_c17 ,open_n3518}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_17  (
    .a(\u2_Display/n434 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c17 ),
    .o({\u2_Display/lt23_c18 ,open_n3519}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_18  (
    .a(\u2_Display/n433 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c18 ),
    .o({\u2_Display/lt23_c19 ,open_n3520}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_19  (
    .a(\u2_Display/n432 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c19 ),
    .o({\u2_Display/lt23_c20 ,open_n3521}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_2  (
    .a(\u2_Display/n449 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c2 ),
    .o({\u2_Display/lt23_c3 ,open_n3522}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_20  (
    .a(\u2_Display/n431 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c20 ),
    .o({\u2_Display/lt23_c21 ,open_n3523}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_21  (
    .a(\u2_Display/n430 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c21 ),
    .o({\u2_Display/lt23_c22 ,open_n3524}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_22  (
    .a(\u2_Display/n429 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c22 ),
    .o({\u2_Display/lt23_c23 ,open_n3525}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_23  (
    .a(\u2_Display/n428 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c23 ),
    .o({\u2_Display/lt23_c24 ,open_n3526}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_24  (
    .a(\u2_Display/n427 ),
    .b(1'b1),
    .c(\u2_Display/lt23_c24 ),
    .o({\u2_Display/lt23_c25 ,open_n3527}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_25  (
    .a(\u2_Display/n426 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c25 ),
    .o({\u2_Display/lt23_c26 ,open_n3528}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_26  (
    .a(\u2_Display/n425 ),
    .b(1'b1),
    .c(\u2_Display/lt23_c26 ),
    .o({\u2_Display/lt23_c27 ,open_n3529}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_27  (
    .a(\u2_Display/n424 ),
    .b(1'b1),
    .c(\u2_Display/lt23_c27 ),
    .o({\u2_Display/lt23_c28 ,open_n3530}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_28  (
    .a(\u2_Display/n423 ),
    .b(1'b1),
    .c(\u2_Display/lt23_c28 ),
    .o({\u2_Display/lt23_c29 ,open_n3531}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_29  (
    .a(\u2_Display/n422 ),
    .b(1'b1),
    .c(\u2_Display/lt23_c29 ),
    .o({\u2_Display/lt23_c30 ,open_n3532}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_3  (
    .a(\u2_Display/n448 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c3 ),
    .o({\u2_Display/lt23_c4 ,open_n3533}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_30  (
    .a(\u2_Display/n421 ),
    .b(1'b1),
    .c(\u2_Display/lt23_c30 ),
    .o({\u2_Display/lt23_c31 ,open_n3534}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_31  (
    .a(\u2_Display/n420 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c31 ),
    .o({\u2_Display/lt23_c32 ,open_n3535}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_4  (
    .a(\u2_Display/n447 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c4 ),
    .o({\u2_Display/lt23_c5 ,open_n3536}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_5  (
    .a(\u2_Display/n446 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c5 ),
    .o({\u2_Display/lt23_c6 ,open_n3537}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_6  (
    .a(\u2_Display/n445 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c6 ),
    .o({\u2_Display/lt23_c7 ,open_n3538}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_7  (
    .a(\u2_Display/n444 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c7 ),
    .o({\u2_Display/lt23_c8 ,open_n3539}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_8  (
    .a(\u2_Display/n443 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c8 ),
    .o({\u2_Display/lt23_c9 ,open_n3540}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_9  (
    .a(\u2_Display/n442 ),
    .b(1'b0),
    .c(\u2_Display/lt23_c9 ),
    .o({\u2_Display/lt23_c10 ,open_n3541}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt23_cin  (
    .a(1'b0),
    .o({\u2_Display/lt23_c0 ,open_n3544}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt23_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt23_c32 ),
    .o({open_n3545,\u2_Display/n452 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_0  (
    .a(\u2_Display/n486 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c0 ),
    .o({\u2_Display/lt24_c1 ,open_n3546}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_1  (
    .a(\u2_Display/n485 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c1 ),
    .o({\u2_Display/lt24_c2 ,open_n3547}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_10  (
    .a(\u2_Display/n476 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c10 ),
    .o({\u2_Display/lt24_c11 ,open_n3548}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_11  (
    .a(\u2_Display/n475 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c11 ),
    .o({\u2_Display/lt24_c12 ,open_n3549}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_12  (
    .a(\u2_Display/n474 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c12 ),
    .o({\u2_Display/lt24_c13 ,open_n3550}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_13  (
    .a(\u2_Display/n473 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c13 ),
    .o({\u2_Display/lt24_c14 ,open_n3551}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_14  (
    .a(\u2_Display/n472 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c14 ),
    .o({\u2_Display/lt24_c15 ,open_n3552}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_15  (
    .a(\u2_Display/n471 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c15 ),
    .o({\u2_Display/lt24_c16 ,open_n3553}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_16  (
    .a(\u2_Display/n470 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c16 ),
    .o({\u2_Display/lt24_c17 ,open_n3554}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_17  (
    .a(\u2_Display/n469 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c17 ),
    .o({\u2_Display/lt24_c18 ,open_n3555}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_18  (
    .a(\u2_Display/n468 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c18 ),
    .o({\u2_Display/lt24_c19 ,open_n3556}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_19  (
    .a(\u2_Display/n467 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c19 ),
    .o({\u2_Display/lt24_c20 ,open_n3557}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_2  (
    .a(\u2_Display/n484 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c2 ),
    .o({\u2_Display/lt24_c3 ,open_n3558}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_20  (
    .a(\u2_Display/n466 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c20 ),
    .o({\u2_Display/lt24_c21 ,open_n3559}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_21  (
    .a(\u2_Display/n465 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c21 ),
    .o({\u2_Display/lt24_c22 ,open_n3560}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_22  (
    .a(\u2_Display/n464 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c22 ),
    .o({\u2_Display/lt24_c23 ,open_n3561}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_23  (
    .a(\u2_Display/n463 ),
    .b(1'b1),
    .c(\u2_Display/lt24_c23 ),
    .o({\u2_Display/lt24_c24 ,open_n3562}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_24  (
    .a(\u2_Display/n462 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c24 ),
    .o({\u2_Display/lt24_c25 ,open_n3563}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_25  (
    .a(\u2_Display/n461 ),
    .b(1'b1),
    .c(\u2_Display/lt24_c25 ),
    .o({\u2_Display/lt24_c26 ,open_n3564}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_26  (
    .a(\u2_Display/n460 ),
    .b(1'b1),
    .c(\u2_Display/lt24_c26 ),
    .o({\u2_Display/lt24_c27 ,open_n3565}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_27  (
    .a(\u2_Display/n459 ),
    .b(1'b1),
    .c(\u2_Display/lt24_c27 ),
    .o({\u2_Display/lt24_c28 ,open_n3566}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_28  (
    .a(\u2_Display/n458 ),
    .b(1'b1),
    .c(\u2_Display/lt24_c28 ),
    .o({\u2_Display/lt24_c29 ,open_n3567}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_29  (
    .a(\u2_Display/n457 ),
    .b(1'b1),
    .c(\u2_Display/lt24_c29 ),
    .o({\u2_Display/lt24_c30 ,open_n3568}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_3  (
    .a(\u2_Display/n483 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c3 ),
    .o({\u2_Display/lt24_c4 ,open_n3569}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_30  (
    .a(\u2_Display/n456 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c30 ),
    .o({\u2_Display/lt24_c31 ,open_n3570}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_31  (
    .a(\u2_Display/n455 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c31 ),
    .o({\u2_Display/lt24_c32 ,open_n3571}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_4  (
    .a(\u2_Display/n482 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c4 ),
    .o({\u2_Display/lt24_c5 ,open_n3572}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_5  (
    .a(\u2_Display/n481 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c5 ),
    .o({\u2_Display/lt24_c6 ,open_n3573}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_6  (
    .a(\u2_Display/n480 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c6 ),
    .o({\u2_Display/lt24_c7 ,open_n3574}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_7  (
    .a(\u2_Display/n479 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c7 ),
    .o({\u2_Display/lt24_c8 ,open_n3575}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_8  (
    .a(\u2_Display/n478 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c8 ),
    .o({\u2_Display/lt24_c9 ,open_n3576}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_9  (
    .a(\u2_Display/n477 ),
    .b(1'b0),
    .c(\u2_Display/lt24_c9 ),
    .o({\u2_Display/lt24_c10 ,open_n3577}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt24_cin  (
    .a(1'b0),
    .o({\u2_Display/lt24_c0 ,open_n3580}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt24_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt24_c32 ),
    .o({open_n3581,\u2_Display/n487 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_0  (
    .a(\u2_Display/n521 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c0 ),
    .o({\u2_Display/lt25_c1 ,open_n3582}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_1  (
    .a(\u2_Display/n520 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c1 ),
    .o({\u2_Display/lt25_c2 ,open_n3583}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_10  (
    .a(\u2_Display/n511 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c10 ),
    .o({\u2_Display/lt25_c11 ,open_n3584}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_11  (
    .a(\u2_Display/n510 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c11 ),
    .o({\u2_Display/lt25_c12 ,open_n3585}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_12  (
    .a(\u2_Display/n509 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c12 ),
    .o({\u2_Display/lt25_c13 ,open_n3586}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_13  (
    .a(\u2_Display/n508 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c13 ),
    .o({\u2_Display/lt25_c14 ,open_n3587}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_14  (
    .a(\u2_Display/n507 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c14 ),
    .o({\u2_Display/lt25_c15 ,open_n3588}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_15  (
    .a(\u2_Display/n506 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c15 ),
    .o({\u2_Display/lt25_c16 ,open_n3589}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_16  (
    .a(\u2_Display/n505 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c16 ),
    .o({\u2_Display/lt25_c17 ,open_n3590}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_17  (
    .a(\u2_Display/n504 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c17 ),
    .o({\u2_Display/lt25_c18 ,open_n3591}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_18  (
    .a(\u2_Display/n503 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c18 ),
    .o({\u2_Display/lt25_c19 ,open_n3592}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_19  (
    .a(\u2_Display/n502 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c19 ),
    .o({\u2_Display/lt25_c20 ,open_n3593}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_2  (
    .a(\u2_Display/n519 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c2 ),
    .o({\u2_Display/lt25_c3 ,open_n3594}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_20  (
    .a(\u2_Display/n501 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c20 ),
    .o({\u2_Display/lt25_c21 ,open_n3595}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_21  (
    .a(\u2_Display/n500 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c21 ),
    .o({\u2_Display/lt25_c22 ,open_n3596}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_22  (
    .a(\u2_Display/n499 ),
    .b(1'b1),
    .c(\u2_Display/lt25_c22 ),
    .o({\u2_Display/lt25_c23 ,open_n3597}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_23  (
    .a(\u2_Display/n498 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c23 ),
    .o({\u2_Display/lt25_c24 ,open_n3598}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_24  (
    .a(\u2_Display/n497 ),
    .b(1'b1),
    .c(\u2_Display/lt25_c24 ),
    .o({\u2_Display/lt25_c25 ,open_n3599}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_25  (
    .a(\u2_Display/n496 ),
    .b(1'b1),
    .c(\u2_Display/lt25_c25 ),
    .o({\u2_Display/lt25_c26 ,open_n3600}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_26  (
    .a(\u2_Display/n495 ),
    .b(1'b1),
    .c(\u2_Display/lt25_c26 ),
    .o({\u2_Display/lt25_c27 ,open_n3601}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_27  (
    .a(\u2_Display/n494 ),
    .b(1'b1),
    .c(\u2_Display/lt25_c27 ),
    .o({\u2_Display/lt25_c28 ,open_n3602}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_28  (
    .a(\u2_Display/n493 ),
    .b(1'b1),
    .c(\u2_Display/lt25_c28 ),
    .o({\u2_Display/lt25_c29 ,open_n3603}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_29  (
    .a(\u2_Display/n492 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c29 ),
    .o({\u2_Display/lt25_c30 ,open_n3604}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_3  (
    .a(\u2_Display/n518 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c3 ),
    .o({\u2_Display/lt25_c4 ,open_n3605}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_30  (
    .a(\u2_Display/n491 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c30 ),
    .o({\u2_Display/lt25_c31 ,open_n3606}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_31  (
    .a(\u2_Display/n490 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c31 ),
    .o({\u2_Display/lt25_c32 ,open_n3607}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_4  (
    .a(\u2_Display/n517 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c4 ),
    .o({\u2_Display/lt25_c5 ,open_n3608}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_5  (
    .a(\u2_Display/n516 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c5 ),
    .o({\u2_Display/lt25_c6 ,open_n3609}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_6  (
    .a(\u2_Display/n515 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c6 ),
    .o({\u2_Display/lt25_c7 ,open_n3610}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_7  (
    .a(\u2_Display/n514 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c7 ),
    .o({\u2_Display/lt25_c8 ,open_n3611}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_8  (
    .a(\u2_Display/n513 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c8 ),
    .o({\u2_Display/lt25_c9 ,open_n3612}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_9  (
    .a(\u2_Display/n512 ),
    .b(1'b0),
    .c(\u2_Display/lt25_c9 ),
    .o({\u2_Display/lt25_c10 ,open_n3613}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt25_cin  (
    .a(1'b0),
    .o({\u2_Display/lt25_c0 ,open_n3616}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt25_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt25_c32 ),
    .o({open_n3617,\u2_Display/n522 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_0  (
    .a(\u2_Display/n556 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c0 ),
    .o({\u2_Display/lt26_c1 ,open_n3618}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_1  (
    .a(\u2_Display/n555 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c1 ),
    .o({\u2_Display/lt26_c2 ,open_n3619}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_10  (
    .a(\u2_Display/n546 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c10 ),
    .o({\u2_Display/lt26_c11 ,open_n3620}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_11  (
    .a(\u2_Display/n545 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c11 ),
    .o({\u2_Display/lt26_c12 ,open_n3621}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_12  (
    .a(\u2_Display/n544 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c12 ),
    .o({\u2_Display/lt26_c13 ,open_n3622}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_13  (
    .a(\u2_Display/n543 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c13 ),
    .o({\u2_Display/lt26_c14 ,open_n3623}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_14  (
    .a(\u2_Display/n542 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c14 ),
    .o({\u2_Display/lt26_c15 ,open_n3624}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_15  (
    .a(\u2_Display/n541 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c15 ),
    .o({\u2_Display/lt26_c16 ,open_n3625}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_16  (
    .a(\u2_Display/n540 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c16 ),
    .o({\u2_Display/lt26_c17 ,open_n3626}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_17  (
    .a(\u2_Display/n539 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c17 ),
    .o({\u2_Display/lt26_c18 ,open_n3627}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_18  (
    .a(\u2_Display/n538 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c18 ),
    .o({\u2_Display/lt26_c19 ,open_n3628}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_19  (
    .a(\u2_Display/n537 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c19 ),
    .o({\u2_Display/lt26_c20 ,open_n3629}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_2  (
    .a(\u2_Display/n554 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c2 ),
    .o({\u2_Display/lt26_c3 ,open_n3630}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_20  (
    .a(\u2_Display/n536 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c20 ),
    .o({\u2_Display/lt26_c21 ,open_n3631}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_21  (
    .a(\u2_Display/n535 ),
    .b(1'b1),
    .c(\u2_Display/lt26_c21 ),
    .o({\u2_Display/lt26_c22 ,open_n3632}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_22  (
    .a(\u2_Display/n534 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c22 ),
    .o({\u2_Display/lt26_c23 ,open_n3633}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_23  (
    .a(\u2_Display/n533 ),
    .b(1'b1),
    .c(\u2_Display/lt26_c23 ),
    .o({\u2_Display/lt26_c24 ,open_n3634}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_24  (
    .a(\u2_Display/n532 ),
    .b(1'b1),
    .c(\u2_Display/lt26_c24 ),
    .o({\u2_Display/lt26_c25 ,open_n3635}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_25  (
    .a(\u2_Display/n531 ),
    .b(1'b1),
    .c(\u2_Display/lt26_c25 ),
    .o({\u2_Display/lt26_c26 ,open_n3636}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_26  (
    .a(\u2_Display/n530 ),
    .b(1'b1),
    .c(\u2_Display/lt26_c26 ),
    .o({\u2_Display/lt26_c27 ,open_n3637}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_27  (
    .a(\u2_Display/n529 ),
    .b(1'b1),
    .c(\u2_Display/lt26_c27 ),
    .o({\u2_Display/lt26_c28 ,open_n3638}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_28  (
    .a(\u2_Display/n528 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c28 ),
    .o({\u2_Display/lt26_c29 ,open_n3639}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_29  (
    .a(\u2_Display/n527 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c29 ),
    .o({\u2_Display/lt26_c30 ,open_n3640}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_3  (
    .a(\u2_Display/n553 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c3 ),
    .o({\u2_Display/lt26_c4 ,open_n3641}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_30  (
    .a(\u2_Display/n526 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c30 ),
    .o({\u2_Display/lt26_c31 ,open_n3642}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_31  (
    .a(\u2_Display/n525 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c31 ),
    .o({\u2_Display/lt26_c32 ,open_n3643}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_4  (
    .a(\u2_Display/n552 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c4 ),
    .o({\u2_Display/lt26_c5 ,open_n3644}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_5  (
    .a(\u2_Display/n551 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c5 ),
    .o({\u2_Display/lt26_c6 ,open_n3645}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_6  (
    .a(\u2_Display/n550 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c6 ),
    .o({\u2_Display/lt26_c7 ,open_n3646}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_7  (
    .a(\u2_Display/n549 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c7 ),
    .o({\u2_Display/lt26_c8 ,open_n3647}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_8  (
    .a(\u2_Display/n548 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c8 ),
    .o({\u2_Display/lt26_c9 ,open_n3648}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_9  (
    .a(\u2_Display/n547 ),
    .b(1'b0),
    .c(\u2_Display/lt26_c9 ),
    .o({\u2_Display/lt26_c10 ,open_n3649}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt26_cin  (
    .a(1'b0),
    .o({\u2_Display/lt26_c0 ,open_n3652}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt26_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt26_c32 ),
    .o({open_n3653,\u2_Display/n557 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_0  (
    .a(\u2_Display/n591 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c0 ),
    .o({\u2_Display/lt27_c1 ,open_n3654}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_1  (
    .a(\u2_Display/n590 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c1 ),
    .o({\u2_Display/lt27_c2 ,open_n3655}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_10  (
    .a(\u2_Display/n581 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c10 ),
    .o({\u2_Display/lt27_c11 ,open_n3656}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_11  (
    .a(\u2_Display/n580 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c11 ),
    .o({\u2_Display/lt27_c12 ,open_n3657}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_12  (
    .a(\u2_Display/n579 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c12 ),
    .o({\u2_Display/lt27_c13 ,open_n3658}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_13  (
    .a(\u2_Display/n578 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c13 ),
    .o({\u2_Display/lt27_c14 ,open_n3659}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_14  (
    .a(\u2_Display/n577 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c14 ),
    .o({\u2_Display/lt27_c15 ,open_n3660}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_15  (
    .a(\u2_Display/n576 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c15 ),
    .o({\u2_Display/lt27_c16 ,open_n3661}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_16  (
    .a(\u2_Display/n575 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c16 ),
    .o({\u2_Display/lt27_c17 ,open_n3662}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_17  (
    .a(\u2_Display/n574 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c17 ),
    .o({\u2_Display/lt27_c18 ,open_n3663}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_18  (
    .a(\u2_Display/n573 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c18 ),
    .o({\u2_Display/lt27_c19 ,open_n3664}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_19  (
    .a(\u2_Display/n572 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c19 ),
    .o({\u2_Display/lt27_c20 ,open_n3665}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_2  (
    .a(\u2_Display/n589 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c2 ),
    .o({\u2_Display/lt27_c3 ,open_n3666}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_20  (
    .a(\u2_Display/n571 ),
    .b(1'b1),
    .c(\u2_Display/lt27_c20 ),
    .o({\u2_Display/lt27_c21 ,open_n3667}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_21  (
    .a(\u2_Display/n570 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c21 ),
    .o({\u2_Display/lt27_c22 ,open_n3668}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_22  (
    .a(\u2_Display/n569 ),
    .b(1'b1),
    .c(\u2_Display/lt27_c22 ),
    .o({\u2_Display/lt27_c23 ,open_n3669}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_23  (
    .a(\u2_Display/n568 ),
    .b(1'b1),
    .c(\u2_Display/lt27_c23 ),
    .o({\u2_Display/lt27_c24 ,open_n3670}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_24  (
    .a(\u2_Display/n567 ),
    .b(1'b1),
    .c(\u2_Display/lt27_c24 ),
    .o({\u2_Display/lt27_c25 ,open_n3671}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_25  (
    .a(\u2_Display/n566 ),
    .b(1'b1),
    .c(\u2_Display/lt27_c25 ),
    .o({\u2_Display/lt27_c26 ,open_n3672}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_26  (
    .a(\u2_Display/n565 ),
    .b(1'b1),
    .c(\u2_Display/lt27_c26 ),
    .o({\u2_Display/lt27_c27 ,open_n3673}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_27  (
    .a(\u2_Display/n564 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c27 ),
    .o({\u2_Display/lt27_c28 ,open_n3674}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_28  (
    .a(\u2_Display/n563 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c28 ),
    .o({\u2_Display/lt27_c29 ,open_n3675}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_29  (
    .a(\u2_Display/n562 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c29 ),
    .o({\u2_Display/lt27_c30 ,open_n3676}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_3  (
    .a(\u2_Display/n588 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c3 ),
    .o({\u2_Display/lt27_c4 ,open_n3677}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_30  (
    .a(\u2_Display/n561 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c30 ),
    .o({\u2_Display/lt27_c31 ,open_n3678}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_31  (
    .a(\u2_Display/n560 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c31 ),
    .o({\u2_Display/lt27_c32 ,open_n3679}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_4  (
    .a(\u2_Display/n587 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c4 ),
    .o({\u2_Display/lt27_c5 ,open_n3680}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_5  (
    .a(\u2_Display/n586 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c5 ),
    .o({\u2_Display/lt27_c6 ,open_n3681}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_6  (
    .a(\u2_Display/n585 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c6 ),
    .o({\u2_Display/lt27_c7 ,open_n3682}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_7  (
    .a(\u2_Display/n584 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c7 ),
    .o({\u2_Display/lt27_c8 ,open_n3683}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_8  (
    .a(\u2_Display/n583 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c8 ),
    .o({\u2_Display/lt27_c9 ,open_n3684}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_9  (
    .a(\u2_Display/n582 ),
    .b(1'b0),
    .c(\u2_Display/lt27_c9 ),
    .o({\u2_Display/lt27_c10 ,open_n3685}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt27_cin  (
    .a(1'b0),
    .o({\u2_Display/lt27_c0 ,open_n3688}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt27_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt27_c32 ),
    .o({open_n3689,\u2_Display/n592 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_0  (
    .a(\u2_Display/n626 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c0 ),
    .o({\u2_Display/lt28_c1 ,open_n3690}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_1  (
    .a(\u2_Display/n625 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c1 ),
    .o({\u2_Display/lt28_c2 ,open_n3691}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_10  (
    .a(\u2_Display/n616 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c10 ),
    .o({\u2_Display/lt28_c11 ,open_n3692}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_11  (
    .a(\u2_Display/n615 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c11 ),
    .o({\u2_Display/lt28_c12 ,open_n3693}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_12  (
    .a(\u2_Display/n614 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c12 ),
    .o({\u2_Display/lt28_c13 ,open_n3694}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_13  (
    .a(\u2_Display/n613 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c13 ),
    .o({\u2_Display/lt28_c14 ,open_n3695}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_14  (
    .a(\u2_Display/n612 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c14 ),
    .o({\u2_Display/lt28_c15 ,open_n3696}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_15  (
    .a(\u2_Display/n611 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c15 ),
    .o({\u2_Display/lt28_c16 ,open_n3697}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_16  (
    .a(\u2_Display/n610 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c16 ),
    .o({\u2_Display/lt28_c17 ,open_n3698}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_17  (
    .a(\u2_Display/n609 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c17 ),
    .o({\u2_Display/lt28_c18 ,open_n3699}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_18  (
    .a(\u2_Display/n608 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c18 ),
    .o({\u2_Display/lt28_c19 ,open_n3700}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_19  (
    .a(\u2_Display/n607 ),
    .b(1'b1),
    .c(\u2_Display/lt28_c19 ),
    .o({\u2_Display/lt28_c20 ,open_n3701}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_2  (
    .a(\u2_Display/n624 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c2 ),
    .o({\u2_Display/lt28_c3 ,open_n3702}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_20  (
    .a(\u2_Display/n606 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c20 ),
    .o({\u2_Display/lt28_c21 ,open_n3703}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_21  (
    .a(\u2_Display/n605 ),
    .b(1'b1),
    .c(\u2_Display/lt28_c21 ),
    .o({\u2_Display/lt28_c22 ,open_n3704}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_22  (
    .a(\u2_Display/n604 ),
    .b(1'b1),
    .c(\u2_Display/lt28_c22 ),
    .o({\u2_Display/lt28_c23 ,open_n3705}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_23  (
    .a(\u2_Display/n603 ),
    .b(1'b1),
    .c(\u2_Display/lt28_c23 ),
    .o({\u2_Display/lt28_c24 ,open_n3706}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_24  (
    .a(\u2_Display/n602 ),
    .b(1'b1),
    .c(\u2_Display/lt28_c24 ),
    .o({\u2_Display/lt28_c25 ,open_n3707}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_25  (
    .a(\u2_Display/n601 ),
    .b(1'b1),
    .c(\u2_Display/lt28_c25 ),
    .o({\u2_Display/lt28_c26 ,open_n3708}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_26  (
    .a(\u2_Display/n600 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c26 ),
    .o({\u2_Display/lt28_c27 ,open_n3709}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_27  (
    .a(\u2_Display/n599 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c27 ),
    .o({\u2_Display/lt28_c28 ,open_n3710}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_28  (
    .a(\u2_Display/n598 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c28 ),
    .o({\u2_Display/lt28_c29 ,open_n3711}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_29  (
    .a(\u2_Display/n597 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c29 ),
    .o({\u2_Display/lt28_c30 ,open_n3712}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_3  (
    .a(\u2_Display/n623 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c3 ),
    .o({\u2_Display/lt28_c4 ,open_n3713}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_30  (
    .a(\u2_Display/n596 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c30 ),
    .o({\u2_Display/lt28_c31 ,open_n3714}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_31  (
    .a(\u2_Display/n595 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c31 ),
    .o({\u2_Display/lt28_c32 ,open_n3715}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_4  (
    .a(\u2_Display/n622 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c4 ),
    .o({\u2_Display/lt28_c5 ,open_n3716}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_5  (
    .a(\u2_Display/n621 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c5 ),
    .o({\u2_Display/lt28_c6 ,open_n3717}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_6  (
    .a(\u2_Display/n620 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c6 ),
    .o({\u2_Display/lt28_c7 ,open_n3718}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_7  (
    .a(\u2_Display/n619 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c7 ),
    .o({\u2_Display/lt28_c8 ,open_n3719}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_8  (
    .a(\u2_Display/n618 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c8 ),
    .o({\u2_Display/lt28_c9 ,open_n3720}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_9  (
    .a(\u2_Display/n617 ),
    .b(1'b0),
    .c(\u2_Display/lt28_c9 ),
    .o({\u2_Display/lt28_c10 ,open_n3721}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt28_cin  (
    .a(1'b0),
    .o({\u2_Display/lt28_c0 ,open_n3724}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt28_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt28_c32 ),
    .o({open_n3725,\u2_Display/n627 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_0  (
    .a(\u2_Display/n661 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c0 ),
    .o({\u2_Display/lt29_c1 ,open_n3726}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_1  (
    .a(\u2_Display/n660 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c1 ),
    .o({\u2_Display/lt29_c2 ,open_n3727}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_10  (
    .a(\u2_Display/n651 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c10 ),
    .o({\u2_Display/lt29_c11 ,open_n3728}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_11  (
    .a(\u2_Display/n650 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c11 ),
    .o({\u2_Display/lt29_c12 ,open_n3729}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_12  (
    .a(\u2_Display/n649 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c12 ),
    .o({\u2_Display/lt29_c13 ,open_n3730}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_13  (
    .a(\u2_Display/n648 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c13 ),
    .o({\u2_Display/lt29_c14 ,open_n3731}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_14  (
    .a(\u2_Display/n647 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c14 ),
    .o({\u2_Display/lt29_c15 ,open_n3732}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_15  (
    .a(\u2_Display/n646 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c15 ),
    .o({\u2_Display/lt29_c16 ,open_n3733}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_16  (
    .a(\u2_Display/n645 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c16 ),
    .o({\u2_Display/lt29_c17 ,open_n3734}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_17  (
    .a(\u2_Display/n644 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c17 ),
    .o({\u2_Display/lt29_c18 ,open_n3735}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_18  (
    .a(\u2_Display/n643 ),
    .b(1'b1),
    .c(\u2_Display/lt29_c18 ),
    .o({\u2_Display/lt29_c19 ,open_n3736}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_19  (
    .a(\u2_Display/n642 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c19 ),
    .o({\u2_Display/lt29_c20 ,open_n3737}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_2  (
    .a(\u2_Display/n659 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c2 ),
    .o({\u2_Display/lt29_c3 ,open_n3738}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_20  (
    .a(\u2_Display/n641 ),
    .b(1'b1),
    .c(\u2_Display/lt29_c20 ),
    .o({\u2_Display/lt29_c21 ,open_n3739}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_21  (
    .a(\u2_Display/n640 ),
    .b(1'b1),
    .c(\u2_Display/lt29_c21 ),
    .o({\u2_Display/lt29_c22 ,open_n3740}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_22  (
    .a(\u2_Display/n639 ),
    .b(1'b1),
    .c(\u2_Display/lt29_c22 ),
    .o({\u2_Display/lt29_c23 ,open_n3741}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_23  (
    .a(\u2_Display/n638 ),
    .b(1'b1),
    .c(\u2_Display/lt29_c23 ),
    .o({\u2_Display/lt29_c24 ,open_n3742}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_24  (
    .a(\u2_Display/n637 ),
    .b(1'b1),
    .c(\u2_Display/lt29_c24 ),
    .o({\u2_Display/lt29_c25 ,open_n3743}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_25  (
    .a(\u2_Display/n636 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c25 ),
    .o({\u2_Display/lt29_c26 ,open_n3744}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_26  (
    .a(\u2_Display/n635 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c26 ),
    .o({\u2_Display/lt29_c27 ,open_n3745}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_27  (
    .a(\u2_Display/n634 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c27 ),
    .o({\u2_Display/lt29_c28 ,open_n3746}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_28  (
    .a(\u2_Display/n633 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c28 ),
    .o({\u2_Display/lt29_c29 ,open_n3747}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_29  (
    .a(\u2_Display/n632 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c29 ),
    .o({\u2_Display/lt29_c30 ,open_n3748}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_3  (
    .a(\u2_Display/n658 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c3 ),
    .o({\u2_Display/lt29_c4 ,open_n3749}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_30  (
    .a(\u2_Display/n631 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c30 ),
    .o({\u2_Display/lt29_c31 ,open_n3750}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_31  (
    .a(\u2_Display/n630 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c31 ),
    .o({\u2_Display/lt29_c32 ,open_n3751}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_4  (
    .a(\u2_Display/n657 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c4 ),
    .o({\u2_Display/lt29_c5 ,open_n3752}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_5  (
    .a(\u2_Display/n656 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c5 ),
    .o({\u2_Display/lt29_c6 ,open_n3753}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_6  (
    .a(\u2_Display/n655 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c6 ),
    .o({\u2_Display/lt29_c7 ,open_n3754}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_7  (
    .a(\u2_Display/n654 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c7 ),
    .o({\u2_Display/lt29_c8 ,open_n3755}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_8  (
    .a(\u2_Display/n653 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c8 ),
    .o({\u2_Display/lt29_c9 ,open_n3756}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_9  (
    .a(\u2_Display/n652 ),
    .b(1'b0),
    .c(\u2_Display/lt29_c9 ),
    .o({\u2_Display/lt29_c10 ,open_n3757}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt29_cin  (
    .a(1'b0),
    .o({\u2_Display/lt29_c0 ,open_n3760}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt29_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt29_c32 ),
    .o({open_n3761,\u2_Display/n662 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt2_2_0  (
    .a(lcd_ypos[0]),
    .b(\u2_Display/j [0]),
    .c(\u2_Display/lt2_2_c0 ),
    .o({\u2_Display/lt2_2_c1 ,open_n3762}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt2_2_1  (
    .a(lcd_ypos[1]),
    .b(\u2_Display/j [1]),
    .c(\u2_Display/lt2_2_c1 ),
    .o({\u2_Display/lt2_2_c2 ,open_n3763}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt2_2_10  (
    .a(lcd_ypos[10]),
    .b(1'b1),
    .c(\u2_Display/lt2_2_c10 ),
    .o({\u2_Display/lt2_2_c11 ,open_n3764}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt2_2_11  (
    .a(lcd_ypos[11]),
    .b(1'b0),
    .c(\u2_Display/lt2_2_c11 ),
    .o({\u2_Display/lt2_2_c12 ,open_n3765}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt2_2_2  (
    .a(lcd_ypos[2]),
    .b(\u2_Display/j [2]),
    .c(\u2_Display/lt2_2_c2 ),
    .o({\u2_Display/lt2_2_c3 ,open_n3766}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt2_2_3  (
    .a(lcd_ypos[3]),
    .b(\u2_Display/j [3]),
    .c(\u2_Display/lt2_2_c3 ),
    .o({\u2_Display/lt2_2_c4 ,open_n3767}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt2_2_4  (
    .a(lcd_ypos[4]),
    .b(\u2_Display/j [4]),
    .c(\u2_Display/lt2_2_c4 ),
    .o({\u2_Display/lt2_2_c5 ,open_n3768}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt2_2_5  (
    .a(lcd_ypos[5]),
    .b(\u2_Display/j [5]),
    .c(\u2_Display/lt2_2_c5 ),
    .o({\u2_Display/lt2_2_c6 ,open_n3769}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt2_2_6  (
    .a(lcd_ypos[6]),
    .b(\u2_Display/j [6]),
    .c(\u2_Display/lt2_2_c6 ),
    .o({\u2_Display/lt2_2_c7 ,open_n3770}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt2_2_7  (
    .a(lcd_ypos[7]),
    .b(\u2_Display/j [7]),
    .c(\u2_Display/lt2_2_c7 ),
    .o({\u2_Display/lt2_2_c8 ,open_n3771}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt2_2_8  (
    .a(lcd_ypos[8]),
    .b(\u2_Display/j [8]),
    .c(\u2_Display/lt2_2_c8 ),
    .o({\u2_Display/lt2_2_c9 ,open_n3772}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt2_2_9  (
    .a(lcd_ypos[9]),
    .b(\u2_Display/j [9]),
    .c(\u2_Display/lt2_2_c9 ),
    .o({\u2_Display/lt2_2_c10 ,open_n3773}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt2_2_cin  (
    .a(1'b0),
    .o({\u2_Display/lt2_2_c0 ,open_n3776}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt2_2_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt2_2_c12 ),
    .o({open_n3777,\u2_Display/n48 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_0  (
    .a(\u2_Display/n696 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c0 ),
    .o({\u2_Display/lt30_c1 ,open_n3778}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_1  (
    .a(\u2_Display/n695 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c1 ),
    .o({\u2_Display/lt30_c2 ,open_n3779}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_10  (
    .a(\u2_Display/n686 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c10 ),
    .o({\u2_Display/lt30_c11 ,open_n3780}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_11  (
    .a(\u2_Display/n685 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c11 ),
    .o({\u2_Display/lt30_c12 ,open_n3781}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_12  (
    .a(\u2_Display/n684 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c12 ),
    .o({\u2_Display/lt30_c13 ,open_n3782}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_13  (
    .a(\u2_Display/n683 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c13 ),
    .o({\u2_Display/lt30_c14 ,open_n3783}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_14  (
    .a(\u2_Display/n682 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c14 ),
    .o({\u2_Display/lt30_c15 ,open_n3784}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_15  (
    .a(\u2_Display/n681 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c15 ),
    .o({\u2_Display/lt30_c16 ,open_n3785}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_16  (
    .a(\u2_Display/n680 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c16 ),
    .o({\u2_Display/lt30_c17 ,open_n3786}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_17  (
    .a(\u2_Display/n679 ),
    .b(1'b1),
    .c(\u2_Display/lt30_c17 ),
    .o({\u2_Display/lt30_c18 ,open_n3787}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_18  (
    .a(\u2_Display/n678 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c18 ),
    .o({\u2_Display/lt30_c19 ,open_n3788}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_19  (
    .a(\u2_Display/n677 ),
    .b(1'b1),
    .c(\u2_Display/lt30_c19 ),
    .o({\u2_Display/lt30_c20 ,open_n3789}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_2  (
    .a(\u2_Display/n694 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c2 ),
    .o({\u2_Display/lt30_c3 ,open_n3790}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_20  (
    .a(\u2_Display/n676 ),
    .b(1'b1),
    .c(\u2_Display/lt30_c20 ),
    .o({\u2_Display/lt30_c21 ,open_n3791}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_21  (
    .a(\u2_Display/n675 ),
    .b(1'b1),
    .c(\u2_Display/lt30_c21 ),
    .o({\u2_Display/lt30_c22 ,open_n3792}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_22  (
    .a(\u2_Display/n674 ),
    .b(1'b1),
    .c(\u2_Display/lt30_c22 ),
    .o({\u2_Display/lt30_c23 ,open_n3793}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_23  (
    .a(\u2_Display/n673 ),
    .b(1'b1),
    .c(\u2_Display/lt30_c23 ),
    .o({\u2_Display/lt30_c24 ,open_n3794}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_24  (
    .a(\u2_Display/n672 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c24 ),
    .o({\u2_Display/lt30_c25 ,open_n3795}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_25  (
    .a(\u2_Display/n671 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c25 ),
    .o({\u2_Display/lt30_c26 ,open_n3796}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_26  (
    .a(\u2_Display/n670 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c26 ),
    .o({\u2_Display/lt30_c27 ,open_n3797}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_27  (
    .a(\u2_Display/n669 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c27 ),
    .o({\u2_Display/lt30_c28 ,open_n3798}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_28  (
    .a(\u2_Display/n668 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c28 ),
    .o({\u2_Display/lt30_c29 ,open_n3799}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_29  (
    .a(\u2_Display/n667 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c29 ),
    .o({\u2_Display/lt30_c30 ,open_n3800}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_3  (
    .a(\u2_Display/n693 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c3 ),
    .o({\u2_Display/lt30_c4 ,open_n3801}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_30  (
    .a(\u2_Display/n666 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c30 ),
    .o({\u2_Display/lt30_c31 ,open_n3802}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_31  (
    .a(\u2_Display/n665 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c31 ),
    .o({\u2_Display/lt30_c32 ,open_n3803}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_4  (
    .a(\u2_Display/n692 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c4 ),
    .o({\u2_Display/lt30_c5 ,open_n3804}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_5  (
    .a(\u2_Display/n691 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c5 ),
    .o({\u2_Display/lt30_c6 ,open_n3805}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_6  (
    .a(\u2_Display/n690 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c6 ),
    .o({\u2_Display/lt30_c7 ,open_n3806}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_7  (
    .a(\u2_Display/n689 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c7 ),
    .o({\u2_Display/lt30_c8 ,open_n3807}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_8  (
    .a(\u2_Display/n688 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c8 ),
    .o({\u2_Display/lt30_c9 ,open_n3808}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_9  (
    .a(\u2_Display/n687 ),
    .b(1'b0),
    .c(\u2_Display/lt30_c9 ),
    .o({\u2_Display/lt30_c10 ,open_n3809}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt30_cin  (
    .a(1'b0),
    .o({\u2_Display/lt30_c0 ,open_n3812}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt30_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt30_c32 ),
    .o({open_n3813,\u2_Display/n697 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_0  (
    .a(\u2_Display/n731 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c0 ),
    .o({\u2_Display/lt31_c1 ,open_n3814}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_1  (
    .a(\u2_Display/n730 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c1 ),
    .o({\u2_Display/lt31_c2 ,open_n3815}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_10  (
    .a(\u2_Display/n721 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c10 ),
    .o({\u2_Display/lt31_c11 ,open_n3816}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_11  (
    .a(\u2_Display/n720 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c11 ),
    .o({\u2_Display/lt31_c12 ,open_n3817}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_12  (
    .a(\u2_Display/n719 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c12 ),
    .o({\u2_Display/lt31_c13 ,open_n3818}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_13  (
    .a(\u2_Display/n718 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c13 ),
    .o({\u2_Display/lt31_c14 ,open_n3819}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_14  (
    .a(\u2_Display/n717 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c14 ),
    .o({\u2_Display/lt31_c15 ,open_n3820}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_15  (
    .a(\u2_Display/n716 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c15 ),
    .o({\u2_Display/lt31_c16 ,open_n3821}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_16  (
    .a(\u2_Display/n715 ),
    .b(1'b1),
    .c(\u2_Display/lt31_c16 ),
    .o({\u2_Display/lt31_c17 ,open_n3822}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_17  (
    .a(\u2_Display/n714 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c17 ),
    .o({\u2_Display/lt31_c18 ,open_n3823}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_18  (
    .a(\u2_Display/n713 ),
    .b(1'b1),
    .c(\u2_Display/lt31_c18 ),
    .o({\u2_Display/lt31_c19 ,open_n3824}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_19  (
    .a(\u2_Display/n712 ),
    .b(1'b1),
    .c(\u2_Display/lt31_c19 ),
    .o({\u2_Display/lt31_c20 ,open_n3825}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_2  (
    .a(\u2_Display/n729 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c2 ),
    .o({\u2_Display/lt31_c3 ,open_n3826}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_20  (
    .a(\u2_Display/n711 ),
    .b(1'b1),
    .c(\u2_Display/lt31_c20 ),
    .o({\u2_Display/lt31_c21 ,open_n3827}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_21  (
    .a(\u2_Display/n710 ),
    .b(1'b1),
    .c(\u2_Display/lt31_c21 ),
    .o({\u2_Display/lt31_c22 ,open_n3828}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_22  (
    .a(\u2_Display/n709 ),
    .b(1'b1),
    .c(\u2_Display/lt31_c22 ),
    .o({\u2_Display/lt31_c23 ,open_n3829}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_23  (
    .a(\u2_Display/n708 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c23 ),
    .o({\u2_Display/lt31_c24 ,open_n3830}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_24  (
    .a(\u2_Display/n707 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c24 ),
    .o({\u2_Display/lt31_c25 ,open_n3831}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_25  (
    .a(\u2_Display/n706 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c25 ),
    .o({\u2_Display/lt31_c26 ,open_n3832}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_26  (
    .a(\u2_Display/n705 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c26 ),
    .o({\u2_Display/lt31_c27 ,open_n3833}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_27  (
    .a(\u2_Display/n704 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c27 ),
    .o({\u2_Display/lt31_c28 ,open_n3834}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_28  (
    .a(\u2_Display/n703 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c28 ),
    .o({\u2_Display/lt31_c29 ,open_n3835}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_29  (
    .a(\u2_Display/n702 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c29 ),
    .o({\u2_Display/lt31_c30 ,open_n3836}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_3  (
    .a(\u2_Display/n728 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c3 ),
    .o({\u2_Display/lt31_c4 ,open_n3837}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_30  (
    .a(\u2_Display/n701 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c30 ),
    .o({\u2_Display/lt31_c31 ,open_n3838}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_31  (
    .a(\u2_Display/n700 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c31 ),
    .o({\u2_Display/lt31_c32 ,open_n3839}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_4  (
    .a(\u2_Display/n727 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c4 ),
    .o({\u2_Display/lt31_c5 ,open_n3840}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_5  (
    .a(\u2_Display/n726 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c5 ),
    .o({\u2_Display/lt31_c6 ,open_n3841}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_6  (
    .a(\u2_Display/n725 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c6 ),
    .o({\u2_Display/lt31_c7 ,open_n3842}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_7  (
    .a(\u2_Display/n724 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c7 ),
    .o({\u2_Display/lt31_c8 ,open_n3843}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_8  (
    .a(\u2_Display/n723 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c8 ),
    .o({\u2_Display/lt31_c9 ,open_n3844}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_9  (
    .a(\u2_Display/n722 ),
    .b(1'b0),
    .c(\u2_Display/lt31_c9 ),
    .o({\u2_Display/lt31_c10 ,open_n3845}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt31_cin  (
    .a(1'b0),
    .o({\u2_Display/lt31_c0 ,open_n3848}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt31_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt31_c32 ),
    .o({open_n3849,\u2_Display/n732 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_0  (
    .a(\u2_Display/n766 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c0 ),
    .o({\u2_Display/lt32_c1 ,open_n3850}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_1  (
    .a(\u2_Display/n765 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c1 ),
    .o({\u2_Display/lt32_c2 ,open_n3851}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_10  (
    .a(\u2_Display/n756 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c10 ),
    .o({\u2_Display/lt32_c11 ,open_n3852}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_11  (
    .a(\u2_Display/n755 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c11 ),
    .o({\u2_Display/lt32_c12 ,open_n3853}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_12  (
    .a(\u2_Display/n754 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c12 ),
    .o({\u2_Display/lt32_c13 ,open_n3854}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_13  (
    .a(\u2_Display/n753 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c13 ),
    .o({\u2_Display/lt32_c14 ,open_n3855}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_14  (
    .a(\u2_Display/n752 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c14 ),
    .o({\u2_Display/lt32_c15 ,open_n3856}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_15  (
    .a(\u2_Display/n751 ),
    .b(1'b1),
    .c(\u2_Display/lt32_c15 ),
    .o({\u2_Display/lt32_c16 ,open_n3857}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_16  (
    .a(\u2_Display/n750 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c16 ),
    .o({\u2_Display/lt32_c17 ,open_n3858}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_17  (
    .a(\u2_Display/n749 ),
    .b(1'b1),
    .c(\u2_Display/lt32_c17 ),
    .o({\u2_Display/lt32_c18 ,open_n3859}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_18  (
    .a(\u2_Display/n748 ),
    .b(1'b1),
    .c(\u2_Display/lt32_c18 ),
    .o({\u2_Display/lt32_c19 ,open_n3860}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_19  (
    .a(\u2_Display/n747 ),
    .b(1'b1),
    .c(\u2_Display/lt32_c19 ),
    .o({\u2_Display/lt32_c20 ,open_n3861}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_2  (
    .a(\u2_Display/n764 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c2 ),
    .o({\u2_Display/lt32_c3 ,open_n3862}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_20  (
    .a(\u2_Display/n746 ),
    .b(1'b1),
    .c(\u2_Display/lt32_c20 ),
    .o({\u2_Display/lt32_c21 ,open_n3863}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_21  (
    .a(\u2_Display/n745 ),
    .b(1'b1),
    .c(\u2_Display/lt32_c21 ),
    .o({\u2_Display/lt32_c22 ,open_n3864}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_22  (
    .a(\u2_Display/n744 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c22 ),
    .o({\u2_Display/lt32_c23 ,open_n3865}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_23  (
    .a(\u2_Display/n743 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c23 ),
    .o({\u2_Display/lt32_c24 ,open_n3866}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_24  (
    .a(\u2_Display/n742 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c24 ),
    .o({\u2_Display/lt32_c25 ,open_n3867}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_25  (
    .a(\u2_Display/n741 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c25 ),
    .o({\u2_Display/lt32_c26 ,open_n3868}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_26  (
    .a(\u2_Display/n740 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c26 ),
    .o({\u2_Display/lt32_c27 ,open_n3869}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_27  (
    .a(\u2_Display/n739 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c27 ),
    .o({\u2_Display/lt32_c28 ,open_n3870}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_28  (
    .a(\u2_Display/n738 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c28 ),
    .o({\u2_Display/lt32_c29 ,open_n3871}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_29  (
    .a(\u2_Display/n737 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c29 ),
    .o({\u2_Display/lt32_c30 ,open_n3872}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_3  (
    .a(\u2_Display/n763 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c3 ),
    .o({\u2_Display/lt32_c4 ,open_n3873}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_30  (
    .a(\u2_Display/n736 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c30 ),
    .o({\u2_Display/lt32_c31 ,open_n3874}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_31  (
    .a(\u2_Display/n735 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c31 ),
    .o({\u2_Display/lt32_c32 ,open_n3875}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_4  (
    .a(\u2_Display/n762 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c4 ),
    .o({\u2_Display/lt32_c5 ,open_n3876}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_5  (
    .a(\u2_Display/n761 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c5 ),
    .o({\u2_Display/lt32_c6 ,open_n3877}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_6  (
    .a(\u2_Display/n760 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c6 ),
    .o({\u2_Display/lt32_c7 ,open_n3878}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_7  (
    .a(\u2_Display/n759 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c7 ),
    .o({\u2_Display/lt32_c8 ,open_n3879}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_8  (
    .a(\u2_Display/n758 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c8 ),
    .o({\u2_Display/lt32_c9 ,open_n3880}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_9  (
    .a(\u2_Display/n757 ),
    .b(1'b0),
    .c(\u2_Display/lt32_c9 ),
    .o({\u2_Display/lt32_c10 ,open_n3881}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt32_cin  (
    .a(1'b0),
    .o({\u2_Display/lt32_c0 ,open_n3884}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt32_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt32_c32 ),
    .o({open_n3885,\u2_Display/n767 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_0  (
    .a(\u2_Display/n801 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c0 ),
    .o({\u2_Display/lt33_c1 ,open_n3886}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_1  (
    .a(\u2_Display/n800 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c1 ),
    .o({\u2_Display/lt33_c2 ,open_n3887}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_10  (
    .a(\u2_Display/n791 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c10 ),
    .o({\u2_Display/lt33_c11 ,open_n3888}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_11  (
    .a(\u2_Display/n790 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c11 ),
    .o({\u2_Display/lt33_c12 ,open_n3889}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_12  (
    .a(\u2_Display/n789 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c12 ),
    .o({\u2_Display/lt33_c13 ,open_n3890}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_13  (
    .a(\u2_Display/n788 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c13 ),
    .o({\u2_Display/lt33_c14 ,open_n3891}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_14  (
    .a(\u2_Display/n787 ),
    .b(1'b1),
    .c(\u2_Display/lt33_c14 ),
    .o({\u2_Display/lt33_c15 ,open_n3892}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_15  (
    .a(\u2_Display/n786 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c15 ),
    .o({\u2_Display/lt33_c16 ,open_n3893}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_16  (
    .a(\u2_Display/n785 ),
    .b(1'b1),
    .c(\u2_Display/lt33_c16 ),
    .o({\u2_Display/lt33_c17 ,open_n3894}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_17  (
    .a(\u2_Display/n784 ),
    .b(1'b1),
    .c(\u2_Display/lt33_c17 ),
    .o({\u2_Display/lt33_c18 ,open_n3895}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_18  (
    .a(\u2_Display/n783 ),
    .b(1'b1),
    .c(\u2_Display/lt33_c18 ),
    .o({\u2_Display/lt33_c19 ,open_n3896}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_19  (
    .a(\u2_Display/n782 ),
    .b(1'b1),
    .c(\u2_Display/lt33_c19 ),
    .o({\u2_Display/lt33_c20 ,open_n3897}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_2  (
    .a(\u2_Display/n799 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c2 ),
    .o({\u2_Display/lt33_c3 ,open_n3898}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_20  (
    .a(\u2_Display/n781 ),
    .b(1'b1),
    .c(\u2_Display/lt33_c20 ),
    .o({\u2_Display/lt33_c21 ,open_n3899}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_21  (
    .a(\u2_Display/n780 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c21 ),
    .o({\u2_Display/lt33_c22 ,open_n3900}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_22  (
    .a(\u2_Display/n779 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c22 ),
    .o({\u2_Display/lt33_c23 ,open_n3901}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_23  (
    .a(\u2_Display/n778 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c23 ),
    .o({\u2_Display/lt33_c24 ,open_n3902}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_24  (
    .a(\u2_Display/n777 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c24 ),
    .o({\u2_Display/lt33_c25 ,open_n3903}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_25  (
    .a(\u2_Display/n776 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c25 ),
    .o({\u2_Display/lt33_c26 ,open_n3904}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_26  (
    .a(\u2_Display/n775 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c26 ),
    .o({\u2_Display/lt33_c27 ,open_n3905}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_27  (
    .a(\u2_Display/n774 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c27 ),
    .o({\u2_Display/lt33_c28 ,open_n3906}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_28  (
    .a(\u2_Display/n773 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c28 ),
    .o({\u2_Display/lt33_c29 ,open_n3907}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_29  (
    .a(\u2_Display/n772 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c29 ),
    .o({\u2_Display/lt33_c30 ,open_n3908}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_3  (
    .a(\u2_Display/n798 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c3 ),
    .o({\u2_Display/lt33_c4 ,open_n3909}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_30  (
    .a(\u2_Display/n771 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c30 ),
    .o({\u2_Display/lt33_c31 ,open_n3910}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_31  (
    .a(\u2_Display/n770 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c31 ),
    .o({\u2_Display/lt33_c32 ,open_n3911}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_4  (
    .a(\u2_Display/n797 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c4 ),
    .o({\u2_Display/lt33_c5 ,open_n3912}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_5  (
    .a(\u2_Display/n796 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c5 ),
    .o({\u2_Display/lt33_c6 ,open_n3913}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_6  (
    .a(\u2_Display/n795 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c6 ),
    .o({\u2_Display/lt33_c7 ,open_n3914}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_7  (
    .a(\u2_Display/n794 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c7 ),
    .o({\u2_Display/lt33_c8 ,open_n3915}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_8  (
    .a(\u2_Display/n793 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c8 ),
    .o({\u2_Display/lt33_c9 ,open_n3916}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_9  (
    .a(\u2_Display/n792 ),
    .b(1'b0),
    .c(\u2_Display/lt33_c9 ),
    .o({\u2_Display/lt33_c10 ,open_n3917}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt33_cin  (
    .a(1'b0),
    .o({\u2_Display/lt33_c0 ,open_n3920}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt33_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt33_c32 ),
    .o({open_n3921,\u2_Display/n802 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_0  (
    .a(\u2_Display/n836 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c0 ),
    .o({\u2_Display/lt34_c1 ,open_n3922}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_1  (
    .a(\u2_Display/n835 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c1 ),
    .o({\u2_Display/lt34_c2 ,open_n3923}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_10  (
    .a(\u2_Display/n826 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c10 ),
    .o({\u2_Display/lt34_c11 ,open_n3924}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_11  (
    .a(\u2_Display/n825 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c11 ),
    .o({\u2_Display/lt34_c12 ,open_n3925}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_12  (
    .a(\u2_Display/n824 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c12 ),
    .o({\u2_Display/lt34_c13 ,open_n3926}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_13  (
    .a(\u2_Display/n823 ),
    .b(1'b1),
    .c(\u2_Display/lt34_c13 ),
    .o({\u2_Display/lt34_c14 ,open_n3927}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_14  (
    .a(\u2_Display/n822 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c14 ),
    .o({\u2_Display/lt34_c15 ,open_n3928}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_15  (
    .a(\u2_Display/n821 ),
    .b(1'b1),
    .c(\u2_Display/lt34_c15 ),
    .o({\u2_Display/lt34_c16 ,open_n3929}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_16  (
    .a(\u2_Display/n820 ),
    .b(1'b1),
    .c(\u2_Display/lt34_c16 ),
    .o({\u2_Display/lt34_c17 ,open_n3930}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_17  (
    .a(\u2_Display/n819 ),
    .b(1'b1),
    .c(\u2_Display/lt34_c17 ),
    .o({\u2_Display/lt34_c18 ,open_n3931}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_18  (
    .a(\u2_Display/n818 ),
    .b(1'b1),
    .c(\u2_Display/lt34_c18 ),
    .o({\u2_Display/lt34_c19 ,open_n3932}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_19  (
    .a(\u2_Display/n817 ),
    .b(1'b1),
    .c(\u2_Display/lt34_c19 ),
    .o({\u2_Display/lt34_c20 ,open_n3933}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_2  (
    .a(\u2_Display/n834 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c2 ),
    .o({\u2_Display/lt34_c3 ,open_n3934}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_20  (
    .a(\u2_Display/n816 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c20 ),
    .o({\u2_Display/lt34_c21 ,open_n3935}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_21  (
    .a(\u2_Display/n815 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c21 ),
    .o({\u2_Display/lt34_c22 ,open_n3936}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_22  (
    .a(\u2_Display/n814 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c22 ),
    .o({\u2_Display/lt34_c23 ,open_n3937}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_23  (
    .a(\u2_Display/n813 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c23 ),
    .o({\u2_Display/lt34_c24 ,open_n3938}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_24  (
    .a(\u2_Display/n812 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c24 ),
    .o({\u2_Display/lt34_c25 ,open_n3939}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_25  (
    .a(\u2_Display/n811 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c25 ),
    .o({\u2_Display/lt34_c26 ,open_n3940}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_26  (
    .a(\u2_Display/n810 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c26 ),
    .o({\u2_Display/lt34_c27 ,open_n3941}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_27  (
    .a(\u2_Display/n809 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c27 ),
    .o({\u2_Display/lt34_c28 ,open_n3942}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_28  (
    .a(\u2_Display/n808 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c28 ),
    .o({\u2_Display/lt34_c29 ,open_n3943}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_29  (
    .a(\u2_Display/n807 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c29 ),
    .o({\u2_Display/lt34_c30 ,open_n3944}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_3  (
    .a(\u2_Display/n833 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c3 ),
    .o({\u2_Display/lt34_c4 ,open_n3945}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_30  (
    .a(\u2_Display/n806 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c30 ),
    .o({\u2_Display/lt34_c31 ,open_n3946}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_31  (
    .a(\u2_Display/n805 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c31 ),
    .o({\u2_Display/lt34_c32 ,open_n3947}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_4  (
    .a(\u2_Display/n832 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c4 ),
    .o({\u2_Display/lt34_c5 ,open_n3948}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_5  (
    .a(\u2_Display/n831 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c5 ),
    .o({\u2_Display/lt34_c6 ,open_n3949}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_6  (
    .a(\u2_Display/n830 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c6 ),
    .o({\u2_Display/lt34_c7 ,open_n3950}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_7  (
    .a(\u2_Display/n829 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c7 ),
    .o({\u2_Display/lt34_c8 ,open_n3951}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_8  (
    .a(\u2_Display/n828 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c8 ),
    .o({\u2_Display/lt34_c9 ,open_n3952}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_9  (
    .a(\u2_Display/n827 ),
    .b(1'b0),
    .c(\u2_Display/lt34_c9 ),
    .o({\u2_Display/lt34_c10 ,open_n3953}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt34_cin  (
    .a(1'b0),
    .o({\u2_Display/lt34_c0 ,open_n3956}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt34_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt34_c32 ),
    .o({open_n3957,\u2_Display/n837 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_0  (
    .a(\u2_Display/n871 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c0 ),
    .o({\u2_Display/lt35_c1 ,open_n3958}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_1  (
    .a(\u2_Display/n870 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c1 ),
    .o({\u2_Display/lt35_c2 ,open_n3959}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_10  (
    .a(\u2_Display/n861 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c10 ),
    .o({\u2_Display/lt35_c11 ,open_n3960}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_11  (
    .a(\u2_Display/n860 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c11 ),
    .o({\u2_Display/lt35_c12 ,open_n3961}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_12  (
    .a(\u2_Display/n859 ),
    .b(1'b1),
    .c(\u2_Display/lt35_c12 ),
    .o({\u2_Display/lt35_c13 ,open_n3962}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_13  (
    .a(\u2_Display/n858 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c13 ),
    .o({\u2_Display/lt35_c14 ,open_n3963}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_14  (
    .a(\u2_Display/n857 ),
    .b(1'b1),
    .c(\u2_Display/lt35_c14 ),
    .o({\u2_Display/lt35_c15 ,open_n3964}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_15  (
    .a(\u2_Display/n856 ),
    .b(1'b1),
    .c(\u2_Display/lt35_c15 ),
    .o({\u2_Display/lt35_c16 ,open_n3965}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_16  (
    .a(\u2_Display/n855 ),
    .b(1'b1),
    .c(\u2_Display/lt35_c16 ),
    .o({\u2_Display/lt35_c17 ,open_n3966}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_17  (
    .a(\u2_Display/n854 ),
    .b(1'b1),
    .c(\u2_Display/lt35_c17 ),
    .o({\u2_Display/lt35_c18 ,open_n3967}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_18  (
    .a(\u2_Display/n853 ),
    .b(1'b1),
    .c(\u2_Display/lt35_c18 ),
    .o({\u2_Display/lt35_c19 ,open_n3968}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_19  (
    .a(\u2_Display/n852 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c19 ),
    .o({\u2_Display/lt35_c20 ,open_n3969}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_2  (
    .a(\u2_Display/n869 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c2 ),
    .o({\u2_Display/lt35_c3 ,open_n3970}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_20  (
    .a(\u2_Display/n851 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c20 ),
    .o({\u2_Display/lt35_c21 ,open_n3971}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_21  (
    .a(\u2_Display/n850 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c21 ),
    .o({\u2_Display/lt35_c22 ,open_n3972}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_22  (
    .a(\u2_Display/n849 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c22 ),
    .o({\u2_Display/lt35_c23 ,open_n3973}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_23  (
    .a(\u2_Display/n848 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c23 ),
    .o({\u2_Display/lt35_c24 ,open_n3974}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_24  (
    .a(\u2_Display/n847 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c24 ),
    .o({\u2_Display/lt35_c25 ,open_n3975}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_25  (
    .a(\u2_Display/n846 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c25 ),
    .o({\u2_Display/lt35_c26 ,open_n3976}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_26  (
    .a(\u2_Display/n845 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c26 ),
    .o({\u2_Display/lt35_c27 ,open_n3977}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_27  (
    .a(\u2_Display/n844 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c27 ),
    .o({\u2_Display/lt35_c28 ,open_n3978}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_28  (
    .a(\u2_Display/n843 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c28 ),
    .o({\u2_Display/lt35_c29 ,open_n3979}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_29  (
    .a(\u2_Display/n842 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c29 ),
    .o({\u2_Display/lt35_c30 ,open_n3980}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_3  (
    .a(\u2_Display/n868 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c3 ),
    .o({\u2_Display/lt35_c4 ,open_n3981}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_30  (
    .a(\u2_Display/n841 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c30 ),
    .o({\u2_Display/lt35_c31 ,open_n3982}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_31  (
    .a(\u2_Display/n840 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c31 ),
    .o({\u2_Display/lt35_c32 ,open_n3983}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_4  (
    .a(\u2_Display/n867 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c4 ),
    .o({\u2_Display/lt35_c5 ,open_n3984}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_5  (
    .a(\u2_Display/n866 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c5 ),
    .o({\u2_Display/lt35_c6 ,open_n3985}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_6  (
    .a(\u2_Display/n865 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c6 ),
    .o({\u2_Display/lt35_c7 ,open_n3986}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_7  (
    .a(\u2_Display/n864 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c7 ),
    .o({\u2_Display/lt35_c8 ,open_n3987}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_8  (
    .a(\u2_Display/n863 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c8 ),
    .o({\u2_Display/lt35_c9 ,open_n3988}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_9  (
    .a(\u2_Display/n862 ),
    .b(1'b0),
    .c(\u2_Display/lt35_c9 ),
    .o({\u2_Display/lt35_c10 ,open_n3989}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt35_cin  (
    .a(1'b0),
    .o({\u2_Display/lt35_c0 ,open_n3992}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt35_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt35_c32 ),
    .o({open_n3993,\u2_Display/n872 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_0  (
    .a(\u2_Display/n906 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c0 ),
    .o({\u2_Display/lt36_c1 ,open_n3994}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_1  (
    .a(\u2_Display/n905 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c1 ),
    .o({\u2_Display/lt36_c2 ,open_n3995}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_10  (
    .a(\u2_Display/n896 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c10 ),
    .o({\u2_Display/lt36_c11 ,open_n3996}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_11  (
    .a(\u2_Display/n895 ),
    .b(1'b1),
    .c(\u2_Display/lt36_c11 ),
    .o({\u2_Display/lt36_c12 ,open_n3997}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_12  (
    .a(\u2_Display/n894 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c12 ),
    .o({\u2_Display/lt36_c13 ,open_n3998}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_13  (
    .a(\u2_Display/n893 ),
    .b(1'b1),
    .c(\u2_Display/lt36_c13 ),
    .o({\u2_Display/lt36_c14 ,open_n3999}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_14  (
    .a(\u2_Display/n892 ),
    .b(1'b1),
    .c(\u2_Display/lt36_c14 ),
    .o({\u2_Display/lt36_c15 ,open_n4000}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_15  (
    .a(\u2_Display/n891 ),
    .b(1'b1),
    .c(\u2_Display/lt36_c15 ),
    .o({\u2_Display/lt36_c16 ,open_n4001}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_16  (
    .a(\u2_Display/n890 ),
    .b(1'b1),
    .c(\u2_Display/lt36_c16 ),
    .o({\u2_Display/lt36_c17 ,open_n4002}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_17  (
    .a(\u2_Display/n889 ),
    .b(1'b1),
    .c(\u2_Display/lt36_c17 ),
    .o({\u2_Display/lt36_c18 ,open_n4003}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_18  (
    .a(\u2_Display/n888 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c18 ),
    .o({\u2_Display/lt36_c19 ,open_n4004}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_19  (
    .a(\u2_Display/n887 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c19 ),
    .o({\u2_Display/lt36_c20 ,open_n4005}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_2  (
    .a(\u2_Display/n904 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c2 ),
    .o({\u2_Display/lt36_c3 ,open_n4006}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_20  (
    .a(\u2_Display/n886 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c20 ),
    .o({\u2_Display/lt36_c21 ,open_n4007}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_21  (
    .a(\u2_Display/n885 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c21 ),
    .o({\u2_Display/lt36_c22 ,open_n4008}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_22  (
    .a(\u2_Display/n884 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c22 ),
    .o({\u2_Display/lt36_c23 ,open_n4009}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_23  (
    .a(\u2_Display/n883 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c23 ),
    .o({\u2_Display/lt36_c24 ,open_n4010}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_24  (
    .a(\u2_Display/n882 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c24 ),
    .o({\u2_Display/lt36_c25 ,open_n4011}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_25  (
    .a(\u2_Display/n881 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c25 ),
    .o({\u2_Display/lt36_c26 ,open_n4012}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_26  (
    .a(\u2_Display/n880 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c26 ),
    .o({\u2_Display/lt36_c27 ,open_n4013}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_27  (
    .a(\u2_Display/n879 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c27 ),
    .o({\u2_Display/lt36_c28 ,open_n4014}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_28  (
    .a(\u2_Display/n878 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c28 ),
    .o({\u2_Display/lt36_c29 ,open_n4015}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_29  (
    .a(\u2_Display/n877 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c29 ),
    .o({\u2_Display/lt36_c30 ,open_n4016}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_3  (
    .a(\u2_Display/n903 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c3 ),
    .o({\u2_Display/lt36_c4 ,open_n4017}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_30  (
    .a(\u2_Display/n876 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c30 ),
    .o({\u2_Display/lt36_c31 ,open_n4018}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_31  (
    .a(\u2_Display/n875 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c31 ),
    .o({\u2_Display/lt36_c32 ,open_n4019}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_4  (
    .a(\u2_Display/n902 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c4 ),
    .o({\u2_Display/lt36_c5 ,open_n4020}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_5  (
    .a(\u2_Display/n901 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c5 ),
    .o({\u2_Display/lt36_c6 ,open_n4021}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_6  (
    .a(\u2_Display/n900 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c6 ),
    .o({\u2_Display/lt36_c7 ,open_n4022}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_7  (
    .a(\u2_Display/n899 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c7 ),
    .o({\u2_Display/lt36_c8 ,open_n4023}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_8  (
    .a(\u2_Display/n898 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c8 ),
    .o({\u2_Display/lt36_c9 ,open_n4024}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_9  (
    .a(\u2_Display/n897 ),
    .b(1'b0),
    .c(\u2_Display/lt36_c9 ),
    .o({\u2_Display/lt36_c10 ,open_n4025}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt36_cin  (
    .a(1'b0),
    .o({\u2_Display/lt36_c0 ,open_n4028}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt36_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt36_c32 ),
    .o({open_n4029,\u2_Display/n907 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_0  (
    .a(\u2_Display/n941 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c0 ),
    .o({\u2_Display/lt37_c1 ,open_n4030}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_1  (
    .a(\u2_Display/n940 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c1 ),
    .o({\u2_Display/lt37_c2 ,open_n4031}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_10  (
    .a(\u2_Display/n931 ),
    .b(1'b1),
    .c(\u2_Display/lt37_c10 ),
    .o({\u2_Display/lt37_c11 ,open_n4032}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_11  (
    .a(\u2_Display/n930 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c11 ),
    .o({\u2_Display/lt37_c12 ,open_n4033}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_12  (
    .a(\u2_Display/n929 ),
    .b(1'b1),
    .c(\u2_Display/lt37_c12 ),
    .o({\u2_Display/lt37_c13 ,open_n4034}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_13  (
    .a(\u2_Display/n928 ),
    .b(1'b1),
    .c(\u2_Display/lt37_c13 ),
    .o({\u2_Display/lt37_c14 ,open_n4035}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_14  (
    .a(\u2_Display/n927 ),
    .b(1'b1),
    .c(\u2_Display/lt37_c14 ),
    .o({\u2_Display/lt37_c15 ,open_n4036}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_15  (
    .a(\u2_Display/n926 ),
    .b(1'b1),
    .c(\u2_Display/lt37_c15 ),
    .o({\u2_Display/lt37_c16 ,open_n4037}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_16  (
    .a(\u2_Display/n925 ),
    .b(1'b1),
    .c(\u2_Display/lt37_c16 ),
    .o({\u2_Display/lt37_c17 ,open_n4038}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_17  (
    .a(\u2_Display/n924 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c17 ),
    .o({\u2_Display/lt37_c18 ,open_n4039}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_18  (
    .a(\u2_Display/n923 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c18 ),
    .o({\u2_Display/lt37_c19 ,open_n4040}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_19  (
    .a(\u2_Display/n922 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c19 ),
    .o({\u2_Display/lt37_c20 ,open_n4041}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_2  (
    .a(\u2_Display/n939 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c2 ),
    .o({\u2_Display/lt37_c3 ,open_n4042}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_20  (
    .a(\u2_Display/n921 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c20 ),
    .o({\u2_Display/lt37_c21 ,open_n4043}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_21  (
    .a(\u2_Display/n920 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c21 ),
    .o({\u2_Display/lt37_c22 ,open_n4044}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_22  (
    .a(\u2_Display/n919 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c22 ),
    .o({\u2_Display/lt37_c23 ,open_n4045}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_23  (
    .a(\u2_Display/n918 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c23 ),
    .o({\u2_Display/lt37_c24 ,open_n4046}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_24  (
    .a(\u2_Display/n917 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c24 ),
    .o({\u2_Display/lt37_c25 ,open_n4047}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_25  (
    .a(\u2_Display/n916 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c25 ),
    .o({\u2_Display/lt37_c26 ,open_n4048}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_26  (
    .a(\u2_Display/n915 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c26 ),
    .o({\u2_Display/lt37_c27 ,open_n4049}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_27  (
    .a(\u2_Display/n914 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c27 ),
    .o({\u2_Display/lt37_c28 ,open_n4050}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_28  (
    .a(\u2_Display/n913 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c28 ),
    .o({\u2_Display/lt37_c29 ,open_n4051}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_29  (
    .a(\u2_Display/n912 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c29 ),
    .o({\u2_Display/lt37_c30 ,open_n4052}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_3  (
    .a(\u2_Display/n938 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c3 ),
    .o({\u2_Display/lt37_c4 ,open_n4053}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_30  (
    .a(\u2_Display/n911 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c30 ),
    .o({\u2_Display/lt37_c31 ,open_n4054}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_31  (
    .a(\u2_Display/n910 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c31 ),
    .o({\u2_Display/lt37_c32 ,open_n4055}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_4  (
    .a(\u2_Display/n937 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c4 ),
    .o({\u2_Display/lt37_c5 ,open_n4056}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_5  (
    .a(\u2_Display/n936 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c5 ),
    .o({\u2_Display/lt37_c6 ,open_n4057}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_6  (
    .a(\u2_Display/n935 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c6 ),
    .o({\u2_Display/lt37_c7 ,open_n4058}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_7  (
    .a(\u2_Display/n934 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c7 ),
    .o({\u2_Display/lt37_c8 ,open_n4059}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_8  (
    .a(\u2_Display/n933 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c8 ),
    .o({\u2_Display/lt37_c9 ,open_n4060}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_9  (
    .a(\u2_Display/n932 ),
    .b(1'b0),
    .c(\u2_Display/lt37_c9 ),
    .o({\u2_Display/lt37_c10 ,open_n4061}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt37_cin  (
    .a(1'b0),
    .o({\u2_Display/lt37_c0 ,open_n4064}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt37_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt37_c32 ),
    .o({open_n4065,\u2_Display/n942 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_0  (
    .a(\u2_Display/n976 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c0 ),
    .o({\u2_Display/lt38_c1 ,open_n4066}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_1  (
    .a(\u2_Display/n975 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c1 ),
    .o({\u2_Display/lt38_c2 ,open_n4067}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_10  (
    .a(\u2_Display/n966 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c10 ),
    .o({\u2_Display/lt38_c11 ,open_n4068}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_11  (
    .a(\u2_Display/n965 ),
    .b(1'b1),
    .c(\u2_Display/lt38_c11 ),
    .o({\u2_Display/lt38_c12 ,open_n4069}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_12  (
    .a(\u2_Display/n964 ),
    .b(1'b1),
    .c(\u2_Display/lt38_c12 ),
    .o({\u2_Display/lt38_c13 ,open_n4070}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_13  (
    .a(\u2_Display/n963 ),
    .b(1'b1),
    .c(\u2_Display/lt38_c13 ),
    .o({\u2_Display/lt38_c14 ,open_n4071}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_14  (
    .a(\u2_Display/n962 ),
    .b(1'b1),
    .c(\u2_Display/lt38_c14 ),
    .o({\u2_Display/lt38_c15 ,open_n4072}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_15  (
    .a(\u2_Display/n961 ),
    .b(1'b1),
    .c(\u2_Display/lt38_c15 ),
    .o({\u2_Display/lt38_c16 ,open_n4073}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_16  (
    .a(\u2_Display/n960 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c16 ),
    .o({\u2_Display/lt38_c17 ,open_n4074}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_17  (
    .a(\u2_Display/n959 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c17 ),
    .o({\u2_Display/lt38_c18 ,open_n4075}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_18  (
    .a(\u2_Display/n958 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c18 ),
    .o({\u2_Display/lt38_c19 ,open_n4076}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_19  (
    .a(\u2_Display/n957 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c19 ),
    .o({\u2_Display/lt38_c20 ,open_n4077}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_2  (
    .a(\u2_Display/n974 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c2 ),
    .o({\u2_Display/lt38_c3 ,open_n4078}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_20  (
    .a(\u2_Display/n956 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c20 ),
    .o({\u2_Display/lt38_c21 ,open_n4079}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_21  (
    .a(\u2_Display/n955 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c21 ),
    .o({\u2_Display/lt38_c22 ,open_n4080}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_22  (
    .a(\u2_Display/n954 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c22 ),
    .o({\u2_Display/lt38_c23 ,open_n4081}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_23  (
    .a(\u2_Display/n953 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c23 ),
    .o({\u2_Display/lt38_c24 ,open_n4082}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_24  (
    .a(\u2_Display/n952 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c24 ),
    .o({\u2_Display/lt38_c25 ,open_n4083}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_25  (
    .a(\u2_Display/n951 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c25 ),
    .o({\u2_Display/lt38_c26 ,open_n4084}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_26  (
    .a(\u2_Display/n950 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c26 ),
    .o({\u2_Display/lt38_c27 ,open_n4085}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_27  (
    .a(\u2_Display/n949 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c27 ),
    .o({\u2_Display/lt38_c28 ,open_n4086}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_28  (
    .a(\u2_Display/n948 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c28 ),
    .o({\u2_Display/lt38_c29 ,open_n4087}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_29  (
    .a(\u2_Display/n947 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c29 ),
    .o({\u2_Display/lt38_c30 ,open_n4088}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_3  (
    .a(\u2_Display/n973 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c3 ),
    .o({\u2_Display/lt38_c4 ,open_n4089}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_30  (
    .a(\u2_Display/n946 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c30 ),
    .o({\u2_Display/lt38_c31 ,open_n4090}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_31  (
    .a(\u2_Display/n945 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c31 ),
    .o({\u2_Display/lt38_c32 ,open_n4091}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_4  (
    .a(\u2_Display/n972 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c4 ),
    .o({\u2_Display/lt38_c5 ,open_n4092}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_5  (
    .a(\u2_Display/n971 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c5 ),
    .o({\u2_Display/lt38_c6 ,open_n4093}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_6  (
    .a(\u2_Display/n970 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c6 ),
    .o({\u2_Display/lt38_c7 ,open_n4094}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_7  (
    .a(\u2_Display/n969 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c7 ),
    .o({\u2_Display/lt38_c8 ,open_n4095}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_8  (
    .a(\u2_Display/n968 ),
    .b(1'b0),
    .c(\u2_Display/lt38_c8 ),
    .o({\u2_Display/lt38_c9 ,open_n4096}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_9  (
    .a(\u2_Display/n967 ),
    .b(1'b1),
    .c(\u2_Display/lt38_c9 ),
    .o({\u2_Display/lt38_c10 ,open_n4097}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt38_cin  (
    .a(1'b0),
    .o({\u2_Display/lt38_c0 ,open_n4100}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt38_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt38_c32 ),
    .o({open_n4101,\u2_Display/n977 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_0  (
    .a(\u2_Display/n1011 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c0 ),
    .o({\u2_Display/lt39_c1 ,open_n4102}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_1  (
    .a(\u2_Display/n1010 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c1 ),
    .o({\u2_Display/lt39_c2 ,open_n4103}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_10  (
    .a(\u2_Display/n1001 ),
    .b(1'b1),
    .c(\u2_Display/lt39_c10 ),
    .o({\u2_Display/lt39_c11 ,open_n4104}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_11  (
    .a(\u2_Display/n1000 ),
    .b(1'b1),
    .c(\u2_Display/lt39_c11 ),
    .o({\u2_Display/lt39_c12 ,open_n4105}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_12  (
    .a(\u2_Display/n999 ),
    .b(1'b1),
    .c(\u2_Display/lt39_c12 ),
    .o({\u2_Display/lt39_c13 ,open_n4106}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_13  (
    .a(\u2_Display/n998 ),
    .b(1'b1),
    .c(\u2_Display/lt39_c13 ),
    .o({\u2_Display/lt39_c14 ,open_n4107}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_14  (
    .a(\u2_Display/n997 ),
    .b(1'b1),
    .c(\u2_Display/lt39_c14 ),
    .o({\u2_Display/lt39_c15 ,open_n4108}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_15  (
    .a(\u2_Display/n996 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c15 ),
    .o({\u2_Display/lt39_c16 ,open_n4109}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_16  (
    .a(\u2_Display/n995 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c16 ),
    .o({\u2_Display/lt39_c17 ,open_n4110}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_17  (
    .a(\u2_Display/n994 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c17 ),
    .o({\u2_Display/lt39_c18 ,open_n4111}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_18  (
    .a(\u2_Display/n993 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c18 ),
    .o({\u2_Display/lt39_c19 ,open_n4112}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_19  (
    .a(\u2_Display/n992 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c19 ),
    .o({\u2_Display/lt39_c20 ,open_n4113}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_2  (
    .a(\u2_Display/n1009 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c2 ),
    .o({\u2_Display/lt39_c3 ,open_n4114}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_20  (
    .a(\u2_Display/n991 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c20 ),
    .o({\u2_Display/lt39_c21 ,open_n4115}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_21  (
    .a(\u2_Display/n990 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c21 ),
    .o({\u2_Display/lt39_c22 ,open_n4116}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_22  (
    .a(\u2_Display/n989 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c22 ),
    .o({\u2_Display/lt39_c23 ,open_n4117}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_23  (
    .a(\u2_Display/n988 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c23 ),
    .o({\u2_Display/lt39_c24 ,open_n4118}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_24  (
    .a(\u2_Display/n987 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c24 ),
    .o({\u2_Display/lt39_c25 ,open_n4119}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_25  (
    .a(\u2_Display/n986 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c25 ),
    .o({\u2_Display/lt39_c26 ,open_n4120}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_26  (
    .a(\u2_Display/n985 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c26 ),
    .o({\u2_Display/lt39_c27 ,open_n4121}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_27  (
    .a(\u2_Display/n984 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c27 ),
    .o({\u2_Display/lt39_c28 ,open_n4122}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_28  (
    .a(\u2_Display/n983 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c28 ),
    .o({\u2_Display/lt39_c29 ,open_n4123}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_29  (
    .a(\u2_Display/n982 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c29 ),
    .o({\u2_Display/lt39_c30 ,open_n4124}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_3  (
    .a(\u2_Display/n1008 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c3 ),
    .o({\u2_Display/lt39_c4 ,open_n4125}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_30  (
    .a(\u2_Display/n981 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c30 ),
    .o({\u2_Display/lt39_c31 ,open_n4126}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_31  (
    .a(\u2_Display/n980 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c31 ),
    .o({\u2_Display/lt39_c32 ,open_n4127}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_4  (
    .a(\u2_Display/n1007 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c4 ),
    .o({\u2_Display/lt39_c5 ,open_n4128}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_5  (
    .a(\u2_Display/n1006 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c5 ),
    .o({\u2_Display/lt39_c6 ,open_n4129}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_6  (
    .a(\u2_Display/n1005 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c6 ),
    .o({\u2_Display/lt39_c7 ,open_n4130}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_7  (
    .a(\u2_Display/n1004 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c7 ),
    .o({\u2_Display/lt39_c8 ,open_n4131}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_8  (
    .a(\u2_Display/n1003 ),
    .b(1'b1),
    .c(\u2_Display/lt39_c8 ),
    .o({\u2_Display/lt39_c9 ,open_n4132}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_9  (
    .a(\u2_Display/n1002 ),
    .b(1'b0),
    .c(\u2_Display/lt39_c9 ),
    .o({\u2_Display/lt39_c10 ,open_n4133}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt39_cin  (
    .a(1'b0),
    .o({\u2_Display/lt39_c0 ,open_n4136}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt39_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt39_c32 ),
    .o({open_n4137,\u2_Display/n1012 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt3_0  (
    .a(\u2_Display/j [0]),
    .b(lcd_ypos[0]),
    .c(\u2_Display/lt3_c0 ),
    .o({\u2_Display/lt3_c1 ,open_n4138}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt3_1  (
    .a(\u2_Display/j [1]),
    .b(lcd_ypos[1]),
    .c(\u2_Display/lt3_c1 ),
    .o({\u2_Display/lt3_c2 ,open_n4139}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt3_10  (
    .a(1'b0),
    .b(lcd_ypos[10]),
    .c(\u2_Display/lt3_c10 ),
    .o({\u2_Display/lt3_c11 ,open_n4140}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt3_11  (
    .a(1'b0),
    .b(lcd_ypos[11]),
    .c(\u2_Display/lt3_c11 ),
    .o({\u2_Display/lt3_c12 ,open_n4141}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt3_2  (
    .a(\u2_Display/j [2]),
    .b(lcd_ypos[2]),
    .c(\u2_Display/lt3_c2 ),
    .o({\u2_Display/lt3_c3 ,open_n4142}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt3_3  (
    .a(\u2_Display/j [3]),
    .b(lcd_ypos[3]),
    .c(\u2_Display/lt3_c3 ),
    .o({\u2_Display/lt3_c4 ,open_n4143}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt3_4  (
    .a(\u2_Display/j [4]),
    .b(lcd_ypos[4]),
    .c(\u2_Display/lt3_c4 ),
    .o({\u2_Display/lt3_c5 ,open_n4144}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt3_5  (
    .a(\u2_Display/j [5]),
    .b(lcd_ypos[5]),
    .c(\u2_Display/lt3_c5 ),
    .o({\u2_Display/lt3_c6 ,open_n4145}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt3_6  (
    .a(\u2_Display/j [6]),
    .b(lcd_ypos[6]),
    .c(\u2_Display/lt3_c6 ),
    .o({\u2_Display/lt3_c7 ,open_n4146}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt3_7  (
    .a(\u2_Display/j [7]),
    .b(lcd_ypos[7]),
    .c(\u2_Display/lt3_c7 ),
    .o({\u2_Display/lt3_c8 ,open_n4147}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt3_8  (
    .a(\u2_Display/j [8]),
    .b(lcd_ypos[8]),
    .c(\u2_Display/lt3_c8 ),
    .o({\u2_Display/lt3_c9 ,open_n4148}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt3_9  (
    .a(\u2_Display/j [9]),
    .b(lcd_ypos[9]),
    .c(\u2_Display/lt3_c9 ),
    .o({\u2_Display/lt3_c10 ,open_n4149}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt3_cin  (
    .a(1'b0),
    .o({\u2_Display/lt3_c0 ,open_n4152}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt3_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt3_c12 ),
    .o({open_n4153,\u2_Display/n50 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_0  (
    .a(\u2_Display/n1046 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c0 ),
    .o({\u2_Display/lt40_c1 ,open_n4154}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_1  (
    .a(\u2_Display/n1045 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c1 ),
    .o({\u2_Display/lt40_c2 ,open_n4155}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_10  (
    .a(\u2_Display/n1036 ),
    .b(1'b1),
    .c(\u2_Display/lt40_c10 ),
    .o({\u2_Display/lt40_c11 ,open_n4156}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_11  (
    .a(\u2_Display/n1035 ),
    .b(1'b1),
    .c(\u2_Display/lt40_c11 ),
    .o({\u2_Display/lt40_c12 ,open_n4157}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_12  (
    .a(\u2_Display/n1034 ),
    .b(1'b1),
    .c(\u2_Display/lt40_c12 ),
    .o({\u2_Display/lt40_c13 ,open_n4158}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_13  (
    .a(\u2_Display/n1033 ),
    .b(1'b1),
    .c(\u2_Display/lt40_c13 ),
    .o({\u2_Display/lt40_c14 ,open_n4159}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_14  (
    .a(\u2_Display/n1032 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c14 ),
    .o({\u2_Display/lt40_c15 ,open_n4160}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_15  (
    .a(\u2_Display/n1031 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c15 ),
    .o({\u2_Display/lt40_c16 ,open_n4161}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_16  (
    .a(\u2_Display/n1030 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c16 ),
    .o({\u2_Display/lt40_c17 ,open_n4162}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_17  (
    .a(\u2_Display/n1029 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c17 ),
    .o({\u2_Display/lt40_c18 ,open_n4163}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_18  (
    .a(\u2_Display/n1028 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c18 ),
    .o({\u2_Display/lt40_c19 ,open_n4164}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_19  (
    .a(\u2_Display/n1027 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c19 ),
    .o({\u2_Display/lt40_c20 ,open_n4165}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_2  (
    .a(\u2_Display/n1044 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c2 ),
    .o({\u2_Display/lt40_c3 ,open_n4166}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_20  (
    .a(\u2_Display/n1026 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c20 ),
    .o({\u2_Display/lt40_c21 ,open_n4167}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_21  (
    .a(\u2_Display/n1025 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c21 ),
    .o({\u2_Display/lt40_c22 ,open_n4168}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_22  (
    .a(\u2_Display/n1024 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c22 ),
    .o({\u2_Display/lt40_c23 ,open_n4169}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_23  (
    .a(\u2_Display/n1023 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c23 ),
    .o({\u2_Display/lt40_c24 ,open_n4170}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_24  (
    .a(\u2_Display/n1022 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c24 ),
    .o({\u2_Display/lt40_c25 ,open_n4171}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_25  (
    .a(\u2_Display/n1021 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c25 ),
    .o({\u2_Display/lt40_c26 ,open_n4172}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_26  (
    .a(\u2_Display/n1020 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c26 ),
    .o({\u2_Display/lt40_c27 ,open_n4173}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_27  (
    .a(\u2_Display/n1019 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c27 ),
    .o({\u2_Display/lt40_c28 ,open_n4174}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_28  (
    .a(\u2_Display/n1018 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c28 ),
    .o({\u2_Display/lt40_c29 ,open_n4175}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_29  (
    .a(\u2_Display/n1017 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c29 ),
    .o({\u2_Display/lt40_c30 ,open_n4176}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_3  (
    .a(\u2_Display/n1043 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c3 ),
    .o({\u2_Display/lt40_c4 ,open_n4177}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_30  (
    .a(\u2_Display/n1016 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c30 ),
    .o({\u2_Display/lt40_c31 ,open_n4178}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_31  (
    .a(\u2_Display/n1015 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c31 ),
    .o({\u2_Display/lt40_c32 ,open_n4179}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_4  (
    .a(\u2_Display/n1042 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c4 ),
    .o({\u2_Display/lt40_c5 ,open_n4180}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_5  (
    .a(\u2_Display/n1041 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c5 ),
    .o({\u2_Display/lt40_c6 ,open_n4181}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_6  (
    .a(\u2_Display/n1040 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c6 ),
    .o({\u2_Display/lt40_c7 ,open_n4182}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_7  (
    .a(\u2_Display/n1039 ),
    .b(1'b1),
    .c(\u2_Display/lt40_c7 ),
    .o({\u2_Display/lt40_c8 ,open_n4183}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_8  (
    .a(\u2_Display/n1038 ),
    .b(1'b0),
    .c(\u2_Display/lt40_c8 ),
    .o({\u2_Display/lt40_c9 ,open_n4184}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_9  (
    .a(\u2_Display/n1037 ),
    .b(1'b1),
    .c(\u2_Display/lt40_c9 ),
    .o({\u2_Display/lt40_c10 ,open_n4185}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt40_cin  (
    .a(1'b0),
    .o({\u2_Display/lt40_c0 ,open_n4188}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt40_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt40_c32 ),
    .o({open_n4189,\u2_Display/n1047 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_0  (
    .a(\u2_Display/n1081 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c0 ),
    .o({\u2_Display/lt41_c1 ,open_n4190}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_1  (
    .a(\u2_Display/n1080 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c1 ),
    .o({\u2_Display/lt41_c2 ,open_n4191}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_10  (
    .a(\u2_Display/n1071 ),
    .b(1'b1),
    .c(\u2_Display/lt41_c10 ),
    .o({\u2_Display/lt41_c11 ,open_n4192}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_11  (
    .a(\u2_Display/n1070 ),
    .b(1'b1),
    .c(\u2_Display/lt41_c11 ),
    .o({\u2_Display/lt41_c12 ,open_n4193}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_12  (
    .a(\u2_Display/n1069 ),
    .b(1'b1),
    .c(\u2_Display/lt41_c12 ),
    .o({\u2_Display/lt41_c13 ,open_n4194}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_13  (
    .a(\u2_Display/n1068 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c13 ),
    .o({\u2_Display/lt41_c14 ,open_n4195}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_14  (
    .a(\u2_Display/n1067 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c14 ),
    .o({\u2_Display/lt41_c15 ,open_n4196}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_15  (
    .a(\u2_Display/n1066 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c15 ),
    .o({\u2_Display/lt41_c16 ,open_n4197}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_16  (
    .a(\u2_Display/n1065 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c16 ),
    .o({\u2_Display/lt41_c17 ,open_n4198}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_17  (
    .a(\u2_Display/n1064 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c17 ),
    .o({\u2_Display/lt41_c18 ,open_n4199}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_18  (
    .a(\u2_Display/n1063 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c18 ),
    .o({\u2_Display/lt41_c19 ,open_n4200}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_19  (
    .a(\u2_Display/n1062 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c19 ),
    .o({\u2_Display/lt41_c20 ,open_n4201}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_2  (
    .a(\u2_Display/n1079 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c2 ),
    .o({\u2_Display/lt41_c3 ,open_n4202}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_20  (
    .a(\u2_Display/n1061 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c20 ),
    .o({\u2_Display/lt41_c21 ,open_n4203}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_21  (
    .a(\u2_Display/n1060 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c21 ),
    .o({\u2_Display/lt41_c22 ,open_n4204}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_22  (
    .a(\u2_Display/n1059 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c22 ),
    .o({\u2_Display/lt41_c23 ,open_n4205}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_23  (
    .a(\u2_Display/n1058 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c23 ),
    .o({\u2_Display/lt41_c24 ,open_n4206}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_24  (
    .a(\u2_Display/n1057 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c24 ),
    .o({\u2_Display/lt41_c25 ,open_n4207}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_25  (
    .a(\u2_Display/n1056 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c25 ),
    .o({\u2_Display/lt41_c26 ,open_n4208}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_26  (
    .a(\u2_Display/n1055 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c26 ),
    .o({\u2_Display/lt41_c27 ,open_n4209}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_27  (
    .a(\u2_Display/n1054 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c27 ),
    .o({\u2_Display/lt41_c28 ,open_n4210}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_28  (
    .a(\u2_Display/n1053 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c28 ),
    .o({\u2_Display/lt41_c29 ,open_n4211}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_29  (
    .a(\u2_Display/n1052 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c29 ),
    .o({\u2_Display/lt41_c30 ,open_n4212}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_3  (
    .a(\u2_Display/n1078 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c3 ),
    .o({\u2_Display/lt41_c4 ,open_n4213}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_30  (
    .a(\u2_Display/n1051 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c30 ),
    .o({\u2_Display/lt41_c31 ,open_n4214}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_31  (
    .a(\u2_Display/n1050 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c31 ),
    .o({\u2_Display/lt41_c32 ,open_n4215}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_4  (
    .a(\u2_Display/n1077 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c4 ),
    .o({\u2_Display/lt41_c5 ,open_n4216}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_5  (
    .a(\u2_Display/n1076 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c5 ),
    .o({\u2_Display/lt41_c6 ,open_n4217}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_6  (
    .a(\u2_Display/n1075 ),
    .b(1'b1),
    .c(\u2_Display/lt41_c6 ),
    .o({\u2_Display/lt41_c7 ,open_n4218}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_7  (
    .a(\u2_Display/n1074 ),
    .b(1'b0),
    .c(\u2_Display/lt41_c7 ),
    .o({\u2_Display/lt41_c8 ,open_n4219}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_8  (
    .a(\u2_Display/n1073 ),
    .b(1'b1),
    .c(\u2_Display/lt41_c8 ),
    .o({\u2_Display/lt41_c9 ,open_n4220}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_9  (
    .a(\u2_Display/n1072 ),
    .b(1'b1),
    .c(\u2_Display/lt41_c9 ),
    .o({\u2_Display/lt41_c10 ,open_n4221}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt41_cin  (
    .a(1'b0),
    .o({\u2_Display/lt41_c0 ,open_n4224}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt41_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt41_c32 ),
    .o({open_n4225,\u2_Display/n1082 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_0  (
    .a(\u2_Display/n1116 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c0 ),
    .o({\u2_Display/lt42_c1 ,open_n4226}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_1  (
    .a(\u2_Display/n1115 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c1 ),
    .o({\u2_Display/lt42_c2 ,open_n4227}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_10  (
    .a(\u2_Display/n1106 ),
    .b(1'b1),
    .c(\u2_Display/lt42_c10 ),
    .o({\u2_Display/lt42_c11 ,open_n4228}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_11  (
    .a(\u2_Display/n1105 ),
    .b(1'b1),
    .c(\u2_Display/lt42_c11 ),
    .o({\u2_Display/lt42_c12 ,open_n4229}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_12  (
    .a(\u2_Display/n1104 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c12 ),
    .o({\u2_Display/lt42_c13 ,open_n4230}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_13  (
    .a(\u2_Display/n1103 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c13 ),
    .o({\u2_Display/lt42_c14 ,open_n4231}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_14  (
    .a(\u2_Display/n1102 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c14 ),
    .o({\u2_Display/lt42_c15 ,open_n4232}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_15  (
    .a(\u2_Display/n1101 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c15 ),
    .o({\u2_Display/lt42_c16 ,open_n4233}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_16  (
    .a(\u2_Display/n1100 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c16 ),
    .o({\u2_Display/lt42_c17 ,open_n4234}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_17  (
    .a(\u2_Display/n1099 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c17 ),
    .o({\u2_Display/lt42_c18 ,open_n4235}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_18  (
    .a(\u2_Display/n1098 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c18 ),
    .o({\u2_Display/lt42_c19 ,open_n4236}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_19  (
    .a(\u2_Display/n1097 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c19 ),
    .o({\u2_Display/lt42_c20 ,open_n4237}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_2  (
    .a(\u2_Display/n1114 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c2 ),
    .o({\u2_Display/lt42_c3 ,open_n4238}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_20  (
    .a(\u2_Display/n1096 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c20 ),
    .o({\u2_Display/lt42_c21 ,open_n4239}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_21  (
    .a(\u2_Display/n1095 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c21 ),
    .o({\u2_Display/lt42_c22 ,open_n4240}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_22  (
    .a(\u2_Display/n1094 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c22 ),
    .o({\u2_Display/lt42_c23 ,open_n4241}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_23  (
    .a(\u2_Display/n1093 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c23 ),
    .o({\u2_Display/lt42_c24 ,open_n4242}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_24  (
    .a(\u2_Display/n1092 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c24 ),
    .o({\u2_Display/lt42_c25 ,open_n4243}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_25  (
    .a(\u2_Display/n1091 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c25 ),
    .o({\u2_Display/lt42_c26 ,open_n4244}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_26  (
    .a(\u2_Display/n1090 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c26 ),
    .o({\u2_Display/lt42_c27 ,open_n4245}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_27  (
    .a(\u2_Display/n1089 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c27 ),
    .o({\u2_Display/lt42_c28 ,open_n4246}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_28  (
    .a(\u2_Display/n1088 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c28 ),
    .o({\u2_Display/lt42_c29 ,open_n4247}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_29  (
    .a(\u2_Display/n1087 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c29 ),
    .o({\u2_Display/lt42_c30 ,open_n4248}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_3  (
    .a(\u2_Display/n1113 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c3 ),
    .o({\u2_Display/lt42_c4 ,open_n4249}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_30  (
    .a(\u2_Display/n1086 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c30 ),
    .o({\u2_Display/lt42_c31 ,open_n4250}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_31  (
    .a(\u2_Display/n1085 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c31 ),
    .o({\u2_Display/lt42_c32 ,open_n4251}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_4  (
    .a(\u2_Display/n1112 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c4 ),
    .o({\u2_Display/lt42_c5 ,open_n4252}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_5  (
    .a(\u2_Display/n1111 ),
    .b(1'b1),
    .c(\u2_Display/lt42_c5 ),
    .o({\u2_Display/lt42_c6 ,open_n4253}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_6  (
    .a(\u2_Display/n1110 ),
    .b(1'b0),
    .c(\u2_Display/lt42_c6 ),
    .o({\u2_Display/lt42_c7 ,open_n4254}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_7  (
    .a(\u2_Display/n1109 ),
    .b(1'b1),
    .c(\u2_Display/lt42_c7 ),
    .o({\u2_Display/lt42_c8 ,open_n4255}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_8  (
    .a(\u2_Display/n1108 ),
    .b(1'b1),
    .c(\u2_Display/lt42_c8 ),
    .o({\u2_Display/lt42_c9 ,open_n4256}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_9  (
    .a(\u2_Display/n1107 ),
    .b(1'b1),
    .c(\u2_Display/lt42_c9 ),
    .o({\u2_Display/lt42_c10 ,open_n4257}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt42_cin  (
    .a(1'b0),
    .o({\u2_Display/lt42_c0 ,open_n4260}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt42_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt42_c32 ),
    .o({open_n4261,\u2_Display/n1117 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_0  (
    .a(\u2_Display/n1151 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c0 ),
    .o({\u2_Display/lt43_c1 ,open_n4262}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_1  (
    .a(\u2_Display/n1150 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c1 ),
    .o({\u2_Display/lt43_c2 ,open_n4263}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_10  (
    .a(\u2_Display/n1141 ),
    .b(1'b1),
    .c(\u2_Display/lt43_c10 ),
    .o({\u2_Display/lt43_c11 ,open_n4264}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_11  (
    .a(\u2_Display/n1140 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c11 ),
    .o({\u2_Display/lt43_c12 ,open_n4265}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_12  (
    .a(\u2_Display/n1139 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c12 ),
    .o({\u2_Display/lt43_c13 ,open_n4266}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_13  (
    .a(\u2_Display/n1138 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c13 ),
    .o({\u2_Display/lt43_c14 ,open_n4267}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_14  (
    .a(\u2_Display/n1137 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c14 ),
    .o({\u2_Display/lt43_c15 ,open_n4268}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_15  (
    .a(\u2_Display/n1136 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c15 ),
    .o({\u2_Display/lt43_c16 ,open_n4269}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_16  (
    .a(\u2_Display/n1135 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c16 ),
    .o({\u2_Display/lt43_c17 ,open_n4270}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_17  (
    .a(\u2_Display/n1134 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c17 ),
    .o({\u2_Display/lt43_c18 ,open_n4271}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_18  (
    .a(\u2_Display/n1133 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c18 ),
    .o({\u2_Display/lt43_c19 ,open_n4272}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_19  (
    .a(\u2_Display/n1132 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c19 ),
    .o({\u2_Display/lt43_c20 ,open_n4273}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_2  (
    .a(\u2_Display/n1149 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c2 ),
    .o({\u2_Display/lt43_c3 ,open_n4274}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_20  (
    .a(\u2_Display/n1131 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c20 ),
    .o({\u2_Display/lt43_c21 ,open_n4275}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_21  (
    .a(\u2_Display/n1130 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c21 ),
    .o({\u2_Display/lt43_c22 ,open_n4276}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_22  (
    .a(\u2_Display/n1129 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c22 ),
    .o({\u2_Display/lt43_c23 ,open_n4277}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_23  (
    .a(\u2_Display/n1128 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c23 ),
    .o({\u2_Display/lt43_c24 ,open_n4278}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_24  (
    .a(\u2_Display/n1127 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c24 ),
    .o({\u2_Display/lt43_c25 ,open_n4279}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_25  (
    .a(\u2_Display/n1126 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c25 ),
    .o({\u2_Display/lt43_c26 ,open_n4280}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_26  (
    .a(\u2_Display/n1125 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c26 ),
    .o({\u2_Display/lt43_c27 ,open_n4281}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_27  (
    .a(\u2_Display/n1124 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c27 ),
    .o({\u2_Display/lt43_c28 ,open_n4282}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_28  (
    .a(\u2_Display/n1123 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c28 ),
    .o({\u2_Display/lt43_c29 ,open_n4283}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_29  (
    .a(\u2_Display/n1122 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c29 ),
    .o({\u2_Display/lt43_c30 ,open_n4284}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_3  (
    .a(\u2_Display/n1148 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c3 ),
    .o({\u2_Display/lt43_c4 ,open_n4285}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_30  (
    .a(\u2_Display/n1121 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c30 ),
    .o({\u2_Display/lt43_c31 ,open_n4286}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_31  (
    .a(\u2_Display/n1120 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c31 ),
    .o({\u2_Display/lt43_c32 ,open_n4287}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_4  (
    .a(\u2_Display/n1147 ),
    .b(1'b1),
    .c(\u2_Display/lt43_c4 ),
    .o({\u2_Display/lt43_c5 ,open_n4288}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_5  (
    .a(\u2_Display/n1146 ),
    .b(1'b0),
    .c(\u2_Display/lt43_c5 ),
    .o({\u2_Display/lt43_c6 ,open_n4289}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_6  (
    .a(\u2_Display/n1145 ),
    .b(1'b1),
    .c(\u2_Display/lt43_c6 ),
    .o({\u2_Display/lt43_c7 ,open_n4290}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_7  (
    .a(\u2_Display/n1144 ),
    .b(1'b1),
    .c(\u2_Display/lt43_c7 ),
    .o({\u2_Display/lt43_c8 ,open_n4291}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_8  (
    .a(\u2_Display/n1143 ),
    .b(1'b1),
    .c(\u2_Display/lt43_c8 ),
    .o({\u2_Display/lt43_c9 ,open_n4292}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_9  (
    .a(\u2_Display/n1142 ),
    .b(1'b1),
    .c(\u2_Display/lt43_c9 ),
    .o({\u2_Display/lt43_c10 ,open_n4293}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt43_cin  (
    .a(1'b0),
    .o({\u2_Display/lt43_c0 ,open_n4296}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt43_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt43_c32 ),
    .o({open_n4297,\u2_Display/n1152 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_0  (
    .a(\u2_Display/n1186 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c0 ),
    .o({\u2_Display/lt44_c1 ,open_n4298}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_1  (
    .a(\u2_Display/n1185 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c1 ),
    .o({\u2_Display/lt44_c2 ,open_n4299}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_10  (
    .a(\u2_Display/n1176 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c10 ),
    .o({\u2_Display/lt44_c11 ,open_n4300}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_11  (
    .a(\u2_Display/n1175 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c11 ),
    .o({\u2_Display/lt44_c12 ,open_n4301}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_12  (
    .a(\u2_Display/n1174 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c12 ),
    .o({\u2_Display/lt44_c13 ,open_n4302}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_13  (
    .a(\u2_Display/n1173 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c13 ),
    .o({\u2_Display/lt44_c14 ,open_n4303}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_14  (
    .a(\u2_Display/n1172 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c14 ),
    .o({\u2_Display/lt44_c15 ,open_n4304}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_15  (
    .a(\u2_Display/n1171 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c15 ),
    .o({\u2_Display/lt44_c16 ,open_n4305}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_16  (
    .a(\u2_Display/n1170 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c16 ),
    .o({\u2_Display/lt44_c17 ,open_n4306}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_17  (
    .a(\u2_Display/n1169 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c17 ),
    .o({\u2_Display/lt44_c18 ,open_n4307}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_18  (
    .a(\u2_Display/n1168 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c18 ),
    .o({\u2_Display/lt44_c19 ,open_n4308}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_19  (
    .a(\u2_Display/n1167 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c19 ),
    .o({\u2_Display/lt44_c20 ,open_n4309}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_2  (
    .a(\u2_Display/n1184 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c2 ),
    .o({\u2_Display/lt44_c3 ,open_n4310}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_20  (
    .a(\u2_Display/n1166 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c20 ),
    .o({\u2_Display/lt44_c21 ,open_n4311}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_21  (
    .a(\u2_Display/n1165 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c21 ),
    .o({\u2_Display/lt44_c22 ,open_n4312}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_22  (
    .a(\u2_Display/n1164 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c22 ),
    .o({\u2_Display/lt44_c23 ,open_n4313}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_23  (
    .a(\u2_Display/n1163 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c23 ),
    .o({\u2_Display/lt44_c24 ,open_n4314}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_24  (
    .a(\u2_Display/n1162 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c24 ),
    .o({\u2_Display/lt44_c25 ,open_n4315}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_25  (
    .a(\u2_Display/n1161 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c25 ),
    .o({\u2_Display/lt44_c26 ,open_n4316}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_26  (
    .a(\u2_Display/n1160 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c26 ),
    .o({\u2_Display/lt44_c27 ,open_n4317}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_27  (
    .a(\u2_Display/n1159 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c27 ),
    .o({\u2_Display/lt44_c28 ,open_n4318}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_28  (
    .a(\u2_Display/n1158 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c28 ),
    .o({\u2_Display/lt44_c29 ,open_n4319}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_29  (
    .a(\u2_Display/n1157 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c29 ),
    .o({\u2_Display/lt44_c30 ,open_n4320}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_3  (
    .a(\u2_Display/n1183 ),
    .b(1'b1),
    .c(\u2_Display/lt44_c3 ),
    .o({\u2_Display/lt44_c4 ,open_n4321}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_30  (
    .a(\u2_Display/n1156 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c30 ),
    .o({\u2_Display/lt44_c31 ,open_n4322}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_31  (
    .a(\u2_Display/n1155 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c31 ),
    .o({\u2_Display/lt44_c32 ,open_n4323}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_4  (
    .a(\u2_Display/n1182 ),
    .b(1'b0),
    .c(\u2_Display/lt44_c4 ),
    .o({\u2_Display/lt44_c5 ,open_n4324}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_5  (
    .a(\u2_Display/n1181 ),
    .b(1'b1),
    .c(\u2_Display/lt44_c5 ),
    .o({\u2_Display/lt44_c6 ,open_n4325}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_6  (
    .a(\u2_Display/n1180 ),
    .b(1'b1),
    .c(\u2_Display/lt44_c6 ),
    .o({\u2_Display/lt44_c7 ,open_n4326}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_7  (
    .a(\u2_Display/n1179 ),
    .b(1'b1),
    .c(\u2_Display/lt44_c7 ),
    .o({\u2_Display/lt44_c8 ,open_n4327}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_8  (
    .a(\u2_Display/n1178 ),
    .b(1'b1),
    .c(\u2_Display/lt44_c8 ),
    .o({\u2_Display/lt44_c9 ,open_n4328}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_9  (
    .a(\u2_Display/n1177 ),
    .b(1'b1),
    .c(\u2_Display/lt44_c9 ),
    .o({\u2_Display/lt44_c10 ,open_n4329}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt44_cin  (
    .a(1'b0),
    .o({\u2_Display/lt44_c0 ,open_n4332}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt44_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt44_c32 ),
    .o({open_n4333,\u2_Display/n1187 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt4_2_0  (
    .a(lcd_xpos[0]),
    .b(\u2_Display/i [0]),
    .c(\u2_Display/lt4_2_c0 ),
    .o({\u2_Display/lt4_2_c1 ,open_n4334}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt4_2_1  (
    .a(lcd_xpos[1]),
    .b(\u2_Display/i [1]),
    .c(\u2_Display/lt4_2_c1 ),
    .o({\u2_Display/lt4_2_c2 ,open_n4335}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt4_2_10  (
    .a(lcd_xpos[10]),
    .b(\u2_Display/n94 [3]),
    .c(\u2_Display/lt4_2_c10 ),
    .o({\u2_Display/lt4_2_c11 ,open_n4336}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt4_2_11  (
    .a(lcd_xpos[11]),
    .b(\u2_Display/add4_2_co ),
    .c(\u2_Display/lt4_2_c11 ),
    .o({\u2_Display/lt4_2_c12 ,open_n4337}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt4_2_2  (
    .a(lcd_xpos[2]),
    .b(\u2_Display/i [2]),
    .c(\u2_Display/lt4_2_c2 ),
    .o({\u2_Display/lt4_2_c3 ,open_n4338}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt4_2_3  (
    .a(lcd_xpos[3]),
    .b(\u2_Display/i [3]),
    .c(\u2_Display/lt4_2_c3 ),
    .o({\u2_Display/lt4_2_c4 ,open_n4339}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt4_2_4  (
    .a(lcd_xpos[4]),
    .b(\u2_Display/i [4]),
    .c(\u2_Display/lt4_2_c4 ),
    .o({\u2_Display/lt4_2_c5 ,open_n4340}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt4_2_5  (
    .a(lcd_xpos[5]),
    .b(\u2_Display/i [5]),
    .c(\u2_Display/lt4_2_c5 ),
    .o({\u2_Display/lt4_2_c6 ,open_n4341}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt4_2_6  (
    .a(lcd_xpos[6]),
    .b(\u2_Display/i [6]),
    .c(\u2_Display/lt4_2_c6 ),
    .o({\u2_Display/lt4_2_c7 ,open_n4342}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt4_2_7  (
    .a(lcd_xpos[7]),
    .b(\u2_Display/n94 [0]),
    .c(\u2_Display/lt4_2_c7 ),
    .o({\u2_Display/lt4_2_c8 ,open_n4343}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt4_2_8  (
    .a(lcd_xpos[8]),
    .b(\u2_Display/n94 [1]),
    .c(\u2_Display/lt4_2_c8 ),
    .o({\u2_Display/lt4_2_c9 ,open_n4344}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt4_2_9  (
    .a(lcd_xpos[9]),
    .b(\u2_Display/n94 [2]),
    .c(\u2_Display/lt4_2_c9 ),
    .o({\u2_Display/lt4_2_c10 ,open_n4345}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt4_2_cin  (
    .a(1'b0),
    .o({\u2_Display/lt4_2_c0 ,open_n4348}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt4_2_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt4_2_c12 ),
    .o({open_n4349,\u2_Display/n95 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_0  (
    .a(\u2_Display/counta [0]),
    .b(1'b0),
    .c(\u2_Display/lt55_c0 ),
    .o({\u2_Display/lt55_c1 ,open_n4350}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_1  (
    .a(\u2_Display/counta [1]),
    .b(1'b0),
    .c(\u2_Display/lt55_c1 ),
    .o({\u2_Display/lt55_c2 ,open_n4351}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_10  (
    .a(\u2_Display/counta [10]),
    .b(1'b0),
    .c(\u2_Display/lt55_c10 ),
    .o({\u2_Display/lt55_c11 ,open_n4352}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_11  (
    .a(\u2_Display/counta [11]),
    .b(1'b0),
    .c(\u2_Display/lt55_c11 ),
    .o({\u2_Display/lt55_c12 ,open_n4353}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_12  (
    .a(\u2_Display/counta [12]),
    .b(1'b0),
    .c(\u2_Display/lt55_c12 ),
    .o({\u2_Display/lt55_c13 ,open_n4354}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_13  (
    .a(\u2_Display/counta [13]),
    .b(1'b0),
    .c(\u2_Display/lt55_c13 ),
    .o({\u2_Display/lt55_c14 ,open_n4355}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_14  (
    .a(\u2_Display/counta [14]),
    .b(1'b0),
    .c(\u2_Display/lt55_c14 ),
    .o({\u2_Display/lt55_c15 ,open_n4356}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_15  (
    .a(\u2_Display/counta [15]),
    .b(1'b0),
    .c(\u2_Display/lt55_c15 ),
    .o({\u2_Display/lt55_c16 ,open_n4357}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_16  (
    .a(\u2_Display/counta [16]),
    .b(1'b0),
    .c(\u2_Display/lt55_c16 ),
    .o({\u2_Display/lt55_c17 ,open_n4358}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_17  (
    .a(\u2_Display/counta [17]),
    .b(1'b0),
    .c(\u2_Display/lt55_c17 ),
    .o({\u2_Display/lt55_c18 ,open_n4359}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_18  (
    .a(\u2_Display/counta [18]),
    .b(1'b0),
    .c(\u2_Display/lt55_c18 ),
    .o({\u2_Display/lt55_c19 ,open_n4360}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_19  (
    .a(\u2_Display/counta [19]),
    .b(1'b0),
    .c(\u2_Display/lt55_c19 ),
    .o({\u2_Display/lt55_c20 ,open_n4361}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_2  (
    .a(\u2_Display/counta [2]),
    .b(1'b0),
    .c(\u2_Display/lt55_c2 ),
    .o({\u2_Display/lt55_c3 ,open_n4362}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_20  (
    .a(\u2_Display/counta [20]),
    .b(1'b0),
    .c(\u2_Display/lt55_c20 ),
    .o({\u2_Display/lt55_c21 ,open_n4363}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_21  (
    .a(\u2_Display/counta [21]),
    .b(1'b0),
    .c(\u2_Display/lt55_c21 ),
    .o({\u2_Display/lt55_c22 ,open_n4364}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_22  (
    .a(\u2_Display/counta [22]),
    .b(1'b0),
    .c(\u2_Display/lt55_c22 ),
    .o({\u2_Display/lt55_c23 ,open_n4365}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_23  (
    .a(\u2_Display/counta [23]),
    .b(1'b0),
    .c(\u2_Display/lt55_c23 ),
    .o({\u2_Display/lt55_c24 ,open_n4366}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_24  (
    .a(\u2_Display/counta [24]),
    .b(1'b1),
    .c(\u2_Display/lt55_c24 ),
    .o({\u2_Display/lt55_c25 ,open_n4367}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_25  (
    .a(\u2_Display/counta [25]),
    .b(1'b0),
    .c(\u2_Display/lt55_c25 ),
    .o({\u2_Display/lt55_c26 ,open_n4368}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_26  (
    .a(\u2_Display/counta [26]),
    .b(1'b0),
    .c(\u2_Display/lt55_c26 ),
    .o({\u2_Display/lt55_c27 ,open_n4369}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_27  (
    .a(\u2_Display/counta [27]),
    .b(1'b0),
    .c(\u2_Display/lt55_c27 ),
    .o({\u2_Display/lt55_c28 ,open_n4370}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_28  (
    .a(\u2_Display/counta [28]),
    .b(1'b0),
    .c(\u2_Display/lt55_c28 ),
    .o({\u2_Display/lt55_c29 ,open_n4371}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_29  (
    .a(\u2_Display/counta [29]),
    .b(1'b1),
    .c(\u2_Display/lt55_c29 ),
    .o({\u2_Display/lt55_c30 ,open_n4372}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_3  (
    .a(\u2_Display/counta [3]),
    .b(1'b0),
    .c(\u2_Display/lt55_c3 ),
    .o({\u2_Display/lt55_c4 ,open_n4373}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_30  (
    .a(\u2_Display/counta [30]),
    .b(1'b1),
    .c(\u2_Display/lt55_c30 ),
    .o({\u2_Display/lt55_c31 ,open_n4374}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_31  (
    .a(\u2_Display/counta [31]),
    .b(1'b1),
    .c(\u2_Display/lt55_c31 ),
    .o({\u2_Display/lt55_c32 ,open_n4375}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_4  (
    .a(\u2_Display/counta [4]),
    .b(1'b0),
    .c(\u2_Display/lt55_c4 ),
    .o({\u2_Display/lt55_c5 ,open_n4376}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_5  (
    .a(\u2_Display/counta [5]),
    .b(1'b0),
    .c(\u2_Display/lt55_c5 ),
    .o({\u2_Display/lt55_c6 ,open_n4377}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_6  (
    .a(\u2_Display/counta [6]),
    .b(1'b0),
    .c(\u2_Display/lt55_c6 ),
    .o({\u2_Display/lt55_c7 ,open_n4378}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_7  (
    .a(\u2_Display/counta [7]),
    .b(1'b0),
    .c(\u2_Display/lt55_c7 ),
    .o({\u2_Display/lt55_c8 ,open_n4379}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_8  (
    .a(\u2_Display/counta [8]),
    .b(1'b0),
    .c(\u2_Display/lt55_c8 ),
    .o({\u2_Display/lt55_c9 ,open_n4380}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_9  (
    .a(\u2_Display/counta [9]),
    .b(1'b0),
    .c(\u2_Display/lt55_c9 ),
    .o({\u2_Display/lt55_c10 ,open_n4381}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt55_cin  (
    .a(1'b0),
    .o({\u2_Display/lt55_c0 ,open_n4384}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt55_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt55_c32 ),
    .o({open_n4385,\u2_Display/n1540 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_0  (
    .a(\u2_Display/n1574 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c0 ),
    .o({\u2_Display/lt56_c1 ,open_n4386}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_1  (
    .a(\u2_Display/n1573 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c1 ),
    .o({\u2_Display/lt56_c2 ,open_n4387}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_10  (
    .a(\u2_Display/n1564 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c10 ),
    .o({\u2_Display/lt56_c11 ,open_n4388}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_11  (
    .a(\u2_Display/n1563 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c11 ),
    .o({\u2_Display/lt56_c12 ,open_n4389}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_12  (
    .a(\u2_Display/n1562 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c12 ),
    .o({\u2_Display/lt56_c13 ,open_n4390}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_13  (
    .a(\u2_Display/n1561 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c13 ),
    .o({\u2_Display/lt56_c14 ,open_n4391}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_14  (
    .a(\u2_Display/n1560 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c14 ),
    .o({\u2_Display/lt56_c15 ,open_n4392}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_15  (
    .a(\u2_Display/n1559 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c15 ),
    .o({\u2_Display/lt56_c16 ,open_n4393}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_16  (
    .a(\u2_Display/n1558 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c16 ),
    .o({\u2_Display/lt56_c17 ,open_n4394}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_17  (
    .a(\u2_Display/n1557 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c17 ),
    .o({\u2_Display/lt56_c18 ,open_n4395}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_18  (
    .a(\u2_Display/n1556 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c18 ),
    .o({\u2_Display/lt56_c19 ,open_n4396}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_19  (
    .a(\u2_Display/n1555 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c19 ),
    .o({\u2_Display/lt56_c20 ,open_n4397}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_2  (
    .a(\u2_Display/n1572 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c2 ),
    .o({\u2_Display/lt56_c3 ,open_n4398}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_20  (
    .a(\u2_Display/n1554 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c20 ),
    .o({\u2_Display/lt56_c21 ,open_n4399}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_21  (
    .a(\u2_Display/n1553 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c21 ),
    .o({\u2_Display/lt56_c22 ,open_n4400}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_22  (
    .a(\u2_Display/n1552 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c22 ),
    .o({\u2_Display/lt56_c23 ,open_n4401}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_23  (
    .a(\u2_Display/n1551 ),
    .b(1'b1),
    .c(\u2_Display/lt56_c23 ),
    .o({\u2_Display/lt56_c24 ,open_n4402}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_24  (
    .a(\u2_Display/n1550 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c24 ),
    .o({\u2_Display/lt56_c25 ,open_n4403}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_25  (
    .a(\u2_Display/n1549 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c25 ),
    .o({\u2_Display/lt56_c26 ,open_n4404}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_26  (
    .a(\u2_Display/n1548 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c26 ),
    .o({\u2_Display/lt56_c27 ,open_n4405}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_27  (
    .a(\u2_Display/n1547 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c27 ),
    .o({\u2_Display/lt56_c28 ,open_n4406}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_28  (
    .a(\u2_Display/n1546 ),
    .b(1'b1),
    .c(\u2_Display/lt56_c28 ),
    .o({\u2_Display/lt56_c29 ,open_n4407}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_29  (
    .a(\u2_Display/n1545 ),
    .b(1'b1),
    .c(\u2_Display/lt56_c29 ),
    .o({\u2_Display/lt56_c30 ,open_n4408}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_3  (
    .a(\u2_Display/n1571 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c3 ),
    .o({\u2_Display/lt56_c4 ,open_n4409}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_30  (
    .a(\u2_Display/n1544 ),
    .b(1'b1),
    .c(\u2_Display/lt56_c30 ),
    .o({\u2_Display/lt56_c31 ,open_n4410}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_31  (
    .a(\u2_Display/n1543 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c31 ),
    .o({\u2_Display/lt56_c32 ,open_n4411}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_4  (
    .a(\u2_Display/n1570 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c4 ),
    .o({\u2_Display/lt56_c5 ,open_n4412}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_5  (
    .a(\u2_Display/n1569 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c5 ),
    .o({\u2_Display/lt56_c6 ,open_n4413}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_6  (
    .a(\u2_Display/n1568 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c6 ),
    .o({\u2_Display/lt56_c7 ,open_n4414}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_7  (
    .a(\u2_Display/n1567 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c7 ),
    .o({\u2_Display/lt56_c8 ,open_n4415}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_8  (
    .a(\u2_Display/n1566 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c8 ),
    .o({\u2_Display/lt56_c9 ,open_n4416}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_9  (
    .a(\u2_Display/n1565 ),
    .b(1'b0),
    .c(\u2_Display/lt56_c9 ),
    .o({\u2_Display/lt56_c10 ,open_n4417}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt56_cin  (
    .a(1'b0),
    .o({\u2_Display/lt56_c0 ,open_n4420}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt56_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt56_c32 ),
    .o({open_n4421,\u2_Display/n1575 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_0  (
    .a(\u2_Display/n1609 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c0 ),
    .o({\u2_Display/lt57_c1 ,open_n4422}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_1  (
    .a(\u2_Display/n1608 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c1 ),
    .o({\u2_Display/lt57_c2 ,open_n4423}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_10  (
    .a(\u2_Display/n1599 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c10 ),
    .o({\u2_Display/lt57_c11 ,open_n4424}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_11  (
    .a(\u2_Display/n1598 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c11 ),
    .o({\u2_Display/lt57_c12 ,open_n4425}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_12  (
    .a(\u2_Display/n1597 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c12 ),
    .o({\u2_Display/lt57_c13 ,open_n4426}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_13  (
    .a(\u2_Display/n1596 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c13 ),
    .o({\u2_Display/lt57_c14 ,open_n4427}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_14  (
    .a(\u2_Display/n1595 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c14 ),
    .o({\u2_Display/lt57_c15 ,open_n4428}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_15  (
    .a(\u2_Display/n1594 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c15 ),
    .o({\u2_Display/lt57_c16 ,open_n4429}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_16  (
    .a(\u2_Display/n1593 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c16 ),
    .o({\u2_Display/lt57_c17 ,open_n4430}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_17  (
    .a(\u2_Display/n1592 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c17 ),
    .o({\u2_Display/lt57_c18 ,open_n4431}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_18  (
    .a(\u2_Display/n1591 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c18 ),
    .o({\u2_Display/lt57_c19 ,open_n4432}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_19  (
    .a(\u2_Display/n1590 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c19 ),
    .o({\u2_Display/lt57_c20 ,open_n4433}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_2  (
    .a(\u2_Display/n1607 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c2 ),
    .o({\u2_Display/lt57_c3 ,open_n4434}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_20  (
    .a(\u2_Display/n1589 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c20 ),
    .o({\u2_Display/lt57_c21 ,open_n4435}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_21  (
    .a(\u2_Display/n1588 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c21 ),
    .o({\u2_Display/lt57_c22 ,open_n4436}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_22  (
    .a(\u2_Display/n1587 ),
    .b(1'b1),
    .c(\u2_Display/lt57_c22 ),
    .o({\u2_Display/lt57_c23 ,open_n4437}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_23  (
    .a(\u2_Display/n1586 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c23 ),
    .o({\u2_Display/lt57_c24 ,open_n4438}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_24  (
    .a(\u2_Display/n1585 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c24 ),
    .o({\u2_Display/lt57_c25 ,open_n4439}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_25  (
    .a(\u2_Display/n1584 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c25 ),
    .o({\u2_Display/lt57_c26 ,open_n4440}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_26  (
    .a(\u2_Display/n1583 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c26 ),
    .o({\u2_Display/lt57_c27 ,open_n4441}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_27  (
    .a(\u2_Display/n1582 ),
    .b(1'b1),
    .c(\u2_Display/lt57_c27 ),
    .o({\u2_Display/lt57_c28 ,open_n4442}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_28  (
    .a(\u2_Display/n1581 ),
    .b(1'b1),
    .c(\u2_Display/lt57_c28 ),
    .o({\u2_Display/lt57_c29 ,open_n4443}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_29  (
    .a(\u2_Display/n1580 ),
    .b(1'b1),
    .c(\u2_Display/lt57_c29 ),
    .o({\u2_Display/lt57_c30 ,open_n4444}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_3  (
    .a(\u2_Display/n1606 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c3 ),
    .o({\u2_Display/lt57_c4 ,open_n4445}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_30  (
    .a(\u2_Display/n1579 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c30 ),
    .o({\u2_Display/lt57_c31 ,open_n4446}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_31  (
    .a(\u2_Display/n1578 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c31 ),
    .o({\u2_Display/lt57_c32 ,open_n4447}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_4  (
    .a(\u2_Display/n1605 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c4 ),
    .o({\u2_Display/lt57_c5 ,open_n4448}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_5  (
    .a(\u2_Display/n1604 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c5 ),
    .o({\u2_Display/lt57_c6 ,open_n4449}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_6  (
    .a(\u2_Display/n1603 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c6 ),
    .o({\u2_Display/lt57_c7 ,open_n4450}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_7  (
    .a(\u2_Display/n1602 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c7 ),
    .o({\u2_Display/lt57_c8 ,open_n4451}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_8  (
    .a(\u2_Display/n1601 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c8 ),
    .o({\u2_Display/lt57_c9 ,open_n4452}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_9  (
    .a(\u2_Display/n1600 ),
    .b(1'b0),
    .c(\u2_Display/lt57_c9 ),
    .o({\u2_Display/lt57_c10 ,open_n4453}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt57_cin  (
    .a(1'b0),
    .o({\u2_Display/lt57_c0 ,open_n4456}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt57_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt57_c32 ),
    .o({open_n4457,\u2_Display/n1610 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_0  (
    .a(\u2_Display/n1644 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c0 ),
    .o({\u2_Display/lt58_c1 ,open_n4458}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_1  (
    .a(\u2_Display/n1643 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c1 ),
    .o({\u2_Display/lt58_c2 ,open_n4459}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_10  (
    .a(\u2_Display/n1634 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c10 ),
    .o({\u2_Display/lt58_c11 ,open_n4460}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_11  (
    .a(\u2_Display/n1633 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c11 ),
    .o({\u2_Display/lt58_c12 ,open_n4461}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_12  (
    .a(\u2_Display/n1632 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c12 ),
    .o({\u2_Display/lt58_c13 ,open_n4462}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_13  (
    .a(\u2_Display/n1631 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c13 ),
    .o({\u2_Display/lt58_c14 ,open_n4463}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_14  (
    .a(\u2_Display/n1630 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c14 ),
    .o({\u2_Display/lt58_c15 ,open_n4464}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_15  (
    .a(\u2_Display/n1629 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c15 ),
    .o({\u2_Display/lt58_c16 ,open_n4465}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_16  (
    .a(\u2_Display/n1628 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c16 ),
    .o({\u2_Display/lt58_c17 ,open_n4466}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_17  (
    .a(\u2_Display/n1627 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c17 ),
    .o({\u2_Display/lt58_c18 ,open_n4467}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_18  (
    .a(\u2_Display/n1626 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c18 ),
    .o({\u2_Display/lt58_c19 ,open_n4468}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_19  (
    .a(\u2_Display/n1625 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c19 ),
    .o({\u2_Display/lt58_c20 ,open_n4469}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_2  (
    .a(\u2_Display/n1642 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c2 ),
    .o({\u2_Display/lt58_c3 ,open_n4470}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_20  (
    .a(\u2_Display/n1624 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c20 ),
    .o({\u2_Display/lt58_c21 ,open_n4471}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_21  (
    .a(\u2_Display/n1623 ),
    .b(1'b1),
    .c(\u2_Display/lt58_c21 ),
    .o({\u2_Display/lt58_c22 ,open_n4472}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_22  (
    .a(\u2_Display/n1622 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c22 ),
    .o({\u2_Display/lt58_c23 ,open_n4473}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_23  (
    .a(\u2_Display/n1621 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c23 ),
    .o({\u2_Display/lt58_c24 ,open_n4474}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_24  (
    .a(\u2_Display/n1620 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c24 ),
    .o({\u2_Display/lt58_c25 ,open_n4475}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_25  (
    .a(\u2_Display/n1619 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c25 ),
    .o({\u2_Display/lt58_c26 ,open_n4476}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_26  (
    .a(\u2_Display/n1618 ),
    .b(1'b1),
    .c(\u2_Display/lt58_c26 ),
    .o({\u2_Display/lt58_c27 ,open_n4477}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_27  (
    .a(\u2_Display/n1617 ),
    .b(1'b1),
    .c(\u2_Display/lt58_c27 ),
    .o({\u2_Display/lt58_c28 ,open_n4478}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_28  (
    .a(\u2_Display/n1616 ),
    .b(1'b1),
    .c(\u2_Display/lt58_c28 ),
    .o({\u2_Display/lt58_c29 ,open_n4479}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_29  (
    .a(\u2_Display/n1615 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c29 ),
    .o({\u2_Display/lt58_c30 ,open_n4480}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_3  (
    .a(\u2_Display/n1641 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c3 ),
    .o({\u2_Display/lt58_c4 ,open_n4481}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_30  (
    .a(\u2_Display/n1614 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c30 ),
    .o({\u2_Display/lt58_c31 ,open_n4482}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_31  (
    .a(\u2_Display/n1613 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c31 ),
    .o({\u2_Display/lt58_c32 ,open_n4483}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_4  (
    .a(\u2_Display/n1640 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c4 ),
    .o({\u2_Display/lt58_c5 ,open_n4484}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_5  (
    .a(\u2_Display/n1639 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c5 ),
    .o({\u2_Display/lt58_c6 ,open_n4485}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_6  (
    .a(\u2_Display/n1638 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c6 ),
    .o({\u2_Display/lt58_c7 ,open_n4486}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_7  (
    .a(\u2_Display/n1637 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c7 ),
    .o({\u2_Display/lt58_c8 ,open_n4487}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_8  (
    .a(\u2_Display/n1636 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c8 ),
    .o({\u2_Display/lt58_c9 ,open_n4488}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_9  (
    .a(\u2_Display/n1635 ),
    .b(1'b0),
    .c(\u2_Display/lt58_c9 ),
    .o({\u2_Display/lt58_c10 ,open_n4489}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt58_cin  (
    .a(1'b0),
    .o({\u2_Display/lt58_c0 ,open_n4492}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt58_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt58_c32 ),
    .o({open_n4493,\u2_Display/n1645 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_0  (
    .a(\u2_Display/n1679 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c0 ),
    .o({\u2_Display/lt59_c1 ,open_n4494}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_1  (
    .a(\u2_Display/n1678 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c1 ),
    .o({\u2_Display/lt59_c2 ,open_n4495}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_10  (
    .a(\u2_Display/n1669 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c10 ),
    .o({\u2_Display/lt59_c11 ,open_n4496}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_11  (
    .a(\u2_Display/n1668 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c11 ),
    .o({\u2_Display/lt59_c12 ,open_n4497}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_12  (
    .a(\u2_Display/n1667 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c12 ),
    .o({\u2_Display/lt59_c13 ,open_n4498}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_13  (
    .a(\u2_Display/n1666 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c13 ),
    .o({\u2_Display/lt59_c14 ,open_n4499}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_14  (
    .a(\u2_Display/n1665 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c14 ),
    .o({\u2_Display/lt59_c15 ,open_n4500}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_15  (
    .a(\u2_Display/n1664 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c15 ),
    .o({\u2_Display/lt59_c16 ,open_n4501}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_16  (
    .a(\u2_Display/n1663 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c16 ),
    .o({\u2_Display/lt59_c17 ,open_n4502}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_17  (
    .a(\u2_Display/n1662 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c17 ),
    .o({\u2_Display/lt59_c18 ,open_n4503}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_18  (
    .a(\u2_Display/n1661 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c18 ),
    .o({\u2_Display/lt59_c19 ,open_n4504}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_19  (
    .a(\u2_Display/n1660 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c19 ),
    .o({\u2_Display/lt59_c20 ,open_n4505}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_2  (
    .a(\u2_Display/n1677 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c2 ),
    .o({\u2_Display/lt59_c3 ,open_n4506}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_20  (
    .a(\u2_Display/n1659 ),
    .b(1'b1),
    .c(\u2_Display/lt59_c20 ),
    .o({\u2_Display/lt59_c21 ,open_n4507}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_21  (
    .a(\u2_Display/n1658 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c21 ),
    .o({\u2_Display/lt59_c22 ,open_n4508}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_22  (
    .a(\u2_Display/n1657 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c22 ),
    .o({\u2_Display/lt59_c23 ,open_n4509}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_23  (
    .a(\u2_Display/n1656 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c23 ),
    .o({\u2_Display/lt59_c24 ,open_n4510}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_24  (
    .a(\u2_Display/n1655 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c24 ),
    .o({\u2_Display/lt59_c25 ,open_n4511}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_25  (
    .a(\u2_Display/n1654 ),
    .b(1'b1),
    .c(\u2_Display/lt59_c25 ),
    .o({\u2_Display/lt59_c26 ,open_n4512}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_26  (
    .a(\u2_Display/n1653 ),
    .b(1'b1),
    .c(\u2_Display/lt59_c26 ),
    .o({\u2_Display/lt59_c27 ,open_n4513}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_27  (
    .a(\u2_Display/n1652 ),
    .b(1'b1),
    .c(\u2_Display/lt59_c27 ),
    .o({\u2_Display/lt59_c28 ,open_n4514}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_28  (
    .a(\u2_Display/n1651 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c28 ),
    .o({\u2_Display/lt59_c29 ,open_n4515}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_29  (
    .a(\u2_Display/n1650 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c29 ),
    .o({\u2_Display/lt59_c30 ,open_n4516}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_3  (
    .a(\u2_Display/n1676 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c3 ),
    .o({\u2_Display/lt59_c4 ,open_n4517}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_30  (
    .a(\u2_Display/n1649 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c30 ),
    .o({\u2_Display/lt59_c31 ,open_n4518}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_31  (
    .a(\u2_Display/n1648 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c31 ),
    .o({\u2_Display/lt59_c32 ,open_n4519}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_4  (
    .a(\u2_Display/n1675 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c4 ),
    .o({\u2_Display/lt59_c5 ,open_n4520}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_5  (
    .a(\u2_Display/n1674 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c5 ),
    .o({\u2_Display/lt59_c6 ,open_n4521}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_6  (
    .a(\u2_Display/n1673 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c6 ),
    .o({\u2_Display/lt59_c7 ,open_n4522}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_7  (
    .a(\u2_Display/n1672 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c7 ),
    .o({\u2_Display/lt59_c8 ,open_n4523}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_8  (
    .a(\u2_Display/n1671 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c8 ),
    .o({\u2_Display/lt59_c9 ,open_n4524}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_9  (
    .a(\u2_Display/n1670 ),
    .b(1'b0),
    .c(\u2_Display/lt59_c9 ),
    .o({\u2_Display/lt59_c10 ,open_n4525}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt59_cin  (
    .a(1'b0),
    .o({\u2_Display/lt59_c0 ,open_n4528}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt59_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt59_c32 ),
    .o({open_n4529,\u2_Display/n1680 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_0  (
    .a(\u2_Display/n96 [0]),
    .b(lcd_xpos[0]),
    .c(\u2_Display/lt5_2_c0 ),
    .o({\u2_Display/lt5_2_c1 ,open_n4530}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_1  (
    .a(\u2_Display/n96 [1]),
    .b(lcd_xpos[1]),
    .c(\u2_Display/lt5_2_c1 ),
    .o({\u2_Display/lt5_2_c2 ,open_n4531}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_10  (
    .a(\u2_Display/n96 [10]),
    .b(lcd_xpos[10]),
    .c(\u2_Display/lt5_2_c10 ),
    .o({\u2_Display/lt5_2_c11 ,open_n4532}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_11  (
    .a(\u2_Display/n96 [31]),
    .b(lcd_xpos[11]),
    .c(\u2_Display/lt5_2_c11 ),
    .o({\u2_Display/lt5_2_c12 ,open_n4533}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_12  (
    .a(\u2_Display/n96 [31]),
    .b(1'b0),
    .c(\u2_Display/lt5_2_c12 ),
    .o({\u2_Display/lt5_2_c13 ,open_n4534}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_2  (
    .a(\u2_Display/n96 [2]),
    .b(lcd_xpos[2]),
    .c(\u2_Display/lt5_2_c2 ),
    .o({\u2_Display/lt5_2_c3 ,open_n4535}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_3  (
    .a(\u2_Display/n96 [3]),
    .b(lcd_xpos[3]),
    .c(\u2_Display/lt5_2_c3 ),
    .o({\u2_Display/lt5_2_c4 ,open_n4536}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_4  (
    .a(\u2_Display/n96 [4]),
    .b(lcd_xpos[4]),
    .c(\u2_Display/lt5_2_c4 ),
    .o({\u2_Display/lt5_2_c5 ,open_n4537}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_5  (
    .a(\u2_Display/n96 [5]),
    .b(lcd_xpos[5]),
    .c(\u2_Display/lt5_2_c5 ),
    .o({\u2_Display/lt5_2_c6 ,open_n4538}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_6  (
    .a(\u2_Display/n96 [6]),
    .b(lcd_xpos[6]),
    .c(\u2_Display/lt5_2_c6 ),
    .o({\u2_Display/lt5_2_c7 ,open_n4539}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_7  (
    .a(\u2_Display/n96 [7]),
    .b(lcd_xpos[7]),
    .c(\u2_Display/lt5_2_c7 ),
    .o({\u2_Display/lt5_2_c8 ,open_n4540}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_8  (
    .a(\u2_Display/n96 [8]),
    .b(lcd_xpos[8]),
    .c(\u2_Display/lt5_2_c8 ),
    .o({\u2_Display/lt5_2_c9 ,open_n4541}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_9  (
    .a(\u2_Display/n96 [9]),
    .b(lcd_xpos[9]),
    .c(\u2_Display/lt5_2_c9 ),
    .o({\u2_Display/lt5_2_c10 ,open_n4542}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt5_2_cin  (
    .a(1'b0),
    .o({\u2_Display/lt5_2_c0 ,open_n4545}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt5_2_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt5_2_c13 ),
    .o({open_n4546,\u2_Display/n97 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_0  (
    .a(\u2_Display/n1714 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c0 ),
    .o({\u2_Display/lt60_c1 ,open_n4547}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_1  (
    .a(\u2_Display/n1713 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c1 ),
    .o({\u2_Display/lt60_c2 ,open_n4548}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_10  (
    .a(\u2_Display/n1704 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c10 ),
    .o({\u2_Display/lt60_c11 ,open_n4549}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_11  (
    .a(\u2_Display/n1703 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c11 ),
    .o({\u2_Display/lt60_c12 ,open_n4550}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_12  (
    .a(\u2_Display/n1702 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c12 ),
    .o({\u2_Display/lt60_c13 ,open_n4551}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_13  (
    .a(\u2_Display/n1701 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c13 ),
    .o({\u2_Display/lt60_c14 ,open_n4552}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_14  (
    .a(\u2_Display/n1700 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c14 ),
    .o({\u2_Display/lt60_c15 ,open_n4553}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_15  (
    .a(\u2_Display/n1699 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c15 ),
    .o({\u2_Display/lt60_c16 ,open_n4554}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_16  (
    .a(\u2_Display/n1698 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c16 ),
    .o({\u2_Display/lt60_c17 ,open_n4555}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_17  (
    .a(\u2_Display/n1697 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c17 ),
    .o({\u2_Display/lt60_c18 ,open_n4556}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_18  (
    .a(\u2_Display/n1696 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c18 ),
    .o({\u2_Display/lt60_c19 ,open_n4557}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_19  (
    .a(\u2_Display/n1695 ),
    .b(1'b1),
    .c(\u2_Display/lt60_c19 ),
    .o({\u2_Display/lt60_c20 ,open_n4558}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_2  (
    .a(\u2_Display/n1712 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c2 ),
    .o({\u2_Display/lt60_c3 ,open_n4559}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_20  (
    .a(\u2_Display/n1694 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c20 ),
    .o({\u2_Display/lt60_c21 ,open_n4560}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_21  (
    .a(\u2_Display/n1693 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c21 ),
    .o({\u2_Display/lt60_c22 ,open_n4561}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_22  (
    .a(\u2_Display/n1692 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c22 ),
    .o({\u2_Display/lt60_c23 ,open_n4562}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_23  (
    .a(\u2_Display/n1691 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c23 ),
    .o({\u2_Display/lt60_c24 ,open_n4563}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_24  (
    .a(\u2_Display/n1690 ),
    .b(1'b1),
    .c(\u2_Display/lt60_c24 ),
    .o({\u2_Display/lt60_c25 ,open_n4564}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_25  (
    .a(\u2_Display/n1689 ),
    .b(1'b1),
    .c(\u2_Display/lt60_c25 ),
    .o({\u2_Display/lt60_c26 ,open_n4565}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_26  (
    .a(\u2_Display/n1688 ),
    .b(1'b1),
    .c(\u2_Display/lt60_c26 ),
    .o({\u2_Display/lt60_c27 ,open_n4566}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_27  (
    .a(\u2_Display/n1687 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c27 ),
    .o({\u2_Display/lt60_c28 ,open_n4567}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_28  (
    .a(\u2_Display/n1686 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c28 ),
    .o({\u2_Display/lt60_c29 ,open_n4568}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_29  (
    .a(\u2_Display/n1685 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c29 ),
    .o({\u2_Display/lt60_c30 ,open_n4569}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_3  (
    .a(\u2_Display/n1711 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c3 ),
    .o({\u2_Display/lt60_c4 ,open_n4570}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_30  (
    .a(\u2_Display/n1684 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c30 ),
    .o({\u2_Display/lt60_c31 ,open_n4571}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_31  (
    .a(\u2_Display/n1683 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c31 ),
    .o({\u2_Display/lt60_c32 ,open_n4572}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_4  (
    .a(\u2_Display/n1710 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c4 ),
    .o({\u2_Display/lt60_c5 ,open_n4573}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_5  (
    .a(\u2_Display/n1709 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c5 ),
    .o({\u2_Display/lt60_c6 ,open_n4574}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_6  (
    .a(\u2_Display/n1708 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c6 ),
    .o({\u2_Display/lt60_c7 ,open_n4575}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_7  (
    .a(\u2_Display/n1707 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c7 ),
    .o({\u2_Display/lt60_c8 ,open_n4576}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_8  (
    .a(\u2_Display/n1706 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c8 ),
    .o({\u2_Display/lt60_c9 ,open_n4577}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_9  (
    .a(\u2_Display/n1705 ),
    .b(1'b0),
    .c(\u2_Display/lt60_c9 ),
    .o({\u2_Display/lt60_c10 ,open_n4578}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt60_cin  (
    .a(1'b0),
    .o({\u2_Display/lt60_c0 ,open_n4581}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt60_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt60_c32 ),
    .o({open_n4582,\u2_Display/n1715 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_0  (
    .a(\u2_Display/n1749 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c0 ),
    .o({\u2_Display/lt61_c1 ,open_n4583}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_1  (
    .a(\u2_Display/n1748 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c1 ),
    .o({\u2_Display/lt61_c2 ,open_n4584}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_10  (
    .a(\u2_Display/n1739 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c10 ),
    .o({\u2_Display/lt61_c11 ,open_n4585}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_11  (
    .a(\u2_Display/n1738 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c11 ),
    .o({\u2_Display/lt61_c12 ,open_n4586}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_12  (
    .a(\u2_Display/n1737 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c12 ),
    .o({\u2_Display/lt61_c13 ,open_n4587}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_13  (
    .a(\u2_Display/n1736 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c13 ),
    .o({\u2_Display/lt61_c14 ,open_n4588}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_14  (
    .a(\u2_Display/n1735 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c14 ),
    .o({\u2_Display/lt61_c15 ,open_n4589}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_15  (
    .a(\u2_Display/n1734 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c15 ),
    .o({\u2_Display/lt61_c16 ,open_n4590}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_16  (
    .a(\u2_Display/n1733 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c16 ),
    .o({\u2_Display/lt61_c17 ,open_n4591}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_17  (
    .a(\u2_Display/n1732 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c17 ),
    .o({\u2_Display/lt61_c18 ,open_n4592}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_18  (
    .a(\u2_Display/n1731 ),
    .b(1'b1),
    .c(\u2_Display/lt61_c18 ),
    .o({\u2_Display/lt61_c19 ,open_n4593}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_19  (
    .a(\u2_Display/n1730 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c19 ),
    .o({\u2_Display/lt61_c20 ,open_n4594}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_2  (
    .a(\u2_Display/n1747 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c2 ),
    .o({\u2_Display/lt61_c3 ,open_n4595}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_20  (
    .a(\u2_Display/n1729 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c20 ),
    .o({\u2_Display/lt61_c21 ,open_n4596}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_21  (
    .a(\u2_Display/n1728 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c21 ),
    .o({\u2_Display/lt61_c22 ,open_n4597}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_22  (
    .a(\u2_Display/n1727 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c22 ),
    .o({\u2_Display/lt61_c23 ,open_n4598}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_23  (
    .a(\u2_Display/n1726 ),
    .b(1'b1),
    .c(\u2_Display/lt61_c23 ),
    .o({\u2_Display/lt61_c24 ,open_n4599}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_24  (
    .a(\u2_Display/n1725 ),
    .b(1'b1),
    .c(\u2_Display/lt61_c24 ),
    .o({\u2_Display/lt61_c25 ,open_n4600}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_25  (
    .a(\u2_Display/n1724 ),
    .b(1'b1),
    .c(\u2_Display/lt61_c25 ),
    .o({\u2_Display/lt61_c26 ,open_n4601}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_26  (
    .a(\u2_Display/n1723 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c26 ),
    .o({\u2_Display/lt61_c27 ,open_n4602}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_27  (
    .a(\u2_Display/n1722 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c27 ),
    .o({\u2_Display/lt61_c28 ,open_n4603}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_28  (
    .a(\u2_Display/n1721 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c28 ),
    .o({\u2_Display/lt61_c29 ,open_n4604}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_29  (
    .a(\u2_Display/n1720 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c29 ),
    .o({\u2_Display/lt61_c30 ,open_n4605}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_3  (
    .a(\u2_Display/n1746 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c3 ),
    .o({\u2_Display/lt61_c4 ,open_n4606}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_30  (
    .a(\u2_Display/n1719 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c30 ),
    .o({\u2_Display/lt61_c31 ,open_n4607}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_31  (
    .a(\u2_Display/n1718 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c31 ),
    .o({\u2_Display/lt61_c32 ,open_n4608}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_4  (
    .a(\u2_Display/n1745 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c4 ),
    .o({\u2_Display/lt61_c5 ,open_n4609}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_5  (
    .a(\u2_Display/n1744 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c5 ),
    .o({\u2_Display/lt61_c6 ,open_n4610}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_6  (
    .a(\u2_Display/n1743 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c6 ),
    .o({\u2_Display/lt61_c7 ,open_n4611}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_7  (
    .a(\u2_Display/n1742 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c7 ),
    .o({\u2_Display/lt61_c8 ,open_n4612}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_8  (
    .a(\u2_Display/n1741 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c8 ),
    .o({\u2_Display/lt61_c9 ,open_n4613}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_9  (
    .a(\u2_Display/n1740 ),
    .b(1'b0),
    .c(\u2_Display/lt61_c9 ),
    .o({\u2_Display/lt61_c10 ,open_n4614}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt61_cin  (
    .a(1'b0),
    .o({\u2_Display/lt61_c0 ,open_n4617}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt61_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt61_c32 ),
    .o({open_n4618,\u2_Display/n1750 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_0  (
    .a(\u2_Display/n1784 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c0 ),
    .o({\u2_Display/lt62_c1 ,open_n4619}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_1  (
    .a(\u2_Display/n1783 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c1 ),
    .o({\u2_Display/lt62_c2 ,open_n4620}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_10  (
    .a(\u2_Display/n1774 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c10 ),
    .o({\u2_Display/lt62_c11 ,open_n4621}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_11  (
    .a(\u2_Display/n1773 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c11 ),
    .o({\u2_Display/lt62_c12 ,open_n4622}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_12  (
    .a(\u2_Display/n1772 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c12 ),
    .o({\u2_Display/lt62_c13 ,open_n4623}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_13  (
    .a(\u2_Display/n1771 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c13 ),
    .o({\u2_Display/lt62_c14 ,open_n4624}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_14  (
    .a(\u2_Display/n1770 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c14 ),
    .o({\u2_Display/lt62_c15 ,open_n4625}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_15  (
    .a(\u2_Display/n1769 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c15 ),
    .o({\u2_Display/lt62_c16 ,open_n4626}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_16  (
    .a(\u2_Display/n1768 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c16 ),
    .o({\u2_Display/lt62_c17 ,open_n4627}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_17  (
    .a(\u2_Display/n1767 ),
    .b(1'b1),
    .c(\u2_Display/lt62_c17 ),
    .o({\u2_Display/lt62_c18 ,open_n4628}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_18  (
    .a(\u2_Display/n1766 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c18 ),
    .o({\u2_Display/lt62_c19 ,open_n4629}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_19  (
    .a(\u2_Display/n1765 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c19 ),
    .o({\u2_Display/lt62_c20 ,open_n4630}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_2  (
    .a(\u2_Display/n1782 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c2 ),
    .o({\u2_Display/lt62_c3 ,open_n4631}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_20  (
    .a(\u2_Display/n1764 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c20 ),
    .o({\u2_Display/lt62_c21 ,open_n4632}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_21  (
    .a(\u2_Display/n1763 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c21 ),
    .o({\u2_Display/lt62_c22 ,open_n4633}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_22  (
    .a(\u2_Display/n1762 ),
    .b(1'b1),
    .c(\u2_Display/lt62_c22 ),
    .o({\u2_Display/lt62_c23 ,open_n4634}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_23  (
    .a(\u2_Display/n1761 ),
    .b(1'b1),
    .c(\u2_Display/lt62_c23 ),
    .o({\u2_Display/lt62_c24 ,open_n4635}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_24  (
    .a(\u2_Display/n1760 ),
    .b(1'b1),
    .c(\u2_Display/lt62_c24 ),
    .o({\u2_Display/lt62_c25 ,open_n4636}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_25  (
    .a(\u2_Display/n1759 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c25 ),
    .o({\u2_Display/lt62_c26 ,open_n4637}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_26  (
    .a(\u2_Display/n1758 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c26 ),
    .o({\u2_Display/lt62_c27 ,open_n4638}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_27  (
    .a(\u2_Display/n1757 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c27 ),
    .o({\u2_Display/lt62_c28 ,open_n4639}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_28  (
    .a(\u2_Display/n1756 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c28 ),
    .o({\u2_Display/lt62_c29 ,open_n4640}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_29  (
    .a(\u2_Display/n1755 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c29 ),
    .o({\u2_Display/lt62_c30 ,open_n4641}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_3  (
    .a(\u2_Display/n1781 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c3 ),
    .o({\u2_Display/lt62_c4 ,open_n4642}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_30  (
    .a(\u2_Display/n1754 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c30 ),
    .o({\u2_Display/lt62_c31 ,open_n4643}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_31  (
    .a(\u2_Display/n1753 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c31 ),
    .o({\u2_Display/lt62_c32 ,open_n4644}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_4  (
    .a(\u2_Display/n1780 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c4 ),
    .o({\u2_Display/lt62_c5 ,open_n4645}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_5  (
    .a(\u2_Display/n1779 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c5 ),
    .o({\u2_Display/lt62_c6 ,open_n4646}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_6  (
    .a(\u2_Display/n1778 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c6 ),
    .o({\u2_Display/lt62_c7 ,open_n4647}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_7  (
    .a(\u2_Display/n1777 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c7 ),
    .o({\u2_Display/lt62_c8 ,open_n4648}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_8  (
    .a(\u2_Display/n1776 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c8 ),
    .o({\u2_Display/lt62_c9 ,open_n4649}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_9  (
    .a(\u2_Display/n1775 ),
    .b(1'b0),
    .c(\u2_Display/lt62_c9 ),
    .o({\u2_Display/lt62_c10 ,open_n4650}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt62_cin  (
    .a(1'b0),
    .o({\u2_Display/lt62_c0 ,open_n4653}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt62_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt62_c32 ),
    .o({open_n4654,\u2_Display/n1785 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_0  (
    .a(\u2_Display/n1819 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c0 ),
    .o({\u2_Display/lt63_c1 ,open_n4655}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_1  (
    .a(\u2_Display/n1818 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c1 ),
    .o({\u2_Display/lt63_c2 ,open_n4656}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_10  (
    .a(\u2_Display/n1809 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c10 ),
    .o({\u2_Display/lt63_c11 ,open_n4657}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_11  (
    .a(\u2_Display/n1808 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c11 ),
    .o({\u2_Display/lt63_c12 ,open_n4658}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_12  (
    .a(\u2_Display/n1807 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c12 ),
    .o({\u2_Display/lt63_c13 ,open_n4659}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_13  (
    .a(\u2_Display/n1806 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c13 ),
    .o({\u2_Display/lt63_c14 ,open_n4660}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_14  (
    .a(\u2_Display/n1805 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c14 ),
    .o({\u2_Display/lt63_c15 ,open_n4661}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_15  (
    .a(\u2_Display/n1804 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c15 ),
    .o({\u2_Display/lt63_c16 ,open_n4662}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_16  (
    .a(\u2_Display/n1803 ),
    .b(1'b1),
    .c(\u2_Display/lt63_c16 ),
    .o({\u2_Display/lt63_c17 ,open_n4663}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_17  (
    .a(\u2_Display/n1802 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c17 ),
    .o({\u2_Display/lt63_c18 ,open_n4664}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_18  (
    .a(\u2_Display/n1801 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c18 ),
    .o({\u2_Display/lt63_c19 ,open_n4665}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_19  (
    .a(\u2_Display/n1800 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c19 ),
    .o({\u2_Display/lt63_c20 ,open_n4666}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_2  (
    .a(\u2_Display/n1817 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c2 ),
    .o({\u2_Display/lt63_c3 ,open_n4667}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_20  (
    .a(\u2_Display/n1799 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c20 ),
    .o({\u2_Display/lt63_c21 ,open_n4668}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_21  (
    .a(\u2_Display/n1798 ),
    .b(1'b1),
    .c(\u2_Display/lt63_c21 ),
    .o({\u2_Display/lt63_c22 ,open_n4669}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_22  (
    .a(\u2_Display/n1797 ),
    .b(1'b1),
    .c(\u2_Display/lt63_c22 ),
    .o({\u2_Display/lt63_c23 ,open_n4670}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_23  (
    .a(\u2_Display/n1796 ),
    .b(1'b1),
    .c(\u2_Display/lt63_c23 ),
    .o({\u2_Display/lt63_c24 ,open_n4671}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_24  (
    .a(\u2_Display/n1795 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c24 ),
    .o({\u2_Display/lt63_c25 ,open_n4672}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_25  (
    .a(\u2_Display/n1794 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c25 ),
    .o({\u2_Display/lt63_c26 ,open_n4673}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_26  (
    .a(\u2_Display/n1793 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c26 ),
    .o({\u2_Display/lt63_c27 ,open_n4674}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_27  (
    .a(\u2_Display/n1792 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c27 ),
    .o({\u2_Display/lt63_c28 ,open_n4675}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_28  (
    .a(\u2_Display/n1791 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c28 ),
    .o({\u2_Display/lt63_c29 ,open_n4676}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_29  (
    .a(\u2_Display/n1790 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c29 ),
    .o({\u2_Display/lt63_c30 ,open_n4677}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_3  (
    .a(\u2_Display/n1816 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c3 ),
    .o({\u2_Display/lt63_c4 ,open_n4678}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_30  (
    .a(\u2_Display/n1789 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c30 ),
    .o({\u2_Display/lt63_c31 ,open_n4679}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_31  (
    .a(\u2_Display/n1788 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c31 ),
    .o({\u2_Display/lt63_c32 ,open_n4680}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_4  (
    .a(\u2_Display/n1815 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c4 ),
    .o({\u2_Display/lt63_c5 ,open_n4681}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_5  (
    .a(\u2_Display/n1814 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c5 ),
    .o({\u2_Display/lt63_c6 ,open_n4682}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_6  (
    .a(\u2_Display/n1813 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c6 ),
    .o({\u2_Display/lt63_c7 ,open_n4683}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_7  (
    .a(\u2_Display/n1812 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c7 ),
    .o({\u2_Display/lt63_c8 ,open_n4684}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_8  (
    .a(\u2_Display/n1811 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c8 ),
    .o({\u2_Display/lt63_c9 ,open_n4685}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_9  (
    .a(\u2_Display/n1810 ),
    .b(1'b0),
    .c(\u2_Display/lt63_c9 ),
    .o({\u2_Display/lt63_c10 ,open_n4686}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt63_cin  (
    .a(1'b0),
    .o({\u2_Display/lt63_c0 ,open_n4689}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt63_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt63_c32 ),
    .o({open_n4690,\u2_Display/n1820 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_0  (
    .a(\u2_Display/n1854 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c0 ),
    .o({\u2_Display/lt64_c1 ,open_n4691}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_1  (
    .a(\u2_Display/n1853 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c1 ),
    .o({\u2_Display/lt64_c2 ,open_n4692}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_10  (
    .a(\u2_Display/n1844 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c10 ),
    .o({\u2_Display/lt64_c11 ,open_n4693}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_11  (
    .a(\u2_Display/n1843 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c11 ),
    .o({\u2_Display/lt64_c12 ,open_n4694}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_12  (
    .a(\u2_Display/n1842 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c12 ),
    .o({\u2_Display/lt64_c13 ,open_n4695}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_13  (
    .a(\u2_Display/n1841 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c13 ),
    .o({\u2_Display/lt64_c14 ,open_n4696}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_14  (
    .a(\u2_Display/n1840 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c14 ),
    .o({\u2_Display/lt64_c15 ,open_n4697}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_15  (
    .a(\u2_Display/n1839 ),
    .b(1'b1),
    .c(\u2_Display/lt64_c15 ),
    .o({\u2_Display/lt64_c16 ,open_n4698}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_16  (
    .a(\u2_Display/n1838 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c16 ),
    .o({\u2_Display/lt64_c17 ,open_n4699}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_17  (
    .a(\u2_Display/n1837 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c17 ),
    .o({\u2_Display/lt64_c18 ,open_n4700}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_18  (
    .a(\u2_Display/n1836 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c18 ),
    .o({\u2_Display/lt64_c19 ,open_n4701}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_19  (
    .a(\u2_Display/n1835 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c19 ),
    .o({\u2_Display/lt64_c20 ,open_n4702}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_2  (
    .a(\u2_Display/n1852 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c2 ),
    .o({\u2_Display/lt64_c3 ,open_n4703}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_20  (
    .a(\u2_Display/n1834 ),
    .b(1'b1),
    .c(\u2_Display/lt64_c20 ),
    .o({\u2_Display/lt64_c21 ,open_n4704}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_21  (
    .a(\u2_Display/n1833 ),
    .b(1'b1),
    .c(\u2_Display/lt64_c21 ),
    .o({\u2_Display/lt64_c22 ,open_n4705}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_22  (
    .a(\u2_Display/n1832 ),
    .b(1'b1),
    .c(\u2_Display/lt64_c22 ),
    .o({\u2_Display/lt64_c23 ,open_n4706}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_23  (
    .a(\u2_Display/n1831 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c23 ),
    .o({\u2_Display/lt64_c24 ,open_n4707}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_24  (
    .a(\u2_Display/n1830 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c24 ),
    .o({\u2_Display/lt64_c25 ,open_n4708}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_25  (
    .a(\u2_Display/n1829 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c25 ),
    .o({\u2_Display/lt64_c26 ,open_n4709}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_26  (
    .a(\u2_Display/n1828 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c26 ),
    .o({\u2_Display/lt64_c27 ,open_n4710}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_27  (
    .a(\u2_Display/n1827 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c27 ),
    .o({\u2_Display/lt64_c28 ,open_n4711}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_28  (
    .a(\u2_Display/n1826 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c28 ),
    .o({\u2_Display/lt64_c29 ,open_n4712}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_29  (
    .a(\u2_Display/n1825 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c29 ),
    .o({\u2_Display/lt64_c30 ,open_n4713}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_3  (
    .a(\u2_Display/n1851 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c3 ),
    .o({\u2_Display/lt64_c4 ,open_n4714}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_30  (
    .a(\u2_Display/n1824 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c30 ),
    .o({\u2_Display/lt64_c31 ,open_n4715}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_31  (
    .a(\u2_Display/n1823 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c31 ),
    .o({\u2_Display/lt64_c32 ,open_n4716}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_4  (
    .a(\u2_Display/n1850 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c4 ),
    .o({\u2_Display/lt64_c5 ,open_n4717}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_5  (
    .a(\u2_Display/n1849 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c5 ),
    .o({\u2_Display/lt64_c6 ,open_n4718}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_6  (
    .a(\u2_Display/n1848 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c6 ),
    .o({\u2_Display/lt64_c7 ,open_n4719}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_7  (
    .a(\u2_Display/n1847 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c7 ),
    .o({\u2_Display/lt64_c8 ,open_n4720}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_8  (
    .a(\u2_Display/n1846 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c8 ),
    .o({\u2_Display/lt64_c9 ,open_n4721}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_9  (
    .a(\u2_Display/n1845 ),
    .b(1'b0),
    .c(\u2_Display/lt64_c9 ),
    .o({\u2_Display/lt64_c10 ,open_n4722}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt64_cin  (
    .a(1'b0),
    .o({\u2_Display/lt64_c0 ,open_n4725}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt64_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt64_c32 ),
    .o({open_n4726,\u2_Display/n1855 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_0  (
    .a(\u2_Display/n1889 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c0 ),
    .o({\u2_Display/lt65_c1 ,open_n4727}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_1  (
    .a(\u2_Display/n1888 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c1 ),
    .o({\u2_Display/lt65_c2 ,open_n4728}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_10  (
    .a(\u2_Display/n1879 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c10 ),
    .o({\u2_Display/lt65_c11 ,open_n4729}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_11  (
    .a(\u2_Display/n1878 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c11 ),
    .o({\u2_Display/lt65_c12 ,open_n4730}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_12  (
    .a(\u2_Display/n1877 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c12 ),
    .o({\u2_Display/lt65_c13 ,open_n4731}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_13  (
    .a(\u2_Display/n1876 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c13 ),
    .o({\u2_Display/lt65_c14 ,open_n4732}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_14  (
    .a(\u2_Display/n1875 ),
    .b(1'b1),
    .c(\u2_Display/lt65_c14 ),
    .o({\u2_Display/lt65_c15 ,open_n4733}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_15  (
    .a(\u2_Display/n1874 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c15 ),
    .o({\u2_Display/lt65_c16 ,open_n4734}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_16  (
    .a(\u2_Display/n1873 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c16 ),
    .o({\u2_Display/lt65_c17 ,open_n4735}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_17  (
    .a(\u2_Display/n1872 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c17 ),
    .o({\u2_Display/lt65_c18 ,open_n4736}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_18  (
    .a(\u2_Display/n1871 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c18 ),
    .o({\u2_Display/lt65_c19 ,open_n4737}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_19  (
    .a(\u2_Display/n1870 ),
    .b(1'b1),
    .c(\u2_Display/lt65_c19 ),
    .o({\u2_Display/lt65_c20 ,open_n4738}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_2  (
    .a(\u2_Display/n1887 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c2 ),
    .o({\u2_Display/lt65_c3 ,open_n4739}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_20  (
    .a(\u2_Display/n1869 ),
    .b(1'b1),
    .c(\u2_Display/lt65_c20 ),
    .o({\u2_Display/lt65_c21 ,open_n4740}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_21  (
    .a(\u2_Display/n1868 ),
    .b(1'b1),
    .c(\u2_Display/lt65_c21 ),
    .o({\u2_Display/lt65_c22 ,open_n4741}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_22  (
    .a(\u2_Display/n1867 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c22 ),
    .o({\u2_Display/lt65_c23 ,open_n4742}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_23  (
    .a(\u2_Display/n1866 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c23 ),
    .o({\u2_Display/lt65_c24 ,open_n4743}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_24  (
    .a(\u2_Display/n1865 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c24 ),
    .o({\u2_Display/lt65_c25 ,open_n4744}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_25  (
    .a(\u2_Display/n1864 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c25 ),
    .o({\u2_Display/lt65_c26 ,open_n4745}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_26  (
    .a(\u2_Display/n1863 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c26 ),
    .o({\u2_Display/lt65_c27 ,open_n4746}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_27  (
    .a(\u2_Display/n1862 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c27 ),
    .o({\u2_Display/lt65_c28 ,open_n4747}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_28  (
    .a(\u2_Display/n1861 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c28 ),
    .o({\u2_Display/lt65_c29 ,open_n4748}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_29  (
    .a(\u2_Display/n1860 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c29 ),
    .o({\u2_Display/lt65_c30 ,open_n4749}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_3  (
    .a(\u2_Display/n1886 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c3 ),
    .o({\u2_Display/lt65_c4 ,open_n4750}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_30  (
    .a(\u2_Display/n1859 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c30 ),
    .o({\u2_Display/lt65_c31 ,open_n4751}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_31  (
    .a(\u2_Display/n1858 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c31 ),
    .o({\u2_Display/lt65_c32 ,open_n4752}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_4  (
    .a(\u2_Display/n1885 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c4 ),
    .o({\u2_Display/lt65_c5 ,open_n4753}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_5  (
    .a(\u2_Display/n1884 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c5 ),
    .o({\u2_Display/lt65_c6 ,open_n4754}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_6  (
    .a(\u2_Display/n1883 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c6 ),
    .o({\u2_Display/lt65_c7 ,open_n4755}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_7  (
    .a(\u2_Display/n1882 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c7 ),
    .o({\u2_Display/lt65_c8 ,open_n4756}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_8  (
    .a(\u2_Display/n1881 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c8 ),
    .o({\u2_Display/lt65_c9 ,open_n4757}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_9  (
    .a(\u2_Display/n1880 ),
    .b(1'b0),
    .c(\u2_Display/lt65_c9 ),
    .o({\u2_Display/lt65_c10 ,open_n4758}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt65_cin  (
    .a(1'b0),
    .o({\u2_Display/lt65_c0 ,open_n4761}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt65_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt65_c32 ),
    .o({open_n4762,\u2_Display/n1890 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_0  (
    .a(\u2_Display/n1924 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c0 ),
    .o({\u2_Display/lt66_c1 ,open_n4763}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_1  (
    .a(\u2_Display/n1923 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c1 ),
    .o({\u2_Display/lt66_c2 ,open_n4764}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_10  (
    .a(\u2_Display/n1914 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c10 ),
    .o({\u2_Display/lt66_c11 ,open_n4765}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_11  (
    .a(\u2_Display/n1913 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c11 ),
    .o({\u2_Display/lt66_c12 ,open_n4766}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_12  (
    .a(\u2_Display/n1912 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c12 ),
    .o({\u2_Display/lt66_c13 ,open_n4767}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_13  (
    .a(\u2_Display/n1911 ),
    .b(1'b1),
    .c(\u2_Display/lt66_c13 ),
    .o({\u2_Display/lt66_c14 ,open_n4768}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_14  (
    .a(\u2_Display/n1910 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c14 ),
    .o({\u2_Display/lt66_c15 ,open_n4769}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_15  (
    .a(\u2_Display/n1909 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c15 ),
    .o({\u2_Display/lt66_c16 ,open_n4770}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_16  (
    .a(\u2_Display/n1908 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c16 ),
    .o({\u2_Display/lt66_c17 ,open_n4771}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_17  (
    .a(\u2_Display/n1907 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c17 ),
    .o({\u2_Display/lt66_c18 ,open_n4772}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_18  (
    .a(\u2_Display/n1906 ),
    .b(1'b1),
    .c(\u2_Display/lt66_c18 ),
    .o({\u2_Display/lt66_c19 ,open_n4773}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_19  (
    .a(\u2_Display/n1905 ),
    .b(1'b1),
    .c(\u2_Display/lt66_c19 ),
    .o({\u2_Display/lt66_c20 ,open_n4774}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_2  (
    .a(\u2_Display/n1922 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c2 ),
    .o({\u2_Display/lt66_c3 ,open_n4775}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_20  (
    .a(\u2_Display/n1904 ),
    .b(1'b1),
    .c(\u2_Display/lt66_c20 ),
    .o({\u2_Display/lt66_c21 ,open_n4776}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_21  (
    .a(\u2_Display/n1903 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c21 ),
    .o({\u2_Display/lt66_c22 ,open_n4777}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_22  (
    .a(\u2_Display/n1902 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c22 ),
    .o({\u2_Display/lt66_c23 ,open_n4778}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_23  (
    .a(\u2_Display/n1901 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c23 ),
    .o({\u2_Display/lt66_c24 ,open_n4779}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_24  (
    .a(\u2_Display/n1900 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c24 ),
    .o({\u2_Display/lt66_c25 ,open_n4780}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_25  (
    .a(\u2_Display/n1899 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c25 ),
    .o({\u2_Display/lt66_c26 ,open_n4781}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_26  (
    .a(\u2_Display/n1898 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c26 ),
    .o({\u2_Display/lt66_c27 ,open_n4782}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_27  (
    .a(\u2_Display/n1897 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c27 ),
    .o({\u2_Display/lt66_c28 ,open_n4783}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_28  (
    .a(\u2_Display/n1896 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c28 ),
    .o({\u2_Display/lt66_c29 ,open_n4784}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_29  (
    .a(\u2_Display/n1895 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c29 ),
    .o({\u2_Display/lt66_c30 ,open_n4785}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_3  (
    .a(\u2_Display/n1921 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c3 ),
    .o({\u2_Display/lt66_c4 ,open_n4786}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_30  (
    .a(\u2_Display/n1894 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c30 ),
    .o({\u2_Display/lt66_c31 ,open_n4787}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_31  (
    .a(\u2_Display/n1893 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c31 ),
    .o({\u2_Display/lt66_c32 ,open_n4788}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_4  (
    .a(\u2_Display/n1920 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c4 ),
    .o({\u2_Display/lt66_c5 ,open_n4789}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_5  (
    .a(\u2_Display/n1919 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c5 ),
    .o({\u2_Display/lt66_c6 ,open_n4790}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_6  (
    .a(\u2_Display/n1918 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c6 ),
    .o({\u2_Display/lt66_c7 ,open_n4791}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_7  (
    .a(\u2_Display/n1917 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c7 ),
    .o({\u2_Display/lt66_c8 ,open_n4792}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_8  (
    .a(\u2_Display/n1916 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c8 ),
    .o({\u2_Display/lt66_c9 ,open_n4793}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_9  (
    .a(\u2_Display/n1915 ),
    .b(1'b0),
    .c(\u2_Display/lt66_c9 ),
    .o({\u2_Display/lt66_c10 ,open_n4794}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt66_cin  (
    .a(1'b0),
    .o({\u2_Display/lt66_c0 ,open_n4797}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt66_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt66_c32 ),
    .o({open_n4798,\u2_Display/n1925 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_0  (
    .a(\u2_Display/n1959 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c0 ),
    .o({\u2_Display/lt67_c1 ,open_n4799}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_1  (
    .a(\u2_Display/n1958 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c1 ),
    .o({\u2_Display/lt67_c2 ,open_n4800}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_10  (
    .a(\u2_Display/n1949 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c10 ),
    .o({\u2_Display/lt67_c11 ,open_n4801}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_11  (
    .a(\u2_Display/n1948 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c11 ),
    .o({\u2_Display/lt67_c12 ,open_n4802}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_12  (
    .a(\u2_Display/n1947 ),
    .b(1'b1),
    .c(\u2_Display/lt67_c12 ),
    .o({\u2_Display/lt67_c13 ,open_n4803}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_13  (
    .a(\u2_Display/n1946 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c13 ),
    .o({\u2_Display/lt67_c14 ,open_n4804}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_14  (
    .a(\u2_Display/n1945 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c14 ),
    .o({\u2_Display/lt67_c15 ,open_n4805}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_15  (
    .a(\u2_Display/n1944 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c15 ),
    .o({\u2_Display/lt67_c16 ,open_n4806}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_16  (
    .a(\u2_Display/n1943 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c16 ),
    .o({\u2_Display/lt67_c17 ,open_n4807}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_17  (
    .a(\u2_Display/n1942 ),
    .b(1'b1),
    .c(\u2_Display/lt67_c17 ),
    .o({\u2_Display/lt67_c18 ,open_n4808}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_18  (
    .a(\u2_Display/n1941 ),
    .b(1'b1),
    .c(\u2_Display/lt67_c18 ),
    .o({\u2_Display/lt67_c19 ,open_n4809}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_19  (
    .a(\u2_Display/n1940 ),
    .b(1'b1),
    .c(\u2_Display/lt67_c19 ),
    .o({\u2_Display/lt67_c20 ,open_n4810}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_2  (
    .a(\u2_Display/n1957 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c2 ),
    .o({\u2_Display/lt67_c3 ,open_n4811}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_20  (
    .a(\u2_Display/n1939 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c20 ),
    .o({\u2_Display/lt67_c21 ,open_n4812}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_21  (
    .a(\u2_Display/n1938 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c21 ),
    .o({\u2_Display/lt67_c22 ,open_n4813}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_22  (
    .a(\u2_Display/n1937 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c22 ),
    .o({\u2_Display/lt67_c23 ,open_n4814}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_23  (
    .a(\u2_Display/n1936 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c23 ),
    .o({\u2_Display/lt67_c24 ,open_n4815}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_24  (
    .a(\u2_Display/n1935 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c24 ),
    .o({\u2_Display/lt67_c25 ,open_n4816}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_25  (
    .a(\u2_Display/n1934 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c25 ),
    .o({\u2_Display/lt67_c26 ,open_n4817}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_26  (
    .a(\u2_Display/n1933 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c26 ),
    .o({\u2_Display/lt67_c27 ,open_n4818}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_27  (
    .a(\u2_Display/n1932 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c27 ),
    .o({\u2_Display/lt67_c28 ,open_n4819}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_28  (
    .a(\u2_Display/n1931 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c28 ),
    .o({\u2_Display/lt67_c29 ,open_n4820}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_29  (
    .a(\u2_Display/n1930 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c29 ),
    .o({\u2_Display/lt67_c30 ,open_n4821}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_3  (
    .a(\u2_Display/n1956 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c3 ),
    .o({\u2_Display/lt67_c4 ,open_n4822}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_30  (
    .a(\u2_Display/n1929 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c30 ),
    .o({\u2_Display/lt67_c31 ,open_n4823}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_31  (
    .a(\u2_Display/n1928 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c31 ),
    .o({\u2_Display/lt67_c32 ,open_n4824}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_4  (
    .a(\u2_Display/n1955 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c4 ),
    .o({\u2_Display/lt67_c5 ,open_n4825}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_5  (
    .a(\u2_Display/n1954 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c5 ),
    .o({\u2_Display/lt67_c6 ,open_n4826}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_6  (
    .a(\u2_Display/n1953 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c6 ),
    .o({\u2_Display/lt67_c7 ,open_n4827}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_7  (
    .a(\u2_Display/n1952 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c7 ),
    .o({\u2_Display/lt67_c8 ,open_n4828}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_8  (
    .a(\u2_Display/n1951 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c8 ),
    .o({\u2_Display/lt67_c9 ,open_n4829}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_9  (
    .a(\u2_Display/n1950 ),
    .b(1'b0),
    .c(\u2_Display/lt67_c9 ),
    .o({\u2_Display/lt67_c10 ,open_n4830}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt67_cin  (
    .a(1'b0),
    .o({\u2_Display/lt67_c0 ,open_n4833}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt67_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt67_c32 ),
    .o({open_n4834,\u2_Display/n1960 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_0  (
    .a(\u2_Display/n1994 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c0 ),
    .o({\u2_Display/lt68_c1 ,open_n4835}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_1  (
    .a(\u2_Display/n1993 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c1 ),
    .o({\u2_Display/lt68_c2 ,open_n4836}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_10  (
    .a(\u2_Display/n1984 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c10 ),
    .o({\u2_Display/lt68_c11 ,open_n4837}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_11  (
    .a(\u2_Display/n1983 ),
    .b(1'b1),
    .c(\u2_Display/lt68_c11 ),
    .o({\u2_Display/lt68_c12 ,open_n4838}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_12  (
    .a(\u2_Display/n1982 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c12 ),
    .o({\u2_Display/lt68_c13 ,open_n4839}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_13  (
    .a(\u2_Display/n1981 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c13 ),
    .o({\u2_Display/lt68_c14 ,open_n4840}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_14  (
    .a(\u2_Display/n1980 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c14 ),
    .o({\u2_Display/lt68_c15 ,open_n4841}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_15  (
    .a(\u2_Display/n1979 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c15 ),
    .o({\u2_Display/lt68_c16 ,open_n4842}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_16  (
    .a(\u2_Display/n1978 ),
    .b(1'b1),
    .c(\u2_Display/lt68_c16 ),
    .o({\u2_Display/lt68_c17 ,open_n4843}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_17  (
    .a(\u2_Display/n1977 ),
    .b(1'b1),
    .c(\u2_Display/lt68_c17 ),
    .o({\u2_Display/lt68_c18 ,open_n4844}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_18  (
    .a(\u2_Display/n1976 ),
    .b(1'b1),
    .c(\u2_Display/lt68_c18 ),
    .o({\u2_Display/lt68_c19 ,open_n4845}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_19  (
    .a(\u2_Display/n1975 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c19 ),
    .o({\u2_Display/lt68_c20 ,open_n4846}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_2  (
    .a(\u2_Display/n1992 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c2 ),
    .o({\u2_Display/lt68_c3 ,open_n4847}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_20  (
    .a(\u2_Display/n1974 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c20 ),
    .o({\u2_Display/lt68_c21 ,open_n4848}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_21  (
    .a(\u2_Display/n1973 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c21 ),
    .o({\u2_Display/lt68_c22 ,open_n4849}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_22  (
    .a(\u2_Display/n1972 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c22 ),
    .o({\u2_Display/lt68_c23 ,open_n4850}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_23  (
    .a(\u2_Display/n1971 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c23 ),
    .o({\u2_Display/lt68_c24 ,open_n4851}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_24  (
    .a(\u2_Display/n1970 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c24 ),
    .o({\u2_Display/lt68_c25 ,open_n4852}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_25  (
    .a(\u2_Display/n1969 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c25 ),
    .o({\u2_Display/lt68_c26 ,open_n4853}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_26  (
    .a(\u2_Display/n1968 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c26 ),
    .o({\u2_Display/lt68_c27 ,open_n4854}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_27  (
    .a(\u2_Display/n1967 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c27 ),
    .o({\u2_Display/lt68_c28 ,open_n4855}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_28  (
    .a(\u2_Display/n1966 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c28 ),
    .o({\u2_Display/lt68_c29 ,open_n4856}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_29  (
    .a(\u2_Display/n1965 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c29 ),
    .o({\u2_Display/lt68_c30 ,open_n4857}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_3  (
    .a(\u2_Display/n1991 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c3 ),
    .o({\u2_Display/lt68_c4 ,open_n4858}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_30  (
    .a(\u2_Display/n1964 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c30 ),
    .o({\u2_Display/lt68_c31 ,open_n4859}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_31  (
    .a(\u2_Display/n1963 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c31 ),
    .o({\u2_Display/lt68_c32 ,open_n4860}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_4  (
    .a(\u2_Display/n1990 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c4 ),
    .o({\u2_Display/lt68_c5 ,open_n4861}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_5  (
    .a(\u2_Display/n1989 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c5 ),
    .o({\u2_Display/lt68_c6 ,open_n4862}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_6  (
    .a(\u2_Display/n1988 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c6 ),
    .o({\u2_Display/lt68_c7 ,open_n4863}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_7  (
    .a(\u2_Display/n1987 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c7 ),
    .o({\u2_Display/lt68_c8 ,open_n4864}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_8  (
    .a(\u2_Display/n1986 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c8 ),
    .o({\u2_Display/lt68_c9 ,open_n4865}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_9  (
    .a(\u2_Display/n1985 ),
    .b(1'b0),
    .c(\u2_Display/lt68_c9 ),
    .o({\u2_Display/lt68_c10 ,open_n4866}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt68_cin  (
    .a(1'b0),
    .o({\u2_Display/lt68_c0 ,open_n4869}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt68_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt68_c32 ),
    .o({open_n4870,\u2_Display/n1995 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_0  (
    .a(\u2_Display/n2029 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c0 ),
    .o({\u2_Display/lt69_c1 ,open_n4871}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_1  (
    .a(\u2_Display/n2028 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c1 ),
    .o({\u2_Display/lt69_c2 ,open_n4872}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_10  (
    .a(\u2_Display/n2019 ),
    .b(1'b1),
    .c(\u2_Display/lt69_c10 ),
    .o({\u2_Display/lt69_c11 ,open_n4873}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_11  (
    .a(\u2_Display/n2018 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c11 ),
    .o({\u2_Display/lt69_c12 ,open_n4874}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_12  (
    .a(\u2_Display/n2017 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c12 ),
    .o({\u2_Display/lt69_c13 ,open_n4875}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_13  (
    .a(\u2_Display/n2016 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c13 ),
    .o({\u2_Display/lt69_c14 ,open_n4876}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_14  (
    .a(\u2_Display/n2015 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c14 ),
    .o({\u2_Display/lt69_c15 ,open_n4877}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_15  (
    .a(\u2_Display/n2014 ),
    .b(1'b1),
    .c(\u2_Display/lt69_c15 ),
    .o({\u2_Display/lt69_c16 ,open_n4878}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_16  (
    .a(\u2_Display/n2013 ),
    .b(1'b1),
    .c(\u2_Display/lt69_c16 ),
    .o({\u2_Display/lt69_c17 ,open_n4879}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_17  (
    .a(\u2_Display/n2012 ),
    .b(1'b1),
    .c(\u2_Display/lt69_c17 ),
    .o({\u2_Display/lt69_c18 ,open_n4880}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_18  (
    .a(\u2_Display/n2011 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c18 ),
    .o({\u2_Display/lt69_c19 ,open_n4881}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_19  (
    .a(\u2_Display/n2010 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c19 ),
    .o({\u2_Display/lt69_c20 ,open_n4882}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_2  (
    .a(\u2_Display/n2027 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c2 ),
    .o({\u2_Display/lt69_c3 ,open_n4883}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_20  (
    .a(\u2_Display/n2009 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c20 ),
    .o({\u2_Display/lt69_c21 ,open_n4884}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_21  (
    .a(\u2_Display/n2008 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c21 ),
    .o({\u2_Display/lt69_c22 ,open_n4885}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_22  (
    .a(\u2_Display/n2007 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c22 ),
    .o({\u2_Display/lt69_c23 ,open_n4886}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_23  (
    .a(\u2_Display/n2006 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c23 ),
    .o({\u2_Display/lt69_c24 ,open_n4887}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_24  (
    .a(\u2_Display/n2005 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c24 ),
    .o({\u2_Display/lt69_c25 ,open_n4888}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_25  (
    .a(\u2_Display/n2004 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c25 ),
    .o({\u2_Display/lt69_c26 ,open_n4889}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_26  (
    .a(\u2_Display/n2003 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c26 ),
    .o({\u2_Display/lt69_c27 ,open_n4890}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_27  (
    .a(\u2_Display/n2002 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c27 ),
    .o({\u2_Display/lt69_c28 ,open_n4891}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_28  (
    .a(\u2_Display/n2001 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c28 ),
    .o({\u2_Display/lt69_c29 ,open_n4892}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_29  (
    .a(\u2_Display/n2000 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c29 ),
    .o({\u2_Display/lt69_c30 ,open_n4893}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_3  (
    .a(\u2_Display/n2026 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c3 ),
    .o({\u2_Display/lt69_c4 ,open_n4894}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_30  (
    .a(\u2_Display/n1999 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c30 ),
    .o({\u2_Display/lt69_c31 ,open_n4895}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_31  (
    .a(\u2_Display/n1998 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c31 ),
    .o({\u2_Display/lt69_c32 ,open_n4896}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_4  (
    .a(\u2_Display/n2025 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c4 ),
    .o({\u2_Display/lt69_c5 ,open_n4897}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_5  (
    .a(\u2_Display/n2024 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c5 ),
    .o({\u2_Display/lt69_c6 ,open_n4898}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_6  (
    .a(\u2_Display/n2023 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c6 ),
    .o({\u2_Display/lt69_c7 ,open_n4899}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_7  (
    .a(\u2_Display/n2022 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c7 ),
    .o({\u2_Display/lt69_c8 ,open_n4900}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_8  (
    .a(\u2_Display/n2021 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c8 ),
    .o({\u2_Display/lt69_c9 ,open_n4901}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_9  (
    .a(\u2_Display/n2020 ),
    .b(1'b0),
    .c(\u2_Display/lt69_c9 ),
    .o({\u2_Display/lt69_c10 ,open_n4902}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt69_cin  (
    .a(1'b0),
    .o({\u2_Display/lt69_c0 ,open_n4905}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt69_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt69_c32 ),
    .o({open_n4906,\u2_Display/n2030 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt6_2_0  (
    .a(lcd_ypos[0]),
    .b(\u2_Display/j [0]),
    .c(\u2_Display/lt6_2_c0 ),
    .o({\u2_Display/lt6_2_c1 ,open_n4907}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt6_2_1  (
    .a(lcd_ypos[1]),
    .b(\u2_Display/j [1]),
    .c(\u2_Display/lt6_2_c1 ),
    .o({\u2_Display/lt6_2_c2 ,open_n4908}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt6_2_10  (
    .a(lcd_ypos[10]),
    .b(\u2_Display/j [9]),
    .c(\u2_Display/lt6_2_c10 ),
    .o({\u2_Display/lt6_2_c11 ,open_n4909}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt6_2_11  (
    .a(lcd_ypos[11]),
    .b(1'b0),
    .c(\u2_Display/lt6_2_c11 ),
    .o({\u2_Display/lt6_2_c12 ,open_n4910}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt6_2_2  (
    .a(lcd_ypos[2]),
    .b(\u2_Display/j [2]),
    .c(\u2_Display/lt6_2_c2 ),
    .o({\u2_Display/lt6_2_c3 ,open_n4911}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt6_2_3  (
    .a(lcd_ypos[3]),
    .b(\u2_Display/j [3]),
    .c(\u2_Display/lt6_2_c3 ),
    .o({\u2_Display/lt6_2_c4 ,open_n4912}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt6_2_4  (
    .a(lcd_ypos[4]),
    .b(\u2_Display/j [4]),
    .c(\u2_Display/lt6_2_c4 ),
    .o({\u2_Display/lt6_2_c5 ,open_n4913}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt6_2_5  (
    .a(lcd_ypos[5]),
    .b(\u2_Display/j [5]),
    .c(\u2_Display/lt6_2_c5 ),
    .o({\u2_Display/lt6_2_c6 ,open_n4914}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt6_2_6  (
    .a(lcd_ypos[6]),
    .b(\u2_Display/j [6]),
    .c(\u2_Display/lt6_2_c6 ),
    .o({\u2_Display/lt6_2_c7 ,open_n4915}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt6_2_7  (
    .a(lcd_ypos[7]),
    .b(\u2_Display/j [7]),
    .c(\u2_Display/lt6_2_c7 ),
    .o({\u2_Display/lt6_2_c8 ,open_n4916}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt6_2_8  (
    .a(lcd_ypos[8]),
    .b(\u2_Display/j [8]),
    .c(\u2_Display/lt6_2_c8 ),
    .o({\u2_Display/lt6_2_c9 ,open_n4917}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt6_2_9  (
    .a(lcd_ypos[9]),
    .b(\u2_Display/n99 [0]),
    .c(\u2_Display/lt6_2_c9 ),
    .o({\u2_Display/lt6_2_c10 ,open_n4918}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt6_2_cin  (
    .a(1'b0),
    .o({\u2_Display/lt6_2_c0 ,open_n4921}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt6_2_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt6_2_c12 ),
    .o({open_n4922,\u2_Display/n100 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_0  (
    .a(\u2_Display/n2064 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c0 ),
    .o({\u2_Display/lt70_c1 ,open_n4923}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_1  (
    .a(\u2_Display/n2063 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c1 ),
    .o({\u2_Display/lt70_c2 ,open_n4924}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_10  (
    .a(\u2_Display/n2054 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c10 ),
    .o({\u2_Display/lt70_c11 ,open_n4925}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_11  (
    .a(\u2_Display/n2053 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c11 ),
    .o({\u2_Display/lt70_c12 ,open_n4926}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_12  (
    .a(\u2_Display/n2052 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c12 ),
    .o({\u2_Display/lt70_c13 ,open_n4927}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_13  (
    .a(\u2_Display/n2051 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c13 ),
    .o({\u2_Display/lt70_c14 ,open_n4928}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_14  (
    .a(\u2_Display/n2050 ),
    .b(1'b1),
    .c(\u2_Display/lt70_c14 ),
    .o({\u2_Display/lt70_c15 ,open_n4929}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_15  (
    .a(\u2_Display/n2049 ),
    .b(1'b1),
    .c(\u2_Display/lt70_c15 ),
    .o({\u2_Display/lt70_c16 ,open_n4930}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_16  (
    .a(\u2_Display/n2048 ),
    .b(1'b1),
    .c(\u2_Display/lt70_c16 ),
    .o({\u2_Display/lt70_c17 ,open_n4931}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_17  (
    .a(\u2_Display/n2047 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c17 ),
    .o({\u2_Display/lt70_c18 ,open_n4932}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_18  (
    .a(\u2_Display/n2046 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c18 ),
    .o({\u2_Display/lt70_c19 ,open_n4933}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_19  (
    .a(\u2_Display/n2045 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c19 ),
    .o({\u2_Display/lt70_c20 ,open_n4934}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_2  (
    .a(\u2_Display/n2062 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c2 ),
    .o({\u2_Display/lt70_c3 ,open_n4935}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_20  (
    .a(\u2_Display/n2044 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c20 ),
    .o({\u2_Display/lt70_c21 ,open_n4936}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_21  (
    .a(\u2_Display/n2043 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c21 ),
    .o({\u2_Display/lt70_c22 ,open_n4937}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_22  (
    .a(\u2_Display/n2042 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c22 ),
    .o({\u2_Display/lt70_c23 ,open_n4938}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_23  (
    .a(\u2_Display/n2041 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c23 ),
    .o({\u2_Display/lt70_c24 ,open_n4939}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_24  (
    .a(\u2_Display/n2040 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c24 ),
    .o({\u2_Display/lt70_c25 ,open_n4940}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_25  (
    .a(\u2_Display/n2039 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c25 ),
    .o({\u2_Display/lt70_c26 ,open_n4941}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_26  (
    .a(\u2_Display/n2038 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c26 ),
    .o({\u2_Display/lt70_c27 ,open_n4942}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_27  (
    .a(\u2_Display/n2037 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c27 ),
    .o({\u2_Display/lt70_c28 ,open_n4943}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_28  (
    .a(\u2_Display/n2036 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c28 ),
    .o({\u2_Display/lt70_c29 ,open_n4944}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_29  (
    .a(\u2_Display/n2035 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c29 ),
    .o({\u2_Display/lt70_c30 ,open_n4945}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_3  (
    .a(\u2_Display/n2061 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c3 ),
    .o({\u2_Display/lt70_c4 ,open_n4946}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_30  (
    .a(\u2_Display/n2034 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c30 ),
    .o({\u2_Display/lt70_c31 ,open_n4947}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_31  (
    .a(\u2_Display/n2033 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c31 ),
    .o({\u2_Display/lt70_c32 ,open_n4948}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_4  (
    .a(\u2_Display/n2060 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c4 ),
    .o({\u2_Display/lt70_c5 ,open_n4949}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_5  (
    .a(\u2_Display/n2059 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c5 ),
    .o({\u2_Display/lt70_c6 ,open_n4950}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_6  (
    .a(\u2_Display/n2058 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c6 ),
    .o({\u2_Display/lt70_c7 ,open_n4951}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_7  (
    .a(\u2_Display/n2057 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c7 ),
    .o({\u2_Display/lt70_c8 ,open_n4952}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_8  (
    .a(\u2_Display/n2056 ),
    .b(1'b0),
    .c(\u2_Display/lt70_c8 ),
    .o({\u2_Display/lt70_c9 ,open_n4953}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_9  (
    .a(\u2_Display/n2055 ),
    .b(1'b1),
    .c(\u2_Display/lt70_c9 ),
    .o({\u2_Display/lt70_c10 ,open_n4954}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt70_cin  (
    .a(1'b0),
    .o({\u2_Display/lt70_c0 ,open_n4957}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt70_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt70_c32 ),
    .o({open_n4958,\u2_Display/n2065 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_0  (
    .a(\u2_Display/n2099 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c0 ),
    .o({\u2_Display/lt71_c1 ,open_n4959}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_1  (
    .a(\u2_Display/n2098 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c1 ),
    .o({\u2_Display/lt71_c2 ,open_n4960}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_10  (
    .a(\u2_Display/n2089 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c10 ),
    .o({\u2_Display/lt71_c11 ,open_n4961}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_11  (
    .a(\u2_Display/n2088 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c11 ),
    .o({\u2_Display/lt71_c12 ,open_n4962}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_12  (
    .a(\u2_Display/n2087 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c12 ),
    .o({\u2_Display/lt71_c13 ,open_n4963}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_13  (
    .a(\u2_Display/n2086 ),
    .b(1'b1),
    .c(\u2_Display/lt71_c13 ),
    .o({\u2_Display/lt71_c14 ,open_n4964}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_14  (
    .a(\u2_Display/n2085 ),
    .b(1'b1),
    .c(\u2_Display/lt71_c14 ),
    .o({\u2_Display/lt71_c15 ,open_n4965}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_15  (
    .a(\u2_Display/n2084 ),
    .b(1'b1),
    .c(\u2_Display/lt71_c15 ),
    .o({\u2_Display/lt71_c16 ,open_n4966}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_16  (
    .a(\u2_Display/n2083 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c16 ),
    .o({\u2_Display/lt71_c17 ,open_n4967}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_17  (
    .a(\u2_Display/n2082 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c17 ),
    .o({\u2_Display/lt71_c18 ,open_n4968}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_18  (
    .a(\u2_Display/n2081 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c18 ),
    .o({\u2_Display/lt71_c19 ,open_n4969}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_19  (
    .a(\u2_Display/n2080 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c19 ),
    .o({\u2_Display/lt71_c20 ,open_n4970}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_2  (
    .a(\u2_Display/n2097 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c2 ),
    .o({\u2_Display/lt71_c3 ,open_n4971}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_20  (
    .a(\u2_Display/n2079 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c20 ),
    .o({\u2_Display/lt71_c21 ,open_n4972}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_21  (
    .a(\u2_Display/n2078 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c21 ),
    .o({\u2_Display/lt71_c22 ,open_n4973}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_22  (
    .a(\u2_Display/n2077 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c22 ),
    .o({\u2_Display/lt71_c23 ,open_n4974}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_23  (
    .a(\u2_Display/n2076 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c23 ),
    .o({\u2_Display/lt71_c24 ,open_n4975}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_24  (
    .a(\u2_Display/n2075 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c24 ),
    .o({\u2_Display/lt71_c25 ,open_n4976}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_25  (
    .a(\u2_Display/n2074 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c25 ),
    .o({\u2_Display/lt71_c26 ,open_n4977}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_26  (
    .a(\u2_Display/n2073 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c26 ),
    .o({\u2_Display/lt71_c27 ,open_n4978}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_27  (
    .a(\u2_Display/n2072 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c27 ),
    .o({\u2_Display/lt71_c28 ,open_n4979}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_28  (
    .a(\u2_Display/n2071 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c28 ),
    .o({\u2_Display/lt71_c29 ,open_n4980}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_29  (
    .a(\u2_Display/n2070 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c29 ),
    .o({\u2_Display/lt71_c30 ,open_n4981}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_3  (
    .a(\u2_Display/n2096 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c3 ),
    .o({\u2_Display/lt71_c4 ,open_n4982}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_30  (
    .a(\u2_Display/n2069 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c30 ),
    .o({\u2_Display/lt71_c31 ,open_n4983}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_31  (
    .a(\u2_Display/n2068 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c31 ),
    .o({\u2_Display/lt71_c32 ,open_n4984}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_4  (
    .a(\u2_Display/n2095 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c4 ),
    .o({\u2_Display/lt71_c5 ,open_n4985}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_5  (
    .a(\u2_Display/n2094 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c5 ),
    .o({\u2_Display/lt71_c6 ,open_n4986}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_6  (
    .a(\u2_Display/n2093 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c6 ),
    .o({\u2_Display/lt71_c7 ,open_n4987}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_7  (
    .a(\u2_Display/n2092 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c7 ),
    .o({\u2_Display/lt71_c8 ,open_n4988}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_8  (
    .a(\u2_Display/n2091 ),
    .b(1'b1),
    .c(\u2_Display/lt71_c8 ),
    .o({\u2_Display/lt71_c9 ,open_n4989}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_9  (
    .a(\u2_Display/n2090 ),
    .b(1'b0),
    .c(\u2_Display/lt71_c9 ),
    .o({\u2_Display/lt71_c10 ,open_n4990}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt71_cin  (
    .a(1'b0),
    .o({\u2_Display/lt71_c0 ,open_n4993}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt71_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt71_c32 ),
    .o({open_n4994,\u2_Display/n2100 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_0  (
    .a(\u2_Display/n2134 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c0 ),
    .o({\u2_Display/lt72_c1 ,open_n4995}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_1  (
    .a(\u2_Display/n2133 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c1 ),
    .o({\u2_Display/lt72_c2 ,open_n4996}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_10  (
    .a(\u2_Display/n2124 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c10 ),
    .o({\u2_Display/lt72_c11 ,open_n4997}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_11  (
    .a(\u2_Display/n2123 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c11 ),
    .o({\u2_Display/lt72_c12 ,open_n4998}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_12  (
    .a(\u2_Display/n2122 ),
    .b(1'b1),
    .c(\u2_Display/lt72_c12 ),
    .o({\u2_Display/lt72_c13 ,open_n4999}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_13  (
    .a(\u2_Display/n2121 ),
    .b(1'b1),
    .c(\u2_Display/lt72_c13 ),
    .o({\u2_Display/lt72_c14 ,open_n5000}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_14  (
    .a(\u2_Display/n2120 ),
    .b(1'b1),
    .c(\u2_Display/lt72_c14 ),
    .o({\u2_Display/lt72_c15 ,open_n5001}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_15  (
    .a(\u2_Display/n2119 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c15 ),
    .o({\u2_Display/lt72_c16 ,open_n5002}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_16  (
    .a(\u2_Display/n2118 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c16 ),
    .o({\u2_Display/lt72_c17 ,open_n5003}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_17  (
    .a(\u2_Display/n2117 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c17 ),
    .o({\u2_Display/lt72_c18 ,open_n5004}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_18  (
    .a(\u2_Display/n2116 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c18 ),
    .o({\u2_Display/lt72_c19 ,open_n5005}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_19  (
    .a(\u2_Display/n2115 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c19 ),
    .o({\u2_Display/lt72_c20 ,open_n5006}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_2  (
    .a(\u2_Display/n2132 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c2 ),
    .o({\u2_Display/lt72_c3 ,open_n5007}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_20  (
    .a(\u2_Display/n2114 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c20 ),
    .o({\u2_Display/lt72_c21 ,open_n5008}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_21  (
    .a(\u2_Display/n2113 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c21 ),
    .o({\u2_Display/lt72_c22 ,open_n5009}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_22  (
    .a(\u2_Display/n2112 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c22 ),
    .o({\u2_Display/lt72_c23 ,open_n5010}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_23  (
    .a(\u2_Display/n2111 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c23 ),
    .o({\u2_Display/lt72_c24 ,open_n5011}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_24  (
    .a(\u2_Display/n2110 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c24 ),
    .o({\u2_Display/lt72_c25 ,open_n5012}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_25  (
    .a(\u2_Display/n2109 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c25 ),
    .o({\u2_Display/lt72_c26 ,open_n5013}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_26  (
    .a(\u2_Display/n2108 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c26 ),
    .o({\u2_Display/lt72_c27 ,open_n5014}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_27  (
    .a(\u2_Display/n2107 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c27 ),
    .o({\u2_Display/lt72_c28 ,open_n5015}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_28  (
    .a(\u2_Display/n2106 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c28 ),
    .o({\u2_Display/lt72_c29 ,open_n5016}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_29  (
    .a(\u2_Display/n2105 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c29 ),
    .o({\u2_Display/lt72_c30 ,open_n5017}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_3  (
    .a(\u2_Display/n2131 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c3 ),
    .o({\u2_Display/lt72_c4 ,open_n5018}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_30  (
    .a(\u2_Display/n2104 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c30 ),
    .o({\u2_Display/lt72_c31 ,open_n5019}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_31  (
    .a(\u2_Display/n2103 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c31 ),
    .o({\u2_Display/lt72_c32 ,open_n5020}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_4  (
    .a(\u2_Display/n2130 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c4 ),
    .o({\u2_Display/lt72_c5 ,open_n5021}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_5  (
    .a(\u2_Display/n2129 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c5 ),
    .o({\u2_Display/lt72_c6 ,open_n5022}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_6  (
    .a(\u2_Display/n2128 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c6 ),
    .o({\u2_Display/lt72_c7 ,open_n5023}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_7  (
    .a(\u2_Display/n2127 ),
    .b(1'b1),
    .c(\u2_Display/lt72_c7 ),
    .o({\u2_Display/lt72_c8 ,open_n5024}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_8  (
    .a(\u2_Display/n2126 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c8 ),
    .o({\u2_Display/lt72_c9 ,open_n5025}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_9  (
    .a(\u2_Display/n2125 ),
    .b(1'b0),
    .c(\u2_Display/lt72_c9 ),
    .o({\u2_Display/lt72_c10 ,open_n5026}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt72_cin  (
    .a(1'b0),
    .o({\u2_Display/lt72_c0 ,open_n5029}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt72_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt72_c32 ),
    .o({open_n5030,\u2_Display/n2135 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_0  (
    .a(\u2_Display/n2169 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c0 ),
    .o({\u2_Display/lt73_c1 ,open_n5031}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_1  (
    .a(\u2_Display/n2168 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c1 ),
    .o({\u2_Display/lt73_c2 ,open_n5032}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_10  (
    .a(\u2_Display/n2159 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c10 ),
    .o({\u2_Display/lt73_c11 ,open_n5033}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_11  (
    .a(\u2_Display/n2158 ),
    .b(1'b1),
    .c(\u2_Display/lt73_c11 ),
    .o({\u2_Display/lt73_c12 ,open_n5034}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_12  (
    .a(\u2_Display/n2157 ),
    .b(1'b1),
    .c(\u2_Display/lt73_c12 ),
    .o({\u2_Display/lt73_c13 ,open_n5035}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_13  (
    .a(\u2_Display/n2156 ),
    .b(1'b1),
    .c(\u2_Display/lt73_c13 ),
    .o({\u2_Display/lt73_c14 ,open_n5036}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_14  (
    .a(\u2_Display/n2155 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c14 ),
    .o({\u2_Display/lt73_c15 ,open_n5037}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_15  (
    .a(\u2_Display/n2154 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c15 ),
    .o({\u2_Display/lt73_c16 ,open_n5038}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_16  (
    .a(\u2_Display/n2153 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c16 ),
    .o({\u2_Display/lt73_c17 ,open_n5039}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_17  (
    .a(\u2_Display/n2152 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c17 ),
    .o({\u2_Display/lt73_c18 ,open_n5040}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_18  (
    .a(\u2_Display/n2151 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c18 ),
    .o({\u2_Display/lt73_c19 ,open_n5041}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_19  (
    .a(\u2_Display/n2150 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c19 ),
    .o({\u2_Display/lt73_c20 ,open_n5042}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_2  (
    .a(\u2_Display/n2167 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c2 ),
    .o({\u2_Display/lt73_c3 ,open_n5043}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_20  (
    .a(\u2_Display/n2149 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c20 ),
    .o({\u2_Display/lt73_c21 ,open_n5044}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_21  (
    .a(\u2_Display/n2148 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c21 ),
    .o({\u2_Display/lt73_c22 ,open_n5045}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_22  (
    .a(\u2_Display/n2147 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c22 ),
    .o({\u2_Display/lt73_c23 ,open_n5046}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_23  (
    .a(\u2_Display/n2146 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c23 ),
    .o({\u2_Display/lt73_c24 ,open_n5047}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_24  (
    .a(\u2_Display/n2145 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c24 ),
    .o({\u2_Display/lt73_c25 ,open_n5048}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_25  (
    .a(\u2_Display/n2144 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c25 ),
    .o({\u2_Display/lt73_c26 ,open_n5049}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_26  (
    .a(\u2_Display/n2143 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c26 ),
    .o({\u2_Display/lt73_c27 ,open_n5050}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_27  (
    .a(\u2_Display/n2142 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c27 ),
    .o({\u2_Display/lt73_c28 ,open_n5051}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_28  (
    .a(\u2_Display/n2141 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c28 ),
    .o({\u2_Display/lt73_c29 ,open_n5052}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_29  (
    .a(\u2_Display/n2140 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c29 ),
    .o({\u2_Display/lt73_c30 ,open_n5053}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_3  (
    .a(\u2_Display/n2166 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c3 ),
    .o({\u2_Display/lt73_c4 ,open_n5054}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_30  (
    .a(\u2_Display/n2139 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c30 ),
    .o({\u2_Display/lt73_c31 ,open_n5055}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_31  (
    .a(\u2_Display/n2138 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c31 ),
    .o({\u2_Display/lt73_c32 ,open_n5056}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_4  (
    .a(\u2_Display/n2165 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c4 ),
    .o({\u2_Display/lt73_c5 ,open_n5057}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_5  (
    .a(\u2_Display/n2164 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c5 ),
    .o({\u2_Display/lt73_c6 ,open_n5058}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_6  (
    .a(\u2_Display/n2163 ),
    .b(1'b1),
    .c(\u2_Display/lt73_c6 ),
    .o({\u2_Display/lt73_c7 ,open_n5059}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_7  (
    .a(\u2_Display/n2162 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c7 ),
    .o({\u2_Display/lt73_c8 ,open_n5060}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_8  (
    .a(\u2_Display/n2161 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c8 ),
    .o({\u2_Display/lt73_c9 ,open_n5061}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_9  (
    .a(\u2_Display/n2160 ),
    .b(1'b0),
    .c(\u2_Display/lt73_c9 ),
    .o({\u2_Display/lt73_c10 ,open_n5062}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt73_cin  (
    .a(1'b0),
    .o({\u2_Display/lt73_c0 ,open_n5065}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt73_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt73_c32 ),
    .o({open_n5066,\u2_Display/n2170 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_0  (
    .a(\u2_Display/n2204 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c0 ),
    .o({\u2_Display/lt74_c1 ,open_n5067}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_1  (
    .a(\u2_Display/n2203 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c1 ),
    .o({\u2_Display/lt74_c2 ,open_n5068}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_10  (
    .a(\u2_Display/n2194 ),
    .b(1'b1),
    .c(\u2_Display/lt74_c10 ),
    .o({\u2_Display/lt74_c11 ,open_n5069}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_11  (
    .a(\u2_Display/n2193 ),
    .b(1'b1),
    .c(\u2_Display/lt74_c11 ),
    .o({\u2_Display/lt74_c12 ,open_n5070}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_12  (
    .a(\u2_Display/n2192 ),
    .b(1'b1),
    .c(\u2_Display/lt74_c12 ),
    .o({\u2_Display/lt74_c13 ,open_n5071}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_13  (
    .a(\u2_Display/n2191 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c13 ),
    .o({\u2_Display/lt74_c14 ,open_n5072}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_14  (
    .a(\u2_Display/n2190 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c14 ),
    .o({\u2_Display/lt74_c15 ,open_n5073}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_15  (
    .a(\u2_Display/n2189 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c15 ),
    .o({\u2_Display/lt74_c16 ,open_n5074}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_16  (
    .a(\u2_Display/n2188 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c16 ),
    .o({\u2_Display/lt74_c17 ,open_n5075}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_17  (
    .a(\u2_Display/n2187 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c17 ),
    .o({\u2_Display/lt74_c18 ,open_n5076}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_18  (
    .a(\u2_Display/n2186 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c18 ),
    .o({\u2_Display/lt74_c19 ,open_n5077}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_19  (
    .a(\u2_Display/n2185 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c19 ),
    .o({\u2_Display/lt74_c20 ,open_n5078}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_2  (
    .a(\u2_Display/n2202 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c2 ),
    .o({\u2_Display/lt74_c3 ,open_n5079}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_20  (
    .a(\u2_Display/n2184 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c20 ),
    .o({\u2_Display/lt74_c21 ,open_n5080}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_21  (
    .a(\u2_Display/n2183 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c21 ),
    .o({\u2_Display/lt74_c22 ,open_n5081}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_22  (
    .a(\u2_Display/n2182 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c22 ),
    .o({\u2_Display/lt74_c23 ,open_n5082}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_23  (
    .a(\u2_Display/n2181 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c23 ),
    .o({\u2_Display/lt74_c24 ,open_n5083}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_24  (
    .a(\u2_Display/n2180 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c24 ),
    .o({\u2_Display/lt74_c25 ,open_n5084}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_25  (
    .a(\u2_Display/n2179 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c25 ),
    .o({\u2_Display/lt74_c26 ,open_n5085}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_26  (
    .a(\u2_Display/n2178 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c26 ),
    .o({\u2_Display/lt74_c27 ,open_n5086}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_27  (
    .a(\u2_Display/n2177 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c27 ),
    .o({\u2_Display/lt74_c28 ,open_n5087}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_28  (
    .a(\u2_Display/n2176 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c28 ),
    .o({\u2_Display/lt74_c29 ,open_n5088}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_29  (
    .a(\u2_Display/n2175 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c29 ),
    .o({\u2_Display/lt74_c30 ,open_n5089}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_3  (
    .a(\u2_Display/n2201 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c3 ),
    .o({\u2_Display/lt74_c4 ,open_n5090}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_30  (
    .a(\u2_Display/n2174 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c30 ),
    .o({\u2_Display/lt74_c31 ,open_n5091}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_31  (
    .a(\u2_Display/n2173 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c31 ),
    .o({\u2_Display/lt74_c32 ,open_n5092}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_4  (
    .a(\u2_Display/n2200 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c4 ),
    .o({\u2_Display/lt74_c5 ,open_n5093}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_5  (
    .a(\u2_Display/n2199 ),
    .b(1'b1),
    .c(\u2_Display/lt74_c5 ),
    .o({\u2_Display/lt74_c6 ,open_n5094}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_6  (
    .a(\u2_Display/n2198 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c6 ),
    .o({\u2_Display/lt74_c7 ,open_n5095}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_7  (
    .a(\u2_Display/n2197 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c7 ),
    .o({\u2_Display/lt74_c8 ,open_n5096}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_8  (
    .a(\u2_Display/n2196 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c8 ),
    .o({\u2_Display/lt74_c9 ,open_n5097}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_9  (
    .a(\u2_Display/n2195 ),
    .b(1'b0),
    .c(\u2_Display/lt74_c9 ),
    .o({\u2_Display/lt74_c10 ,open_n5098}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt74_cin  (
    .a(1'b0),
    .o({\u2_Display/lt74_c0 ,open_n5101}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt74_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt74_c32 ),
    .o({open_n5102,\u2_Display/n2205 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_0  (
    .a(\u2_Display/n2239 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c0 ),
    .o({\u2_Display/lt75_c1 ,open_n5103}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_1  (
    .a(\u2_Display/n2238 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c1 ),
    .o({\u2_Display/lt75_c2 ,open_n5104}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_10  (
    .a(\u2_Display/n2229 ),
    .b(1'b1),
    .c(\u2_Display/lt75_c10 ),
    .o({\u2_Display/lt75_c11 ,open_n5105}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_11  (
    .a(\u2_Display/n2228 ),
    .b(1'b1),
    .c(\u2_Display/lt75_c11 ),
    .o({\u2_Display/lt75_c12 ,open_n5106}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_12  (
    .a(\u2_Display/n2227 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c12 ),
    .o({\u2_Display/lt75_c13 ,open_n5107}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_13  (
    .a(\u2_Display/n2226 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c13 ),
    .o({\u2_Display/lt75_c14 ,open_n5108}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_14  (
    .a(\u2_Display/n2225 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c14 ),
    .o({\u2_Display/lt75_c15 ,open_n5109}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_15  (
    .a(\u2_Display/n2224 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c15 ),
    .o({\u2_Display/lt75_c16 ,open_n5110}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_16  (
    .a(\u2_Display/n2223 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c16 ),
    .o({\u2_Display/lt75_c17 ,open_n5111}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_17  (
    .a(\u2_Display/n2222 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c17 ),
    .o({\u2_Display/lt75_c18 ,open_n5112}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_18  (
    .a(\u2_Display/n2221 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c18 ),
    .o({\u2_Display/lt75_c19 ,open_n5113}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_19  (
    .a(\u2_Display/n2220 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c19 ),
    .o({\u2_Display/lt75_c20 ,open_n5114}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_2  (
    .a(\u2_Display/n2237 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c2 ),
    .o({\u2_Display/lt75_c3 ,open_n5115}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_20  (
    .a(\u2_Display/n2219 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c20 ),
    .o({\u2_Display/lt75_c21 ,open_n5116}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_21  (
    .a(\u2_Display/n2218 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c21 ),
    .o({\u2_Display/lt75_c22 ,open_n5117}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_22  (
    .a(\u2_Display/n2217 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c22 ),
    .o({\u2_Display/lt75_c23 ,open_n5118}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_23  (
    .a(\u2_Display/n2216 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c23 ),
    .o({\u2_Display/lt75_c24 ,open_n5119}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_24  (
    .a(\u2_Display/n2215 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c24 ),
    .o({\u2_Display/lt75_c25 ,open_n5120}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_25  (
    .a(\u2_Display/n2214 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c25 ),
    .o({\u2_Display/lt75_c26 ,open_n5121}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_26  (
    .a(\u2_Display/n2213 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c26 ),
    .o({\u2_Display/lt75_c27 ,open_n5122}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_27  (
    .a(\u2_Display/n2212 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c27 ),
    .o({\u2_Display/lt75_c28 ,open_n5123}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_28  (
    .a(\u2_Display/n2211 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c28 ),
    .o({\u2_Display/lt75_c29 ,open_n5124}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_29  (
    .a(\u2_Display/n2210 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c29 ),
    .o({\u2_Display/lt75_c30 ,open_n5125}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_3  (
    .a(\u2_Display/n2236 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c3 ),
    .o({\u2_Display/lt75_c4 ,open_n5126}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_30  (
    .a(\u2_Display/n2209 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c30 ),
    .o({\u2_Display/lt75_c31 ,open_n5127}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_31  (
    .a(\u2_Display/n2208 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c31 ),
    .o({\u2_Display/lt75_c32 ,open_n5128}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_4  (
    .a(\u2_Display/n2235 ),
    .b(1'b1),
    .c(\u2_Display/lt75_c4 ),
    .o({\u2_Display/lt75_c5 ,open_n5129}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_5  (
    .a(\u2_Display/n2234 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c5 ),
    .o({\u2_Display/lt75_c6 ,open_n5130}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_6  (
    .a(\u2_Display/n2233 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c6 ),
    .o({\u2_Display/lt75_c7 ,open_n5131}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_7  (
    .a(\u2_Display/n2232 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c7 ),
    .o({\u2_Display/lt75_c8 ,open_n5132}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_8  (
    .a(\u2_Display/n2231 ),
    .b(1'b0),
    .c(\u2_Display/lt75_c8 ),
    .o({\u2_Display/lt75_c9 ,open_n5133}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_9  (
    .a(\u2_Display/n2230 ),
    .b(1'b1),
    .c(\u2_Display/lt75_c9 ),
    .o({\u2_Display/lt75_c10 ,open_n5134}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt75_cin  (
    .a(1'b0),
    .o({\u2_Display/lt75_c0 ,open_n5137}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt75_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt75_c32 ),
    .o({open_n5138,\u2_Display/n2240 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_0  (
    .a(\u2_Display/n2274 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c0 ),
    .o({\u2_Display/lt76_c1 ,open_n5139}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_1  (
    .a(\u2_Display/n2273 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c1 ),
    .o({\u2_Display/lt76_c2 ,open_n5140}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_10  (
    .a(\u2_Display/n2264 ),
    .b(1'b1),
    .c(\u2_Display/lt76_c10 ),
    .o({\u2_Display/lt76_c11 ,open_n5141}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_11  (
    .a(\u2_Display/n2263 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c11 ),
    .o({\u2_Display/lt76_c12 ,open_n5142}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_12  (
    .a(\u2_Display/n2262 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c12 ),
    .o({\u2_Display/lt76_c13 ,open_n5143}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_13  (
    .a(\u2_Display/n2261 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c13 ),
    .o({\u2_Display/lt76_c14 ,open_n5144}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_14  (
    .a(\u2_Display/n2260 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c14 ),
    .o({\u2_Display/lt76_c15 ,open_n5145}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_15  (
    .a(\u2_Display/n2259 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c15 ),
    .o({\u2_Display/lt76_c16 ,open_n5146}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_16  (
    .a(\u2_Display/n2258 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c16 ),
    .o({\u2_Display/lt76_c17 ,open_n5147}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_17  (
    .a(\u2_Display/n2257 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c17 ),
    .o({\u2_Display/lt76_c18 ,open_n5148}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_18  (
    .a(\u2_Display/n2256 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c18 ),
    .o({\u2_Display/lt76_c19 ,open_n5149}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_19  (
    .a(\u2_Display/n2255 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c19 ),
    .o({\u2_Display/lt76_c20 ,open_n5150}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_2  (
    .a(\u2_Display/n2272 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c2 ),
    .o({\u2_Display/lt76_c3 ,open_n5151}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_20  (
    .a(\u2_Display/n2254 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c20 ),
    .o({\u2_Display/lt76_c21 ,open_n5152}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_21  (
    .a(\u2_Display/n2253 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c21 ),
    .o({\u2_Display/lt76_c22 ,open_n5153}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_22  (
    .a(\u2_Display/n2252 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c22 ),
    .o({\u2_Display/lt76_c23 ,open_n5154}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_23  (
    .a(\u2_Display/n2251 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c23 ),
    .o({\u2_Display/lt76_c24 ,open_n5155}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_24  (
    .a(\u2_Display/n2250 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c24 ),
    .o({\u2_Display/lt76_c25 ,open_n5156}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_25  (
    .a(\u2_Display/n2249 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c25 ),
    .o({\u2_Display/lt76_c26 ,open_n5157}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_26  (
    .a(\u2_Display/n2248 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c26 ),
    .o({\u2_Display/lt76_c27 ,open_n5158}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_27  (
    .a(\u2_Display/n2247 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c27 ),
    .o({\u2_Display/lt76_c28 ,open_n5159}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_28  (
    .a(\u2_Display/n2246 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c28 ),
    .o({\u2_Display/lt76_c29 ,open_n5160}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_29  (
    .a(\u2_Display/n2245 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c29 ),
    .o({\u2_Display/lt76_c30 ,open_n5161}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_3  (
    .a(\u2_Display/n2271 ),
    .b(1'b1),
    .c(\u2_Display/lt76_c3 ),
    .o({\u2_Display/lt76_c4 ,open_n5162}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_30  (
    .a(\u2_Display/n2244 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c30 ),
    .o({\u2_Display/lt76_c31 ,open_n5163}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_31  (
    .a(\u2_Display/n2243 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c31 ),
    .o({\u2_Display/lt76_c32 ,open_n5164}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_4  (
    .a(\u2_Display/n2270 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c4 ),
    .o({\u2_Display/lt76_c5 ,open_n5165}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_5  (
    .a(\u2_Display/n2269 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c5 ),
    .o({\u2_Display/lt76_c6 ,open_n5166}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_6  (
    .a(\u2_Display/n2268 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c6 ),
    .o({\u2_Display/lt76_c7 ,open_n5167}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_7  (
    .a(\u2_Display/n2267 ),
    .b(1'b0),
    .c(\u2_Display/lt76_c7 ),
    .o({\u2_Display/lt76_c8 ,open_n5168}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_8  (
    .a(\u2_Display/n2266 ),
    .b(1'b1),
    .c(\u2_Display/lt76_c8 ),
    .o({\u2_Display/lt76_c9 ,open_n5169}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_9  (
    .a(\u2_Display/n2265 ),
    .b(1'b1),
    .c(\u2_Display/lt76_c9 ),
    .o({\u2_Display/lt76_c10 ,open_n5170}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt76_cin  (
    .a(1'b0),
    .o({\u2_Display/lt76_c0 ,open_n5173}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt76_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt76_c32 ),
    .o({open_n5174,\u2_Display/n2275 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_0  (
    .a(\u2_Display/n2309 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c0 ),
    .o({\u2_Display/lt77_c1 ,open_n5175}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_1  (
    .a(\u2_Display/n2308 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c1 ),
    .o({\u2_Display/lt77_c2 ,open_n5176}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_10  (
    .a(\u2_Display/n2299 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c10 ),
    .o({\u2_Display/lt77_c11 ,open_n5177}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_11  (
    .a(\u2_Display/n2298 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c11 ),
    .o({\u2_Display/lt77_c12 ,open_n5178}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_12  (
    .a(\u2_Display/n2297 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c12 ),
    .o({\u2_Display/lt77_c13 ,open_n5179}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_13  (
    .a(\u2_Display/n2296 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c13 ),
    .o({\u2_Display/lt77_c14 ,open_n5180}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_14  (
    .a(\u2_Display/n2295 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c14 ),
    .o({\u2_Display/lt77_c15 ,open_n5181}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_15  (
    .a(\u2_Display/n2294 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c15 ),
    .o({\u2_Display/lt77_c16 ,open_n5182}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_16  (
    .a(\u2_Display/n2293 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c16 ),
    .o({\u2_Display/lt77_c17 ,open_n5183}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_17  (
    .a(\u2_Display/n2292 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c17 ),
    .o({\u2_Display/lt77_c18 ,open_n5184}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_18  (
    .a(\u2_Display/n2291 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c18 ),
    .o({\u2_Display/lt77_c19 ,open_n5185}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_19  (
    .a(\u2_Display/n2290 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c19 ),
    .o({\u2_Display/lt77_c20 ,open_n5186}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_2  (
    .a(\u2_Display/n2307 ),
    .b(1'b1),
    .c(\u2_Display/lt77_c2 ),
    .o({\u2_Display/lt77_c3 ,open_n5187}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_20  (
    .a(\u2_Display/n2289 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c20 ),
    .o({\u2_Display/lt77_c21 ,open_n5188}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_21  (
    .a(\u2_Display/n2288 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c21 ),
    .o({\u2_Display/lt77_c22 ,open_n5189}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_22  (
    .a(\u2_Display/n2287 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c22 ),
    .o({\u2_Display/lt77_c23 ,open_n5190}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_23  (
    .a(\u2_Display/n2286 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c23 ),
    .o({\u2_Display/lt77_c24 ,open_n5191}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_24  (
    .a(\u2_Display/n2285 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c24 ),
    .o({\u2_Display/lt77_c25 ,open_n5192}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_25  (
    .a(\u2_Display/n2284 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c25 ),
    .o({\u2_Display/lt77_c26 ,open_n5193}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_26  (
    .a(\u2_Display/n2283 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c26 ),
    .o({\u2_Display/lt77_c27 ,open_n5194}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_27  (
    .a(\u2_Display/n2282 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c27 ),
    .o({\u2_Display/lt77_c28 ,open_n5195}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_28  (
    .a(\u2_Display/n2281 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c28 ),
    .o({\u2_Display/lt77_c29 ,open_n5196}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_29  (
    .a(\u2_Display/n2280 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c29 ),
    .o({\u2_Display/lt77_c30 ,open_n5197}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_3  (
    .a(\u2_Display/n2306 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c3 ),
    .o({\u2_Display/lt77_c4 ,open_n5198}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_30  (
    .a(\u2_Display/n2279 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c30 ),
    .o({\u2_Display/lt77_c31 ,open_n5199}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_31  (
    .a(\u2_Display/n2278 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c31 ),
    .o({\u2_Display/lt77_c32 ,open_n5200}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_4  (
    .a(\u2_Display/n2305 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c4 ),
    .o({\u2_Display/lt77_c5 ,open_n5201}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_5  (
    .a(\u2_Display/n2304 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c5 ),
    .o({\u2_Display/lt77_c6 ,open_n5202}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_6  (
    .a(\u2_Display/n2303 ),
    .b(1'b0),
    .c(\u2_Display/lt77_c6 ),
    .o({\u2_Display/lt77_c7 ,open_n5203}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_7  (
    .a(\u2_Display/n2302 ),
    .b(1'b1),
    .c(\u2_Display/lt77_c7 ),
    .o({\u2_Display/lt77_c8 ,open_n5204}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_8  (
    .a(\u2_Display/n2301 ),
    .b(1'b1),
    .c(\u2_Display/lt77_c8 ),
    .o({\u2_Display/lt77_c9 ,open_n5205}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_9  (
    .a(\u2_Display/n2300 ),
    .b(1'b1),
    .c(\u2_Display/lt77_c9 ),
    .o({\u2_Display/lt77_c10 ,open_n5206}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt77_cin  (
    .a(1'b0),
    .o({\u2_Display/lt77_c0 ,open_n5209}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt77_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt77_c32 ),
    .o({open_n5210,\u2_Display/n2310 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_0  (
    .a(\u2_Display/n102 [0]),
    .b(lcd_ypos[0]),
    .c(\u2_Display/lt7_2_c0 ),
    .o({\u2_Display/lt7_2_c1 ,open_n5211}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_1  (
    .a(\u2_Display/n102 [1]),
    .b(lcd_ypos[1]),
    .c(\u2_Display/lt7_2_c1 ),
    .o({\u2_Display/lt7_2_c2 ,open_n5212}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_10  (
    .a(\u2_Display/n102 [31]),
    .b(lcd_ypos[10]),
    .c(\u2_Display/lt7_2_c10 ),
    .o({\u2_Display/lt7_2_c11 ,open_n5213}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_11  (
    .a(\u2_Display/n102 [31]),
    .b(lcd_ypos[11]),
    .c(\u2_Display/lt7_2_c11 ),
    .o({\u2_Display/lt7_2_c12 ,open_n5214}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_12  (
    .a(\u2_Display/n102 [31]),
    .b(1'b0),
    .c(\u2_Display/lt7_2_c12 ),
    .o({\u2_Display/lt7_2_c13 ,open_n5215}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_2  (
    .a(\u2_Display/n102 [2]),
    .b(lcd_ypos[2]),
    .c(\u2_Display/lt7_2_c2 ),
    .o({\u2_Display/lt7_2_c3 ,open_n5216}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_3  (
    .a(\u2_Display/n102 [3]),
    .b(lcd_ypos[3]),
    .c(\u2_Display/lt7_2_c3 ),
    .o({\u2_Display/lt7_2_c4 ,open_n5217}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_4  (
    .a(\u2_Display/n102 [4]),
    .b(lcd_ypos[4]),
    .c(\u2_Display/lt7_2_c4 ),
    .o({\u2_Display/lt7_2_c5 ,open_n5218}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_5  (
    .a(\u2_Display/n102 [5]),
    .b(lcd_ypos[5]),
    .c(\u2_Display/lt7_2_c5 ),
    .o({\u2_Display/lt7_2_c6 ,open_n5219}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_6  (
    .a(\u2_Display/n102 [6]),
    .b(lcd_ypos[6]),
    .c(\u2_Display/lt7_2_c6 ),
    .o({\u2_Display/lt7_2_c7 ,open_n5220}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_7  (
    .a(\u2_Display/n102 [7]),
    .b(lcd_ypos[7]),
    .c(\u2_Display/lt7_2_c7 ),
    .o({\u2_Display/lt7_2_c8 ,open_n5221}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_8  (
    .a(\u2_Display/n102 [8]),
    .b(lcd_ypos[8]),
    .c(\u2_Display/lt7_2_c8 ),
    .o({\u2_Display/lt7_2_c9 ,open_n5222}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_9  (
    .a(\u2_Display/n102 [9]),
    .b(lcd_ypos[9]),
    .c(\u2_Display/lt7_2_c9 ),
    .o({\u2_Display/lt7_2_c10 ,open_n5223}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt7_2_cin  (
    .a(1'b0),
    .o({\u2_Display/lt7_2_c0 ,open_n5226}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt7_2_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt7_2_c13 ),
    .o({open_n5227,\u2_Display/n103 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_0  (
    .a(\u2_Display/counta [0]),
    .b(1'b0),
    .c(\u2_Display/lt88_c0 ),
    .o({\u2_Display/lt88_c1 ,open_n5228}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_1  (
    .a(\u2_Display/counta [1]),
    .b(1'b0),
    .c(\u2_Display/lt88_c1 ),
    .o({\u2_Display/lt88_c2 ,open_n5229}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_10  (
    .a(\u2_Display/counta [10]),
    .b(1'b0),
    .c(\u2_Display/lt88_c10 ),
    .o({\u2_Display/lt88_c11 ,open_n5230}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_11  (
    .a(\u2_Display/counta [11]),
    .b(1'b0),
    .c(\u2_Display/lt88_c11 ),
    .o({\u2_Display/lt88_c12 ,open_n5231}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_12  (
    .a(\u2_Display/counta [12]),
    .b(1'b0),
    .c(\u2_Display/lt88_c12 ),
    .o({\u2_Display/lt88_c13 ,open_n5232}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_13  (
    .a(\u2_Display/counta [13]),
    .b(1'b0),
    .c(\u2_Display/lt88_c13 ),
    .o({\u2_Display/lt88_c14 ,open_n5233}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_14  (
    .a(\u2_Display/counta [14]),
    .b(1'b0),
    .c(\u2_Display/lt88_c14 ),
    .o({\u2_Display/lt88_c15 ,open_n5234}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_15  (
    .a(\u2_Display/counta [15]),
    .b(1'b0),
    .c(\u2_Display/lt88_c15 ),
    .o({\u2_Display/lt88_c16 ,open_n5235}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_16  (
    .a(\u2_Display/counta [16]),
    .b(1'b0),
    .c(\u2_Display/lt88_c16 ),
    .o({\u2_Display/lt88_c17 ,open_n5236}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_17  (
    .a(\u2_Display/counta [17]),
    .b(1'b0),
    .c(\u2_Display/lt88_c17 ),
    .o({\u2_Display/lt88_c18 ,open_n5237}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_18  (
    .a(\u2_Display/counta [18]),
    .b(1'b0),
    .c(\u2_Display/lt88_c18 ),
    .o({\u2_Display/lt88_c19 ,open_n5238}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_19  (
    .a(\u2_Display/counta [19]),
    .b(1'b0),
    .c(\u2_Display/lt88_c19 ),
    .o({\u2_Display/lt88_c20 ,open_n5239}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_2  (
    .a(\u2_Display/counta [2]),
    .b(1'b0),
    .c(\u2_Display/lt88_c2 ),
    .o({\u2_Display/lt88_c3 ,open_n5240}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_20  (
    .a(\u2_Display/counta [20]),
    .b(1'b0),
    .c(\u2_Display/lt88_c20 ),
    .o({\u2_Display/lt88_c21 ,open_n5241}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_21  (
    .a(\u2_Display/counta [21]),
    .b(1'b0),
    .c(\u2_Display/lt88_c21 ),
    .o({\u2_Display/lt88_c22 ,open_n5242}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_22  (
    .a(\u2_Display/counta [22]),
    .b(1'b0),
    .c(\u2_Display/lt88_c22 ),
    .o({\u2_Display/lt88_c23 ,open_n5243}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_23  (
    .a(\u2_Display/counta [23]),
    .b(1'b0),
    .c(\u2_Display/lt88_c23 ),
    .o({\u2_Display/lt88_c24 ,open_n5244}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_24  (
    .a(\u2_Display/counta [24]),
    .b(1'b0),
    .c(\u2_Display/lt88_c24 ),
    .o({\u2_Display/lt88_c25 ,open_n5245}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_25  (
    .a(\u2_Display/counta [25]),
    .b(1'b1),
    .c(\u2_Display/lt88_c25 ),
    .o({\u2_Display/lt88_c26 ,open_n5246}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_26  (
    .a(\u2_Display/counta [26]),
    .b(1'b1),
    .c(\u2_Display/lt88_c26 ),
    .o({\u2_Display/lt88_c27 ,open_n5247}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_27  (
    .a(\u2_Display/counta [27]),
    .b(1'b0),
    .c(\u2_Display/lt88_c27 ),
    .o({\u2_Display/lt88_c28 ,open_n5248}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_28  (
    .a(\u2_Display/counta [28]),
    .b(1'b1),
    .c(\u2_Display/lt88_c28 ),
    .o({\u2_Display/lt88_c29 ,open_n5249}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_29  (
    .a(\u2_Display/counta [29]),
    .b(1'b0),
    .c(\u2_Display/lt88_c29 ),
    .o({\u2_Display/lt88_c30 ,open_n5250}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_3  (
    .a(\u2_Display/counta [3]),
    .b(1'b0),
    .c(\u2_Display/lt88_c3 ),
    .o({\u2_Display/lt88_c4 ,open_n5251}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_30  (
    .a(\u2_Display/counta [30]),
    .b(1'b0),
    .c(\u2_Display/lt88_c30 ),
    .o({\u2_Display/lt88_c31 ,open_n5252}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_31  (
    .a(\u2_Display/counta [31]),
    .b(1'b1),
    .c(\u2_Display/lt88_c31 ),
    .o({\u2_Display/lt88_c32 ,open_n5253}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_4  (
    .a(\u2_Display/counta [4]),
    .b(1'b0),
    .c(\u2_Display/lt88_c4 ),
    .o({\u2_Display/lt88_c5 ,open_n5254}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_5  (
    .a(\u2_Display/counta [5]),
    .b(1'b0),
    .c(\u2_Display/lt88_c5 ),
    .o({\u2_Display/lt88_c6 ,open_n5255}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_6  (
    .a(\u2_Display/counta [6]),
    .b(1'b0),
    .c(\u2_Display/lt88_c6 ),
    .o({\u2_Display/lt88_c7 ,open_n5256}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_7  (
    .a(\u2_Display/counta [7]),
    .b(1'b0),
    .c(\u2_Display/lt88_c7 ),
    .o({\u2_Display/lt88_c8 ,open_n5257}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_8  (
    .a(\u2_Display/counta [8]),
    .b(1'b0),
    .c(\u2_Display/lt88_c8 ),
    .o({\u2_Display/lt88_c9 ,open_n5258}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_9  (
    .a(\u2_Display/counta [9]),
    .b(1'b0),
    .c(\u2_Display/lt88_c9 ),
    .o({\u2_Display/lt88_c10 ,open_n5259}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt88_cin  (
    .a(1'b0),
    .o({\u2_Display/lt88_c0 ,open_n5262}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt88_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt88_c32 ),
    .o({open_n5263,\u2_Display/n2663 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_0  (
    .a(\u2_Display/n2697 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c0 ),
    .o({\u2_Display/lt89_c1 ,open_n5264}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_1  (
    .a(\u2_Display/n2696 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c1 ),
    .o({\u2_Display/lt89_c2 ,open_n5265}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_10  (
    .a(\u2_Display/n2687 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c10 ),
    .o({\u2_Display/lt89_c11 ,open_n5266}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_11  (
    .a(\u2_Display/n2686 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c11 ),
    .o({\u2_Display/lt89_c12 ,open_n5267}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_12  (
    .a(\u2_Display/n2685 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c12 ),
    .o({\u2_Display/lt89_c13 ,open_n5268}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_13  (
    .a(\u2_Display/n2684 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c13 ),
    .o({\u2_Display/lt89_c14 ,open_n5269}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_14  (
    .a(\u2_Display/n2683 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c14 ),
    .o({\u2_Display/lt89_c15 ,open_n5270}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_15  (
    .a(\u2_Display/n2682 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c15 ),
    .o({\u2_Display/lt89_c16 ,open_n5271}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_16  (
    .a(\u2_Display/n2681 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c16 ),
    .o({\u2_Display/lt89_c17 ,open_n5272}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_17  (
    .a(\u2_Display/n2680 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c17 ),
    .o({\u2_Display/lt89_c18 ,open_n5273}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_18  (
    .a(\u2_Display/n2679 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c18 ),
    .o({\u2_Display/lt89_c19 ,open_n5274}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_19  (
    .a(\u2_Display/n2678 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c19 ),
    .o({\u2_Display/lt89_c20 ,open_n5275}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_2  (
    .a(\u2_Display/n2695 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c2 ),
    .o({\u2_Display/lt89_c3 ,open_n5276}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_20  (
    .a(\u2_Display/n2677 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c20 ),
    .o({\u2_Display/lt89_c21 ,open_n5277}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_21  (
    .a(\u2_Display/n2676 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c21 ),
    .o({\u2_Display/lt89_c22 ,open_n5278}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_22  (
    .a(\u2_Display/n2675 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c22 ),
    .o({\u2_Display/lt89_c23 ,open_n5279}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_23  (
    .a(\u2_Display/n2674 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c23 ),
    .o({\u2_Display/lt89_c24 ,open_n5280}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_24  (
    .a(\u2_Display/n2673 ),
    .b(1'b1),
    .c(\u2_Display/lt89_c24 ),
    .o({\u2_Display/lt89_c25 ,open_n5281}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_25  (
    .a(\u2_Display/n2672 ),
    .b(1'b1),
    .c(\u2_Display/lt89_c25 ),
    .o({\u2_Display/lt89_c26 ,open_n5282}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_26  (
    .a(\u2_Display/n2671 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c26 ),
    .o({\u2_Display/lt89_c27 ,open_n5283}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_27  (
    .a(\u2_Display/n2670 ),
    .b(1'b1),
    .c(\u2_Display/lt89_c27 ),
    .o({\u2_Display/lt89_c28 ,open_n5284}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_28  (
    .a(\u2_Display/n2669 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c28 ),
    .o({\u2_Display/lt89_c29 ,open_n5285}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_29  (
    .a(\u2_Display/n2668 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c29 ),
    .o({\u2_Display/lt89_c30 ,open_n5286}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_3  (
    .a(\u2_Display/n2694 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c3 ),
    .o({\u2_Display/lt89_c4 ,open_n5287}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_30  (
    .a(\u2_Display/n2667 ),
    .b(1'b1),
    .c(\u2_Display/lt89_c30 ),
    .o({\u2_Display/lt89_c31 ,open_n5288}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_31  (
    .a(\u2_Display/n2666 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c31 ),
    .o({\u2_Display/lt89_c32 ,open_n5289}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_4  (
    .a(\u2_Display/n2693 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c4 ),
    .o({\u2_Display/lt89_c5 ,open_n5290}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_5  (
    .a(\u2_Display/n2692 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c5 ),
    .o({\u2_Display/lt89_c6 ,open_n5291}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_6  (
    .a(\u2_Display/n2691 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c6 ),
    .o({\u2_Display/lt89_c7 ,open_n5292}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_7  (
    .a(\u2_Display/n2690 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c7 ),
    .o({\u2_Display/lt89_c8 ,open_n5293}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_8  (
    .a(\u2_Display/n2689 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c8 ),
    .o({\u2_Display/lt89_c9 ,open_n5294}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_9  (
    .a(\u2_Display/n2688 ),
    .b(1'b0),
    .c(\u2_Display/lt89_c9 ),
    .o({\u2_Display/lt89_c10 ,open_n5295}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt89_cin  (
    .a(1'b0),
    .o({\u2_Display/lt89_c0 ,open_n5298}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt89_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt89_c32 ),
    .o({open_n5299,\u2_Display/n2698 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt8_2_0  (
    .a(lcd_xpos[0]),
    .b(\u2_Display/j [0]),
    .c(\u2_Display/lt8_2_c0 ),
    .o({\u2_Display/lt8_2_c1 ,open_n5300}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt8_2_1  (
    .a(lcd_xpos[1]),
    .b(\u2_Display/j [1]),
    .c(\u2_Display/lt8_2_c1 ),
    .o({\u2_Display/lt8_2_c2 ,open_n5301}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt8_2_10  (
    .a(lcd_xpos[10]),
    .b(\u2_Display/add6_2_co ),
    .c(\u2_Display/lt8_2_c10 ),
    .o({\u2_Display/lt8_2_c11 ,open_n5302}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt8_2_11  (
    .a(lcd_xpos[11]),
    .b(1'b0),
    .c(\u2_Display/lt8_2_c11 ),
    .o({\u2_Display/lt8_2_c12 ,open_n5303}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt8_2_2  (
    .a(lcd_xpos[2]),
    .b(\u2_Display/j [2]),
    .c(\u2_Display/lt8_2_c2 ),
    .o({\u2_Display/lt8_2_c3 ,open_n5304}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt8_2_3  (
    .a(lcd_xpos[3]),
    .b(\u2_Display/j [3]),
    .c(\u2_Display/lt8_2_c3 ),
    .o({\u2_Display/lt8_2_c4 ,open_n5305}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt8_2_4  (
    .a(lcd_xpos[4]),
    .b(\u2_Display/j [4]),
    .c(\u2_Display/lt8_2_c4 ),
    .o({\u2_Display/lt8_2_c5 ,open_n5306}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt8_2_5  (
    .a(lcd_xpos[5]),
    .b(\u2_Display/j [5]),
    .c(\u2_Display/lt8_2_c5 ),
    .o({\u2_Display/lt8_2_c6 ,open_n5307}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt8_2_6  (
    .a(lcd_xpos[6]),
    .b(\u2_Display/j [6]),
    .c(\u2_Display/lt8_2_c6 ),
    .o({\u2_Display/lt8_2_c7 ,open_n5308}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt8_2_7  (
    .a(lcd_xpos[7]),
    .b(\u2_Display/n135 [0]),
    .c(\u2_Display/lt8_2_c7 ),
    .o({\u2_Display/lt8_2_c8 ,open_n5309}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt8_2_8  (
    .a(lcd_xpos[8]),
    .b(\u2_Display/n135 [1]),
    .c(\u2_Display/lt8_2_c8 ),
    .o({\u2_Display/lt8_2_c9 ,open_n5310}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt8_2_9  (
    .a(lcd_xpos[9]),
    .b(\u2_Display/n135 [2]),
    .c(\u2_Display/lt8_2_c9 ),
    .o({\u2_Display/lt8_2_c10 ,open_n5311}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt8_2_cin  (
    .a(1'b0),
    .o({\u2_Display/lt8_2_c0 ,open_n5314}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt8_2_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt8_2_c12 ),
    .o({open_n5315,\u2_Display/n136 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_0  (
    .a(\u2_Display/n2732 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c0 ),
    .o({\u2_Display/lt90_c1 ,open_n5316}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_1  (
    .a(\u2_Display/n2731 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c1 ),
    .o({\u2_Display/lt90_c2 ,open_n5317}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_10  (
    .a(\u2_Display/n2722 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c10 ),
    .o({\u2_Display/lt90_c11 ,open_n5318}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_11  (
    .a(\u2_Display/n2721 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c11 ),
    .o({\u2_Display/lt90_c12 ,open_n5319}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_12  (
    .a(\u2_Display/n2720 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c12 ),
    .o({\u2_Display/lt90_c13 ,open_n5320}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_13  (
    .a(\u2_Display/n2719 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c13 ),
    .o({\u2_Display/lt90_c14 ,open_n5321}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_14  (
    .a(\u2_Display/n2718 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c14 ),
    .o({\u2_Display/lt90_c15 ,open_n5322}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_15  (
    .a(\u2_Display/n2717 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c15 ),
    .o({\u2_Display/lt90_c16 ,open_n5323}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_16  (
    .a(\u2_Display/n2716 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c16 ),
    .o({\u2_Display/lt90_c17 ,open_n5324}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_17  (
    .a(\u2_Display/n2715 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c17 ),
    .o({\u2_Display/lt90_c18 ,open_n5325}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_18  (
    .a(\u2_Display/n2714 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c18 ),
    .o({\u2_Display/lt90_c19 ,open_n5326}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_19  (
    .a(\u2_Display/n2713 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c19 ),
    .o({\u2_Display/lt90_c20 ,open_n5327}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_2  (
    .a(\u2_Display/n2730 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c2 ),
    .o({\u2_Display/lt90_c3 ,open_n5328}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_20  (
    .a(\u2_Display/n2712 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c20 ),
    .o({\u2_Display/lt90_c21 ,open_n5329}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_21  (
    .a(\u2_Display/n2711 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c21 ),
    .o({\u2_Display/lt90_c22 ,open_n5330}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_22  (
    .a(\u2_Display/n2710 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c22 ),
    .o({\u2_Display/lt90_c23 ,open_n5331}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_23  (
    .a(\u2_Display/n2709 ),
    .b(1'b1),
    .c(\u2_Display/lt90_c23 ),
    .o({\u2_Display/lt90_c24 ,open_n5332}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_24  (
    .a(\u2_Display/n2708 ),
    .b(1'b1),
    .c(\u2_Display/lt90_c24 ),
    .o({\u2_Display/lt90_c25 ,open_n5333}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_25  (
    .a(\u2_Display/n2707 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c25 ),
    .o({\u2_Display/lt90_c26 ,open_n5334}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_26  (
    .a(\u2_Display/n2706 ),
    .b(1'b1),
    .c(\u2_Display/lt90_c26 ),
    .o({\u2_Display/lt90_c27 ,open_n5335}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_27  (
    .a(\u2_Display/n2705 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c27 ),
    .o({\u2_Display/lt90_c28 ,open_n5336}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_28  (
    .a(\u2_Display/n2704 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c28 ),
    .o({\u2_Display/lt90_c29 ,open_n5337}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_29  (
    .a(\u2_Display/n2703 ),
    .b(1'b1),
    .c(\u2_Display/lt90_c29 ),
    .o({\u2_Display/lt90_c30 ,open_n5338}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_3  (
    .a(\u2_Display/n2729 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c3 ),
    .o({\u2_Display/lt90_c4 ,open_n5339}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_30  (
    .a(\u2_Display/n2702 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c30 ),
    .o({\u2_Display/lt90_c31 ,open_n5340}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_31  (
    .a(\u2_Display/n2701 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c31 ),
    .o({\u2_Display/lt90_c32 ,open_n5341}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_4  (
    .a(\u2_Display/n2728 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c4 ),
    .o({\u2_Display/lt90_c5 ,open_n5342}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_5  (
    .a(\u2_Display/n2727 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c5 ),
    .o({\u2_Display/lt90_c6 ,open_n5343}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_6  (
    .a(\u2_Display/n2726 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c6 ),
    .o({\u2_Display/lt90_c7 ,open_n5344}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_7  (
    .a(\u2_Display/n2725 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c7 ),
    .o({\u2_Display/lt90_c8 ,open_n5345}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_8  (
    .a(\u2_Display/n2724 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c8 ),
    .o({\u2_Display/lt90_c9 ,open_n5346}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_9  (
    .a(\u2_Display/n2723 ),
    .b(1'b0),
    .c(\u2_Display/lt90_c9 ),
    .o({\u2_Display/lt90_c10 ,open_n5347}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt90_cin  (
    .a(1'b0),
    .o({\u2_Display/lt90_c0 ,open_n5350}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt90_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt90_c32 ),
    .o({open_n5351,\u2_Display/n2733 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_0  (
    .a(\u2_Display/n2767 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c0 ),
    .o({\u2_Display/lt91_c1 ,open_n5352}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_1  (
    .a(\u2_Display/n2766 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c1 ),
    .o({\u2_Display/lt91_c2 ,open_n5353}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_10  (
    .a(\u2_Display/n2757 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c10 ),
    .o({\u2_Display/lt91_c11 ,open_n5354}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_11  (
    .a(\u2_Display/n2756 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c11 ),
    .o({\u2_Display/lt91_c12 ,open_n5355}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_12  (
    .a(\u2_Display/n2755 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c12 ),
    .o({\u2_Display/lt91_c13 ,open_n5356}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_13  (
    .a(\u2_Display/n2754 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c13 ),
    .o({\u2_Display/lt91_c14 ,open_n5357}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_14  (
    .a(\u2_Display/n2753 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c14 ),
    .o({\u2_Display/lt91_c15 ,open_n5358}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_15  (
    .a(\u2_Display/n2752 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c15 ),
    .o({\u2_Display/lt91_c16 ,open_n5359}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_16  (
    .a(\u2_Display/n2751 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c16 ),
    .o({\u2_Display/lt91_c17 ,open_n5360}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_17  (
    .a(\u2_Display/n2750 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c17 ),
    .o({\u2_Display/lt91_c18 ,open_n5361}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_18  (
    .a(\u2_Display/n2749 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c18 ),
    .o({\u2_Display/lt91_c19 ,open_n5362}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_19  (
    .a(\u2_Display/n2748 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c19 ),
    .o({\u2_Display/lt91_c20 ,open_n5363}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_2  (
    .a(\u2_Display/n2765 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c2 ),
    .o({\u2_Display/lt91_c3 ,open_n5364}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_20  (
    .a(\u2_Display/n2747 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c20 ),
    .o({\u2_Display/lt91_c21 ,open_n5365}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_21  (
    .a(\u2_Display/n2746 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c21 ),
    .o({\u2_Display/lt91_c22 ,open_n5366}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_22  (
    .a(\u2_Display/n2745 ),
    .b(1'b1),
    .c(\u2_Display/lt91_c22 ),
    .o({\u2_Display/lt91_c23 ,open_n5367}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_23  (
    .a(\u2_Display/n2744 ),
    .b(1'b1),
    .c(\u2_Display/lt91_c23 ),
    .o({\u2_Display/lt91_c24 ,open_n5368}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_24  (
    .a(\u2_Display/n2743 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c24 ),
    .o({\u2_Display/lt91_c25 ,open_n5369}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_25  (
    .a(\u2_Display/n2742 ),
    .b(1'b1),
    .c(\u2_Display/lt91_c25 ),
    .o({\u2_Display/lt91_c26 ,open_n5370}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_26  (
    .a(\u2_Display/n2741 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c26 ),
    .o({\u2_Display/lt91_c27 ,open_n5371}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_27  (
    .a(\u2_Display/n2740 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c27 ),
    .o({\u2_Display/lt91_c28 ,open_n5372}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_28  (
    .a(\u2_Display/n2739 ),
    .b(1'b1),
    .c(\u2_Display/lt91_c28 ),
    .o({\u2_Display/lt91_c29 ,open_n5373}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_29  (
    .a(\u2_Display/n2738 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c29 ),
    .o({\u2_Display/lt91_c30 ,open_n5374}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_3  (
    .a(\u2_Display/n2764 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c3 ),
    .o({\u2_Display/lt91_c4 ,open_n5375}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_30  (
    .a(\u2_Display/n2737 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c30 ),
    .o({\u2_Display/lt91_c31 ,open_n5376}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_31  (
    .a(\u2_Display/n2736 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c31 ),
    .o({\u2_Display/lt91_c32 ,open_n5377}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_4  (
    .a(\u2_Display/n2763 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c4 ),
    .o({\u2_Display/lt91_c5 ,open_n5378}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_5  (
    .a(\u2_Display/n2762 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c5 ),
    .o({\u2_Display/lt91_c6 ,open_n5379}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_6  (
    .a(\u2_Display/n2761 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c6 ),
    .o({\u2_Display/lt91_c7 ,open_n5380}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_7  (
    .a(\u2_Display/n2760 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c7 ),
    .o({\u2_Display/lt91_c8 ,open_n5381}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_8  (
    .a(\u2_Display/n2759 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c8 ),
    .o({\u2_Display/lt91_c9 ,open_n5382}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_9  (
    .a(\u2_Display/n2758 ),
    .b(1'b0),
    .c(\u2_Display/lt91_c9 ),
    .o({\u2_Display/lt91_c10 ,open_n5383}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt91_cin  (
    .a(1'b0),
    .o({\u2_Display/lt91_c0 ,open_n5386}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt91_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt91_c32 ),
    .o({open_n5387,\u2_Display/n2768 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_0  (
    .a(\u2_Display/n2802 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c0 ),
    .o({\u2_Display/lt92_c1 ,open_n5388}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_1  (
    .a(\u2_Display/n2801 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c1 ),
    .o({\u2_Display/lt92_c2 ,open_n5389}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_10  (
    .a(\u2_Display/n2792 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c10 ),
    .o({\u2_Display/lt92_c11 ,open_n5390}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_11  (
    .a(\u2_Display/n2791 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c11 ),
    .o({\u2_Display/lt92_c12 ,open_n5391}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_12  (
    .a(\u2_Display/n2790 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c12 ),
    .o({\u2_Display/lt92_c13 ,open_n5392}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_13  (
    .a(\u2_Display/n2789 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c13 ),
    .o({\u2_Display/lt92_c14 ,open_n5393}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_14  (
    .a(\u2_Display/n2788 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c14 ),
    .o({\u2_Display/lt92_c15 ,open_n5394}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_15  (
    .a(\u2_Display/n2787 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c15 ),
    .o({\u2_Display/lt92_c16 ,open_n5395}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_16  (
    .a(\u2_Display/n2786 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c16 ),
    .o({\u2_Display/lt92_c17 ,open_n5396}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_17  (
    .a(\u2_Display/n2785 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c17 ),
    .o({\u2_Display/lt92_c18 ,open_n5397}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_18  (
    .a(\u2_Display/n2784 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c18 ),
    .o({\u2_Display/lt92_c19 ,open_n5398}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_19  (
    .a(\u2_Display/n2783 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c19 ),
    .o({\u2_Display/lt92_c20 ,open_n5399}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_2  (
    .a(\u2_Display/n2800 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c2 ),
    .o({\u2_Display/lt92_c3 ,open_n5400}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_20  (
    .a(\u2_Display/n2782 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c20 ),
    .o({\u2_Display/lt92_c21 ,open_n5401}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_21  (
    .a(\u2_Display/n2781 ),
    .b(1'b1),
    .c(\u2_Display/lt92_c21 ),
    .o({\u2_Display/lt92_c22 ,open_n5402}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_22  (
    .a(\u2_Display/n2780 ),
    .b(1'b1),
    .c(\u2_Display/lt92_c22 ),
    .o({\u2_Display/lt92_c23 ,open_n5403}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_23  (
    .a(\u2_Display/n2779 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c23 ),
    .o({\u2_Display/lt92_c24 ,open_n5404}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_24  (
    .a(\u2_Display/n2778 ),
    .b(1'b1),
    .c(\u2_Display/lt92_c24 ),
    .o({\u2_Display/lt92_c25 ,open_n5405}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_25  (
    .a(\u2_Display/n2777 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c25 ),
    .o({\u2_Display/lt92_c26 ,open_n5406}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_26  (
    .a(\u2_Display/n2776 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c26 ),
    .o({\u2_Display/lt92_c27 ,open_n5407}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_27  (
    .a(\u2_Display/n2775 ),
    .b(1'b1),
    .c(\u2_Display/lt92_c27 ),
    .o({\u2_Display/lt92_c28 ,open_n5408}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_28  (
    .a(\u2_Display/n2774 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c28 ),
    .o({\u2_Display/lt92_c29 ,open_n5409}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_29  (
    .a(\u2_Display/n2773 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c29 ),
    .o({\u2_Display/lt92_c30 ,open_n5410}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_3  (
    .a(\u2_Display/n2799 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c3 ),
    .o({\u2_Display/lt92_c4 ,open_n5411}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_30  (
    .a(\u2_Display/n2772 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c30 ),
    .o({\u2_Display/lt92_c31 ,open_n5412}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_31  (
    .a(\u2_Display/n2771 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c31 ),
    .o({\u2_Display/lt92_c32 ,open_n5413}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_4  (
    .a(\u2_Display/n2798 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c4 ),
    .o({\u2_Display/lt92_c5 ,open_n5414}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_5  (
    .a(\u2_Display/n2797 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c5 ),
    .o({\u2_Display/lt92_c6 ,open_n5415}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_6  (
    .a(\u2_Display/n2796 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c6 ),
    .o({\u2_Display/lt92_c7 ,open_n5416}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_7  (
    .a(\u2_Display/n2795 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c7 ),
    .o({\u2_Display/lt92_c8 ,open_n5417}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_8  (
    .a(\u2_Display/n2794 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c8 ),
    .o({\u2_Display/lt92_c9 ,open_n5418}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_9  (
    .a(\u2_Display/n2793 ),
    .b(1'b0),
    .c(\u2_Display/lt92_c9 ),
    .o({\u2_Display/lt92_c10 ,open_n5419}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt92_cin  (
    .a(1'b0),
    .o({\u2_Display/lt92_c0 ,open_n5422}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt92_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt92_c32 ),
    .o({open_n5423,\u2_Display/n2803 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_0  (
    .a(\u2_Display/n2837 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c0 ),
    .o({\u2_Display/lt93_c1 ,open_n5424}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_1  (
    .a(\u2_Display/n2836 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c1 ),
    .o({\u2_Display/lt93_c2 ,open_n5425}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_10  (
    .a(\u2_Display/n2827 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c10 ),
    .o({\u2_Display/lt93_c11 ,open_n5426}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_11  (
    .a(\u2_Display/n2826 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c11 ),
    .o({\u2_Display/lt93_c12 ,open_n5427}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_12  (
    .a(\u2_Display/n2825 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c12 ),
    .o({\u2_Display/lt93_c13 ,open_n5428}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_13  (
    .a(\u2_Display/n2824 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c13 ),
    .o({\u2_Display/lt93_c14 ,open_n5429}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_14  (
    .a(\u2_Display/n2823 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c14 ),
    .o({\u2_Display/lt93_c15 ,open_n5430}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_15  (
    .a(\u2_Display/n2822 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c15 ),
    .o({\u2_Display/lt93_c16 ,open_n5431}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_16  (
    .a(\u2_Display/n2821 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c16 ),
    .o({\u2_Display/lt93_c17 ,open_n5432}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_17  (
    .a(\u2_Display/n2820 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c17 ),
    .o({\u2_Display/lt93_c18 ,open_n5433}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_18  (
    .a(\u2_Display/n2819 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c18 ),
    .o({\u2_Display/lt93_c19 ,open_n5434}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_19  (
    .a(\u2_Display/n2818 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c19 ),
    .o({\u2_Display/lt93_c20 ,open_n5435}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_2  (
    .a(\u2_Display/n2835 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c2 ),
    .o({\u2_Display/lt93_c3 ,open_n5436}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_20  (
    .a(\u2_Display/n2817 ),
    .b(1'b1),
    .c(\u2_Display/lt93_c20 ),
    .o({\u2_Display/lt93_c21 ,open_n5437}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_21  (
    .a(\u2_Display/n2816 ),
    .b(1'b1),
    .c(\u2_Display/lt93_c21 ),
    .o({\u2_Display/lt93_c22 ,open_n5438}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_22  (
    .a(\u2_Display/n2815 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c22 ),
    .o({\u2_Display/lt93_c23 ,open_n5439}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_23  (
    .a(\u2_Display/n2814 ),
    .b(1'b1),
    .c(\u2_Display/lt93_c23 ),
    .o({\u2_Display/lt93_c24 ,open_n5440}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_24  (
    .a(\u2_Display/n2813 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c24 ),
    .o({\u2_Display/lt93_c25 ,open_n5441}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_25  (
    .a(\u2_Display/n2812 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c25 ),
    .o({\u2_Display/lt93_c26 ,open_n5442}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_26  (
    .a(\u2_Display/n2811 ),
    .b(1'b1),
    .c(\u2_Display/lt93_c26 ),
    .o({\u2_Display/lt93_c27 ,open_n5443}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_27  (
    .a(\u2_Display/n2810 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c27 ),
    .o({\u2_Display/lt93_c28 ,open_n5444}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_28  (
    .a(\u2_Display/n2809 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c28 ),
    .o({\u2_Display/lt93_c29 ,open_n5445}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_29  (
    .a(\u2_Display/n2808 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c29 ),
    .o({\u2_Display/lt93_c30 ,open_n5446}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_3  (
    .a(\u2_Display/n2834 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c3 ),
    .o({\u2_Display/lt93_c4 ,open_n5447}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_30  (
    .a(\u2_Display/n2807 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c30 ),
    .o({\u2_Display/lt93_c31 ,open_n5448}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_31  (
    .a(\u2_Display/n2806 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c31 ),
    .o({\u2_Display/lt93_c32 ,open_n5449}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_4  (
    .a(\u2_Display/n2833 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c4 ),
    .o({\u2_Display/lt93_c5 ,open_n5450}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_5  (
    .a(\u2_Display/n2832 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c5 ),
    .o({\u2_Display/lt93_c6 ,open_n5451}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_6  (
    .a(\u2_Display/n2831 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c6 ),
    .o({\u2_Display/lt93_c7 ,open_n5452}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_7  (
    .a(\u2_Display/n2830 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c7 ),
    .o({\u2_Display/lt93_c8 ,open_n5453}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_8  (
    .a(\u2_Display/n2829 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c8 ),
    .o({\u2_Display/lt93_c9 ,open_n5454}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_9  (
    .a(\u2_Display/n2828 ),
    .b(1'b0),
    .c(\u2_Display/lt93_c9 ),
    .o({\u2_Display/lt93_c10 ,open_n5455}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt93_cin  (
    .a(1'b0),
    .o({\u2_Display/lt93_c0 ,open_n5458}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt93_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt93_c32 ),
    .o({open_n5459,\u2_Display/n2838 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_0  (
    .a(\u2_Display/n2872 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c0 ),
    .o({\u2_Display/lt94_c1 ,open_n5460}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_1  (
    .a(\u2_Display/n2871 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c1 ),
    .o({\u2_Display/lt94_c2 ,open_n5461}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_10  (
    .a(\u2_Display/n2862 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c10 ),
    .o({\u2_Display/lt94_c11 ,open_n5462}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_11  (
    .a(\u2_Display/n2861 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c11 ),
    .o({\u2_Display/lt94_c12 ,open_n5463}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_12  (
    .a(\u2_Display/n2860 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c12 ),
    .o({\u2_Display/lt94_c13 ,open_n5464}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_13  (
    .a(\u2_Display/n2859 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c13 ),
    .o({\u2_Display/lt94_c14 ,open_n5465}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_14  (
    .a(\u2_Display/n2858 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c14 ),
    .o({\u2_Display/lt94_c15 ,open_n5466}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_15  (
    .a(\u2_Display/n2857 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c15 ),
    .o({\u2_Display/lt94_c16 ,open_n5467}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_16  (
    .a(\u2_Display/n2856 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c16 ),
    .o({\u2_Display/lt94_c17 ,open_n5468}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_17  (
    .a(\u2_Display/n2855 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c17 ),
    .o({\u2_Display/lt94_c18 ,open_n5469}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_18  (
    .a(\u2_Display/n2854 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c18 ),
    .o({\u2_Display/lt94_c19 ,open_n5470}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_19  (
    .a(\u2_Display/n2853 ),
    .b(1'b1),
    .c(\u2_Display/lt94_c19 ),
    .o({\u2_Display/lt94_c20 ,open_n5471}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_2  (
    .a(\u2_Display/n2870 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c2 ),
    .o({\u2_Display/lt94_c3 ,open_n5472}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_20  (
    .a(\u2_Display/n2852 ),
    .b(1'b1),
    .c(\u2_Display/lt94_c20 ),
    .o({\u2_Display/lt94_c21 ,open_n5473}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_21  (
    .a(\u2_Display/n2851 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c21 ),
    .o({\u2_Display/lt94_c22 ,open_n5474}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_22  (
    .a(\u2_Display/n2850 ),
    .b(1'b1),
    .c(\u2_Display/lt94_c22 ),
    .o({\u2_Display/lt94_c23 ,open_n5475}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_23  (
    .a(\u2_Display/n2849 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c23 ),
    .o({\u2_Display/lt94_c24 ,open_n5476}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_24  (
    .a(\u2_Display/n2848 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c24 ),
    .o({\u2_Display/lt94_c25 ,open_n5477}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_25  (
    .a(\u2_Display/n2847 ),
    .b(1'b1),
    .c(\u2_Display/lt94_c25 ),
    .o({\u2_Display/lt94_c26 ,open_n5478}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_26  (
    .a(\u2_Display/n2846 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c26 ),
    .o({\u2_Display/lt94_c27 ,open_n5479}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_27  (
    .a(\u2_Display/n2845 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c27 ),
    .o({\u2_Display/lt94_c28 ,open_n5480}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_28  (
    .a(\u2_Display/n2844 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c28 ),
    .o({\u2_Display/lt94_c29 ,open_n5481}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_29  (
    .a(\u2_Display/n2843 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c29 ),
    .o({\u2_Display/lt94_c30 ,open_n5482}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_3  (
    .a(\u2_Display/n2869 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c3 ),
    .o({\u2_Display/lt94_c4 ,open_n5483}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_30  (
    .a(\u2_Display/n2842 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c30 ),
    .o({\u2_Display/lt94_c31 ,open_n5484}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_31  (
    .a(\u2_Display/n2841 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c31 ),
    .o({\u2_Display/lt94_c32 ,open_n5485}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_4  (
    .a(\u2_Display/n2868 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c4 ),
    .o({\u2_Display/lt94_c5 ,open_n5486}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_5  (
    .a(\u2_Display/n2867 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c5 ),
    .o({\u2_Display/lt94_c6 ,open_n5487}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_6  (
    .a(\u2_Display/n2866 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c6 ),
    .o({\u2_Display/lt94_c7 ,open_n5488}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_7  (
    .a(\u2_Display/n2865 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c7 ),
    .o({\u2_Display/lt94_c8 ,open_n5489}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_8  (
    .a(\u2_Display/n2864 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c8 ),
    .o({\u2_Display/lt94_c9 ,open_n5490}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_9  (
    .a(\u2_Display/n2863 ),
    .b(1'b0),
    .c(\u2_Display/lt94_c9 ),
    .o({\u2_Display/lt94_c10 ,open_n5491}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt94_cin  (
    .a(1'b0),
    .o({\u2_Display/lt94_c0 ,open_n5494}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt94_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt94_c32 ),
    .o({open_n5495,\u2_Display/n2873 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_0  (
    .a(\u2_Display/n2907 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c0 ),
    .o({\u2_Display/lt95_c1 ,open_n5496}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_1  (
    .a(\u2_Display/n2906 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c1 ),
    .o({\u2_Display/lt95_c2 ,open_n5497}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_10  (
    .a(\u2_Display/n2897 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c10 ),
    .o({\u2_Display/lt95_c11 ,open_n5498}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_11  (
    .a(\u2_Display/n2896 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c11 ),
    .o({\u2_Display/lt95_c12 ,open_n5499}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_12  (
    .a(\u2_Display/n2895 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c12 ),
    .o({\u2_Display/lt95_c13 ,open_n5500}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_13  (
    .a(\u2_Display/n2894 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c13 ),
    .o({\u2_Display/lt95_c14 ,open_n5501}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_14  (
    .a(\u2_Display/n2893 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c14 ),
    .o({\u2_Display/lt95_c15 ,open_n5502}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_15  (
    .a(\u2_Display/n2892 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c15 ),
    .o({\u2_Display/lt95_c16 ,open_n5503}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_16  (
    .a(\u2_Display/n2891 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c16 ),
    .o({\u2_Display/lt95_c17 ,open_n5504}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_17  (
    .a(\u2_Display/n2890 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c17 ),
    .o({\u2_Display/lt95_c18 ,open_n5505}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_18  (
    .a(\u2_Display/n2889 ),
    .b(1'b1),
    .c(\u2_Display/lt95_c18 ),
    .o({\u2_Display/lt95_c19 ,open_n5506}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_19  (
    .a(\u2_Display/n2888 ),
    .b(1'b1),
    .c(\u2_Display/lt95_c19 ),
    .o({\u2_Display/lt95_c20 ,open_n5507}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_2  (
    .a(\u2_Display/n2905 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c2 ),
    .o({\u2_Display/lt95_c3 ,open_n5508}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_20  (
    .a(\u2_Display/n2887 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c20 ),
    .o({\u2_Display/lt95_c21 ,open_n5509}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_21  (
    .a(\u2_Display/n2886 ),
    .b(1'b1),
    .c(\u2_Display/lt95_c21 ),
    .o({\u2_Display/lt95_c22 ,open_n5510}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_22  (
    .a(\u2_Display/n2885 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c22 ),
    .o({\u2_Display/lt95_c23 ,open_n5511}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_23  (
    .a(\u2_Display/n2884 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c23 ),
    .o({\u2_Display/lt95_c24 ,open_n5512}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_24  (
    .a(\u2_Display/n2883 ),
    .b(1'b1),
    .c(\u2_Display/lt95_c24 ),
    .o({\u2_Display/lt95_c25 ,open_n5513}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_25  (
    .a(\u2_Display/n2882 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c25 ),
    .o({\u2_Display/lt95_c26 ,open_n5514}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_26  (
    .a(\u2_Display/n2881 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c26 ),
    .o({\u2_Display/lt95_c27 ,open_n5515}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_27  (
    .a(\u2_Display/n2880 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c27 ),
    .o({\u2_Display/lt95_c28 ,open_n5516}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_28  (
    .a(\u2_Display/n2879 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c28 ),
    .o({\u2_Display/lt95_c29 ,open_n5517}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_29  (
    .a(\u2_Display/n2878 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c29 ),
    .o({\u2_Display/lt95_c30 ,open_n5518}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_3  (
    .a(\u2_Display/n2904 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c3 ),
    .o({\u2_Display/lt95_c4 ,open_n5519}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_30  (
    .a(\u2_Display/n2877 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c30 ),
    .o({\u2_Display/lt95_c31 ,open_n5520}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_31  (
    .a(\u2_Display/n2876 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c31 ),
    .o({\u2_Display/lt95_c32 ,open_n5521}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_4  (
    .a(\u2_Display/n2903 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c4 ),
    .o({\u2_Display/lt95_c5 ,open_n5522}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_5  (
    .a(\u2_Display/n2902 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c5 ),
    .o({\u2_Display/lt95_c6 ,open_n5523}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_6  (
    .a(\u2_Display/n2901 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c6 ),
    .o({\u2_Display/lt95_c7 ,open_n5524}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_7  (
    .a(\u2_Display/n2900 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c7 ),
    .o({\u2_Display/lt95_c8 ,open_n5525}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_8  (
    .a(\u2_Display/n2899 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c8 ),
    .o({\u2_Display/lt95_c9 ,open_n5526}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_9  (
    .a(\u2_Display/n2898 ),
    .b(1'b0),
    .c(\u2_Display/lt95_c9 ),
    .o({\u2_Display/lt95_c10 ,open_n5527}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt95_cin  (
    .a(1'b0),
    .o({\u2_Display/lt95_c0 ,open_n5530}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt95_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt95_c32 ),
    .o({open_n5531,\u2_Display/n2908 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_0  (
    .a(\u2_Display/n2942 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c0 ),
    .o({\u2_Display/lt96_c1 ,open_n5532}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_1  (
    .a(\u2_Display/n2941 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c1 ),
    .o({\u2_Display/lt96_c2 ,open_n5533}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_10  (
    .a(\u2_Display/n2932 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c10 ),
    .o({\u2_Display/lt96_c11 ,open_n5534}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_11  (
    .a(\u2_Display/n2931 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c11 ),
    .o({\u2_Display/lt96_c12 ,open_n5535}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_12  (
    .a(\u2_Display/n2930 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c12 ),
    .o({\u2_Display/lt96_c13 ,open_n5536}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_13  (
    .a(\u2_Display/n2929 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c13 ),
    .o({\u2_Display/lt96_c14 ,open_n5537}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_14  (
    .a(\u2_Display/n2928 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c14 ),
    .o({\u2_Display/lt96_c15 ,open_n5538}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_15  (
    .a(\u2_Display/n2927 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c15 ),
    .o({\u2_Display/lt96_c16 ,open_n5539}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_16  (
    .a(\u2_Display/n2926 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c16 ),
    .o({\u2_Display/lt96_c17 ,open_n5540}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_17  (
    .a(\u2_Display/n2925 ),
    .b(1'b1),
    .c(\u2_Display/lt96_c17 ),
    .o({\u2_Display/lt96_c18 ,open_n5541}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_18  (
    .a(\u2_Display/n2924 ),
    .b(1'b1),
    .c(\u2_Display/lt96_c18 ),
    .o({\u2_Display/lt96_c19 ,open_n5542}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_19  (
    .a(\u2_Display/n2923 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c19 ),
    .o({\u2_Display/lt96_c20 ,open_n5543}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_2  (
    .a(\u2_Display/n2940 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c2 ),
    .o({\u2_Display/lt96_c3 ,open_n5544}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_20  (
    .a(\u2_Display/n2922 ),
    .b(1'b1),
    .c(\u2_Display/lt96_c20 ),
    .o({\u2_Display/lt96_c21 ,open_n5545}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_21  (
    .a(\u2_Display/n2921 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c21 ),
    .o({\u2_Display/lt96_c22 ,open_n5546}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_22  (
    .a(\u2_Display/n2920 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c22 ),
    .o({\u2_Display/lt96_c23 ,open_n5547}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_23  (
    .a(\u2_Display/n2919 ),
    .b(1'b1),
    .c(\u2_Display/lt96_c23 ),
    .o({\u2_Display/lt96_c24 ,open_n5548}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_24  (
    .a(\u2_Display/n2918 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c24 ),
    .o({\u2_Display/lt96_c25 ,open_n5549}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_25  (
    .a(\u2_Display/n2917 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c25 ),
    .o({\u2_Display/lt96_c26 ,open_n5550}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_26  (
    .a(\u2_Display/n2916 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c26 ),
    .o({\u2_Display/lt96_c27 ,open_n5551}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_27  (
    .a(\u2_Display/n2915 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c27 ),
    .o({\u2_Display/lt96_c28 ,open_n5552}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_28  (
    .a(\u2_Display/n2914 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c28 ),
    .o({\u2_Display/lt96_c29 ,open_n5553}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_29  (
    .a(\u2_Display/n2913 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c29 ),
    .o({\u2_Display/lt96_c30 ,open_n5554}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_3  (
    .a(\u2_Display/n2939 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c3 ),
    .o({\u2_Display/lt96_c4 ,open_n5555}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_30  (
    .a(\u2_Display/n2912 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c30 ),
    .o({\u2_Display/lt96_c31 ,open_n5556}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_31  (
    .a(\u2_Display/n2911 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c31 ),
    .o({\u2_Display/lt96_c32 ,open_n5557}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_4  (
    .a(\u2_Display/n2938 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c4 ),
    .o({\u2_Display/lt96_c5 ,open_n5558}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_5  (
    .a(\u2_Display/n2937 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c5 ),
    .o({\u2_Display/lt96_c6 ,open_n5559}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_6  (
    .a(\u2_Display/n2936 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c6 ),
    .o({\u2_Display/lt96_c7 ,open_n5560}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_7  (
    .a(\u2_Display/n2935 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c7 ),
    .o({\u2_Display/lt96_c8 ,open_n5561}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_8  (
    .a(\u2_Display/n2934 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c8 ),
    .o({\u2_Display/lt96_c9 ,open_n5562}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_9  (
    .a(\u2_Display/n2933 ),
    .b(1'b0),
    .c(\u2_Display/lt96_c9 ),
    .o({\u2_Display/lt96_c10 ,open_n5563}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt96_cin  (
    .a(1'b0),
    .o({\u2_Display/lt96_c0 ,open_n5566}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt96_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt96_c32 ),
    .o({open_n5567,\u2_Display/n2943 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_0  (
    .a(\u2_Display/n2977 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c0 ),
    .o({\u2_Display/lt97_c1 ,open_n5568}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_1  (
    .a(\u2_Display/n2976 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c1 ),
    .o({\u2_Display/lt97_c2 ,open_n5569}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_10  (
    .a(\u2_Display/n2967 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c10 ),
    .o({\u2_Display/lt97_c11 ,open_n5570}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_11  (
    .a(\u2_Display/n2966 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c11 ),
    .o({\u2_Display/lt97_c12 ,open_n5571}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_12  (
    .a(\u2_Display/n2965 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c12 ),
    .o({\u2_Display/lt97_c13 ,open_n5572}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_13  (
    .a(\u2_Display/n2964 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c13 ),
    .o({\u2_Display/lt97_c14 ,open_n5573}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_14  (
    .a(\u2_Display/n2963 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c14 ),
    .o({\u2_Display/lt97_c15 ,open_n5574}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_15  (
    .a(\u2_Display/n2962 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c15 ),
    .o({\u2_Display/lt97_c16 ,open_n5575}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_16  (
    .a(\u2_Display/n2961 ),
    .b(1'b1),
    .c(\u2_Display/lt97_c16 ),
    .o({\u2_Display/lt97_c17 ,open_n5576}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_17  (
    .a(\u2_Display/n2960 ),
    .b(1'b1),
    .c(\u2_Display/lt97_c17 ),
    .o({\u2_Display/lt97_c18 ,open_n5577}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_18  (
    .a(\u2_Display/n2959 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c18 ),
    .o({\u2_Display/lt97_c19 ,open_n5578}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_19  (
    .a(\u2_Display/n2958 ),
    .b(1'b1),
    .c(\u2_Display/lt97_c19 ),
    .o({\u2_Display/lt97_c20 ,open_n5579}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_2  (
    .a(\u2_Display/n2975 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c2 ),
    .o({\u2_Display/lt97_c3 ,open_n5580}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_20  (
    .a(\u2_Display/n2957 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c20 ),
    .o({\u2_Display/lt97_c21 ,open_n5581}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_21  (
    .a(\u2_Display/n2956 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c21 ),
    .o({\u2_Display/lt97_c22 ,open_n5582}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_22  (
    .a(\u2_Display/n2955 ),
    .b(1'b1),
    .c(\u2_Display/lt97_c22 ),
    .o({\u2_Display/lt97_c23 ,open_n5583}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_23  (
    .a(\u2_Display/n2954 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c23 ),
    .o({\u2_Display/lt97_c24 ,open_n5584}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_24  (
    .a(\u2_Display/n2953 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c24 ),
    .o({\u2_Display/lt97_c25 ,open_n5585}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_25  (
    .a(\u2_Display/n2952 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c25 ),
    .o({\u2_Display/lt97_c26 ,open_n5586}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_26  (
    .a(\u2_Display/n2951 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c26 ),
    .o({\u2_Display/lt97_c27 ,open_n5587}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_27  (
    .a(\u2_Display/n2950 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c27 ),
    .o({\u2_Display/lt97_c28 ,open_n5588}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_28  (
    .a(\u2_Display/n2949 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c28 ),
    .o({\u2_Display/lt97_c29 ,open_n5589}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_29  (
    .a(\u2_Display/n2948 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c29 ),
    .o({\u2_Display/lt97_c30 ,open_n5590}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_3  (
    .a(\u2_Display/n2974 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c3 ),
    .o({\u2_Display/lt97_c4 ,open_n5591}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_30  (
    .a(\u2_Display/n2947 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c30 ),
    .o({\u2_Display/lt97_c31 ,open_n5592}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_31  (
    .a(\u2_Display/n2946 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c31 ),
    .o({\u2_Display/lt97_c32 ,open_n5593}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_4  (
    .a(\u2_Display/n2973 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c4 ),
    .o({\u2_Display/lt97_c5 ,open_n5594}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_5  (
    .a(\u2_Display/n2972 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c5 ),
    .o({\u2_Display/lt97_c6 ,open_n5595}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_6  (
    .a(\u2_Display/n2971 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c6 ),
    .o({\u2_Display/lt97_c7 ,open_n5596}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_7  (
    .a(\u2_Display/n2970 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c7 ),
    .o({\u2_Display/lt97_c8 ,open_n5597}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_8  (
    .a(\u2_Display/n2969 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c8 ),
    .o({\u2_Display/lt97_c9 ,open_n5598}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_9  (
    .a(\u2_Display/n2968 ),
    .b(1'b0),
    .c(\u2_Display/lt97_c9 ),
    .o({\u2_Display/lt97_c10 ,open_n5599}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt97_cin  (
    .a(1'b0),
    .o({\u2_Display/lt97_c0 ,open_n5602}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt97_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt97_c32 ),
    .o({open_n5603,\u2_Display/n2978 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_0  (
    .a(\u2_Display/n3012 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c0 ),
    .o({\u2_Display/lt98_c1 ,open_n5604}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_1  (
    .a(\u2_Display/n3011 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c1 ),
    .o({\u2_Display/lt98_c2 ,open_n5605}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_10  (
    .a(\u2_Display/n3002 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c10 ),
    .o({\u2_Display/lt98_c11 ,open_n5606}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_11  (
    .a(\u2_Display/n3001 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c11 ),
    .o({\u2_Display/lt98_c12 ,open_n5607}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_12  (
    .a(\u2_Display/n3000 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c12 ),
    .o({\u2_Display/lt98_c13 ,open_n5608}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_13  (
    .a(\u2_Display/n2999 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c13 ),
    .o({\u2_Display/lt98_c14 ,open_n5609}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_14  (
    .a(\u2_Display/n2998 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c14 ),
    .o({\u2_Display/lt98_c15 ,open_n5610}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_15  (
    .a(\u2_Display/n2997 ),
    .b(1'b1),
    .c(\u2_Display/lt98_c15 ),
    .o({\u2_Display/lt98_c16 ,open_n5611}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_16  (
    .a(\u2_Display/n2996 ),
    .b(1'b1),
    .c(\u2_Display/lt98_c16 ),
    .o({\u2_Display/lt98_c17 ,open_n5612}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_17  (
    .a(\u2_Display/n2995 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c17 ),
    .o({\u2_Display/lt98_c18 ,open_n5613}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_18  (
    .a(\u2_Display/n2994 ),
    .b(1'b1),
    .c(\u2_Display/lt98_c18 ),
    .o({\u2_Display/lt98_c19 ,open_n5614}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_19  (
    .a(\u2_Display/n2993 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c19 ),
    .o({\u2_Display/lt98_c20 ,open_n5615}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_2  (
    .a(\u2_Display/n3010 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c2 ),
    .o({\u2_Display/lt98_c3 ,open_n5616}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_20  (
    .a(\u2_Display/n2992 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c20 ),
    .o({\u2_Display/lt98_c21 ,open_n5617}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_21  (
    .a(\u2_Display/n2991 ),
    .b(1'b1),
    .c(\u2_Display/lt98_c21 ),
    .o({\u2_Display/lt98_c22 ,open_n5618}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_22  (
    .a(\u2_Display/n2990 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c22 ),
    .o({\u2_Display/lt98_c23 ,open_n5619}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_23  (
    .a(\u2_Display/n2989 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c23 ),
    .o({\u2_Display/lt98_c24 ,open_n5620}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_24  (
    .a(\u2_Display/n2988 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c24 ),
    .o({\u2_Display/lt98_c25 ,open_n5621}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_25  (
    .a(\u2_Display/n2987 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c25 ),
    .o({\u2_Display/lt98_c26 ,open_n5622}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_26  (
    .a(\u2_Display/n2986 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c26 ),
    .o({\u2_Display/lt98_c27 ,open_n5623}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_27  (
    .a(\u2_Display/n2985 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c27 ),
    .o({\u2_Display/lt98_c28 ,open_n5624}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_28  (
    .a(\u2_Display/n2984 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c28 ),
    .o({\u2_Display/lt98_c29 ,open_n5625}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_29  (
    .a(\u2_Display/n2983 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c29 ),
    .o({\u2_Display/lt98_c30 ,open_n5626}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_3  (
    .a(\u2_Display/n3009 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c3 ),
    .o({\u2_Display/lt98_c4 ,open_n5627}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_30  (
    .a(\u2_Display/n2982 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c30 ),
    .o({\u2_Display/lt98_c31 ,open_n5628}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_31  (
    .a(\u2_Display/n2981 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c31 ),
    .o({\u2_Display/lt98_c32 ,open_n5629}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_4  (
    .a(\u2_Display/n3008 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c4 ),
    .o({\u2_Display/lt98_c5 ,open_n5630}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_5  (
    .a(\u2_Display/n3007 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c5 ),
    .o({\u2_Display/lt98_c6 ,open_n5631}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_6  (
    .a(\u2_Display/n3006 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c6 ),
    .o({\u2_Display/lt98_c7 ,open_n5632}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_7  (
    .a(\u2_Display/n3005 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c7 ),
    .o({\u2_Display/lt98_c8 ,open_n5633}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_8  (
    .a(\u2_Display/n3004 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c8 ),
    .o({\u2_Display/lt98_c9 ,open_n5634}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_9  (
    .a(\u2_Display/n3003 ),
    .b(1'b0),
    .c(\u2_Display/lt98_c9 ),
    .o({\u2_Display/lt98_c10 ,open_n5635}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt98_cin  (
    .a(1'b0),
    .o({\u2_Display/lt98_c0 ,open_n5638}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt98_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt98_c32 ),
    .o({open_n5639,\u2_Display/n3013 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_0  (
    .a(\u2_Display/n3047 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c0 ),
    .o({\u2_Display/lt99_c1 ,open_n5640}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_1  (
    .a(\u2_Display/n3046 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c1 ),
    .o({\u2_Display/lt99_c2 ,open_n5641}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_10  (
    .a(\u2_Display/n3037 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c10 ),
    .o({\u2_Display/lt99_c11 ,open_n5642}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_11  (
    .a(\u2_Display/n3036 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c11 ),
    .o({\u2_Display/lt99_c12 ,open_n5643}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_12  (
    .a(\u2_Display/n3035 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c12 ),
    .o({\u2_Display/lt99_c13 ,open_n5644}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_13  (
    .a(\u2_Display/n3034 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c13 ),
    .o({\u2_Display/lt99_c14 ,open_n5645}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_14  (
    .a(\u2_Display/n3033 ),
    .b(1'b1),
    .c(\u2_Display/lt99_c14 ),
    .o({\u2_Display/lt99_c15 ,open_n5646}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_15  (
    .a(\u2_Display/n3032 ),
    .b(1'b1),
    .c(\u2_Display/lt99_c15 ),
    .o({\u2_Display/lt99_c16 ,open_n5647}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_16  (
    .a(\u2_Display/n3031 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c16 ),
    .o({\u2_Display/lt99_c17 ,open_n5648}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_17  (
    .a(\u2_Display/n3030 ),
    .b(1'b1),
    .c(\u2_Display/lt99_c17 ),
    .o({\u2_Display/lt99_c18 ,open_n5649}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_18  (
    .a(\u2_Display/n3029 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c18 ),
    .o({\u2_Display/lt99_c19 ,open_n5650}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_19  (
    .a(\u2_Display/n3028 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c19 ),
    .o({\u2_Display/lt99_c20 ,open_n5651}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_2  (
    .a(\u2_Display/n3045 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c2 ),
    .o({\u2_Display/lt99_c3 ,open_n5652}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_20  (
    .a(\u2_Display/n3027 ),
    .b(1'b1),
    .c(\u2_Display/lt99_c20 ),
    .o({\u2_Display/lt99_c21 ,open_n5653}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_21  (
    .a(\u2_Display/n3026 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c21 ),
    .o({\u2_Display/lt99_c22 ,open_n5654}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_22  (
    .a(\u2_Display/n3025 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c22 ),
    .o({\u2_Display/lt99_c23 ,open_n5655}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_23  (
    .a(\u2_Display/n3024 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c23 ),
    .o({\u2_Display/lt99_c24 ,open_n5656}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_24  (
    .a(\u2_Display/n3023 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c24 ),
    .o({\u2_Display/lt99_c25 ,open_n5657}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_25  (
    .a(\u2_Display/n3022 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c25 ),
    .o({\u2_Display/lt99_c26 ,open_n5658}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_26  (
    .a(\u2_Display/n3021 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c26 ),
    .o({\u2_Display/lt99_c27 ,open_n5659}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_27  (
    .a(\u2_Display/n3020 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c27 ),
    .o({\u2_Display/lt99_c28 ,open_n5660}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_28  (
    .a(\u2_Display/n3019 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c28 ),
    .o({\u2_Display/lt99_c29 ,open_n5661}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_29  (
    .a(\u2_Display/n3018 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c29 ),
    .o({\u2_Display/lt99_c30 ,open_n5662}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_3  (
    .a(\u2_Display/n3044 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c3 ),
    .o({\u2_Display/lt99_c4 ,open_n5663}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_30  (
    .a(\u2_Display/n3017 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c30 ),
    .o({\u2_Display/lt99_c31 ,open_n5664}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_31  (
    .a(\u2_Display/n3016 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c31 ),
    .o({\u2_Display/lt99_c32 ,open_n5665}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_4  (
    .a(\u2_Display/n3043 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c4 ),
    .o({\u2_Display/lt99_c5 ,open_n5666}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_5  (
    .a(\u2_Display/n3042 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c5 ),
    .o({\u2_Display/lt99_c6 ,open_n5667}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_6  (
    .a(\u2_Display/n3041 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c6 ),
    .o({\u2_Display/lt99_c7 ,open_n5668}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_7  (
    .a(\u2_Display/n3040 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c7 ),
    .o({\u2_Display/lt99_c8 ,open_n5669}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_8  (
    .a(\u2_Display/n3039 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c8 ),
    .o({\u2_Display/lt99_c9 ,open_n5670}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_9  (
    .a(\u2_Display/n3038 ),
    .b(1'b0),
    .c(\u2_Display/lt99_c9 ),
    .o({\u2_Display/lt99_c10 ,open_n5671}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt99_cin  (
    .a(1'b0),
    .o({\u2_Display/lt99_c0 ,open_n5674}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt99_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt99_c32 ),
    .o({open_n5675,\u2_Display/n3048 }));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_0  (
    .a(\u2_Display/n137 [0]),
    .b(lcd_xpos[0]),
    .c(\u2_Display/lt9_2_c0 ),
    .o({\u2_Display/lt9_2_c1 ,open_n5676}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_1  (
    .a(\u2_Display/n137 [1]),
    .b(lcd_xpos[1]),
    .c(\u2_Display/lt9_2_c1 ),
    .o({\u2_Display/lt9_2_c2 ,open_n5677}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_10  (
    .a(\u2_Display/n137 [31]),
    .b(lcd_xpos[10]),
    .c(\u2_Display/lt9_2_c10 ),
    .o({\u2_Display/lt9_2_c11 ,open_n5678}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_11  (
    .a(\u2_Display/n137 [31]),
    .b(lcd_xpos[11]),
    .c(\u2_Display/lt9_2_c11 ),
    .o({\u2_Display/lt9_2_c12 ,open_n5679}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_12  (
    .a(\u2_Display/n137 [31]),
    .b(1'b0),
    .c(\u2_Display/lt9_2_c12 ),
    .o({\u2_Display/lt9_2_c13 ,open_n5680}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_2  (
    .a(\u2_Display/n137 [2]),
    .b(lcd_xpos[2]),
    .c(\u2_Display/lt9_2_c2 ),
    .o({\u2_Display/lt9_2_c3 ,open_n5681}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_3  (
    .a(\u2_Display/n137 [3]),
    .b(lcd_xpos[3]),
    .c(\u2_Display/lt9_2_c3 ),
    .o({\u2_Display/lt9_2_c4 ,open_n5682}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_4  (
    .a(\u2_Display/n137 [4]),
    .b(lcd_xpos[4]),
    .c(\u2_Display/lt9_2_c4 ),
    .o({\u2_Display/lt9_2_c5 ,open_n5683}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_5  (
    .a(\u2_Display/n137 [5]),
    .b(lcd_xpos[5]),
    .c(\u2_Display/lt9_2_c5 ),
    .o({\u2_Display/lt9_2_c6 ,open_n5684}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_6  (
    .a(\u2_Display/n137 [6]),
    .b(lcd_xpos[6]),
    .c(\u2_Display/lt9_2_c6 ),
    .o({\u2_Display/lt9_2_c7 ,open_n5685}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_7  (
    .a(\u2_Display/n137 [7]),
    .b(lcd_xpos[7]),
    .c(\u2_Display/lt9_2_c7 ),
    .o({\u2_Display/lt9_2_c8 ,open_n5686}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_8  (
    .a(\u2_Display/n137 [8]),
    .b(lcd_xpos[8]),
    .c(\u2_Display/lt9_2_c8 ),
    .o({\u2_Display/lt9_2_c9 ,open_n5687}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_9  (
    .a(\u2_Display/n137 [9]),
    .b(lcd_xpos[9]),
    .c(\u2_Display/lt9_2_c9 ),
    .o({\u2_Display/lt9_2_c10 ,open_n5688}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u2_Display/lt9_2_cin  (
    .a(1'b0),
    .o({\u2_Display/lt9_2_c0 ,open_n5691}));
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u2_Display/lt9_2_cout  (
    .a(1'b0),
    .b(1'b1),
    .c(\u2_Display/lt9_2_c13 ),
    .o({open_n5692,\u2_Display/n138 }));
  reg_sr_as_w1 \u2_Display/reg0_b0  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [0]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [0]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b1  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [1]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [1]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b10  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [10]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [10]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b11  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [11]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [11]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b12  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [12]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [12]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b13  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [13]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [13]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b14  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [14]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [14]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b15  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [15]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [15]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b16  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [16]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [16]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b17  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [17]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [17]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b18  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [18]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [18]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b19  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [19]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [19]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b2  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [2]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [2]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b20  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [20]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [20]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b21  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [21]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [21]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b22  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [22]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [22]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b23  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [23]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [23]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b24  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [24]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [24]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b25  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [25]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [25]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b26  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [26]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [26]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b27  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [27]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [27]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b28  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [28]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [28]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b29  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [29]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [29]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b3  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [3]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [3]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b30  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [30]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [30]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b4  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [4]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [4]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b5  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [5]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [5]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b6  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [6]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [6]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b7  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [7]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [7]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b8  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [8]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [8]));  // source/rtl/Display.v(61)
  reg_sr_as_w1 \u2_Display/reg0_b9  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [9]),
    .en(1'b1),
    .reset(\u2_Display/n35 ),
    .set(1'b0),
    .q(\u2_Display/n [9]));  // source/rtl/Display.v(61)
  reg_ar_as_w1 \u2_Display/reg1_b0  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n240 [0]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(lcd_data[23]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b0  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [0]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [0]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b1  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [1]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [1]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b10  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [10]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [10]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b11  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [11]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [11]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b12  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [12]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [12]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b13  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [13]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [13]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b14  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [14]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [14]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b15  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [15]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [15]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b16  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [16]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [16]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b17  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [17]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [17]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b18  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [18]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [18]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b19  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [19]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [19]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b2  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [2]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [2]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b20  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [20]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [20]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b21  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [21]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [21]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b22  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [22]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [22]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b23  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [23]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [23]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b24  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [24]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [24]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b25  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [25]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [25]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b26  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [26]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [26]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b27  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [27]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [27]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b28  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [28]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [28]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b29  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [29]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [29]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b3  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [3]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [3]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b30  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [30]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [30]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b31  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [31]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [31]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b4  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [4]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [4]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b5  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [5]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [5]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b6  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [6]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [6]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b7  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [7]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [7]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b8  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [8]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [8]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg2_b9  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [9]),
    .en(\u2_Display/mux21_b0_sel_is_0_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/counta [9]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b0  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [0]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [0]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b1  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [1]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [1]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b10  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [10]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [10]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b2  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [2]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [2]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b3  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [3]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [3]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b4  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [4]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [4]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b5  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [5]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [5]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b6  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [6]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [6]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b7  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [7]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [7]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b8  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [8]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [8]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg3_b9  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [9]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/i [9]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b0  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [0]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [0]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b1  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [1]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [1]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b2  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [2]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [2]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b3  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [3]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [3]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b4  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [4]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [4]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b5  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [5]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [5]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b6  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [6]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [6]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b7  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [7]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [7]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b8  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [8]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [8]));  // source/rtl/Display.v(252)
  reg_ar_as_w1 \u2_Display/reg4_b9  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [9]),
    .en(rst_n_pad),
    .reset(1'b0),
    .set(1'b0),
    .q(\u2_Display/j [9]));  // source/rtl/Display.v(252)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub0_2/u0  (
    .a(1'b0),
    .b(\u2_Display/i [0]),
    .c(\u2_Display/sub0_2/c0 ),
    .o({\u2_Display/sub0_2/c1 ,\u2_Display/n96 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub0_2/u1  (
    .a(1'b0),
    .b(\u2_Display/i [1]),
    .c(\u2_Display/sub0_2/c1 ),
    .o({\u2_Display/sub0_2/c2 ,\u2_Display/n96 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub0_2/u10  (
    .a(1'b0),
    .b(\u2_Display/i [10]),
    .c(\u2_Display/sub0_2/c10 ),
    .o({\u2_Display/sub0_2/c11 ,\u2_Display/n96 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub0_2/u2  (
    .a(1'b0),
    .b(\u2_Display/i [2]),
    .c(\u2_Display/sub0_2/c2 ),
    .o({\u2_Display/sub0_2/c3 ,\u2_Display/n96 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub0_2/u3  (
    .a(1'b0),
    .b(\u2_Display/i [3]),
    .c(\u2_Display/sub0_2/c3 ),
    .o({\u2_Display/sub0_2/c4 ,\u2_Display/n96 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub0_2/u4  (
    .a(1'b0),
    .b(\u2_Display/i [4]),
    .c(\u2_Display/sub0_2/c4 ),
    .o({\u2_Display/sub0_2/c5 ,\u2_Display/n96 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub0_2/u5  (
    .a(1'b0),
    .b(\u2_Display/i [5]),
    .c(\u2_Display/sub0_2/c5 ),
    .o({\u2_Display/sub0_2/c6 ,\u2_Display/n96 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub0_2/u6  (
    .a(1'b0),
    .b(\u2_Display/i [6]),
    .c(\u2_Display/sub0_2/c6 ),
    .o({\u2_Display/sub0_2/c7 ,\u2_Display/n96 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub0_2/u7  (
    .a(1'b1),
    .b(\u2_Display/i [7]),
    .c(\u2_Display/sub0_2/c7 ),
    .o({\u2_Display/sub0_2/c8 ,\u2_Display/n96 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub0_2/u8  (
    .a(1'b0),
    .b(\u2_Display/i [8]),
    .c(\u2_Display/sub0_2/c8 ),
    .o({\u2_Display/sub0_2/c9 ,\u2_Display/n96 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub0_2/u9  (
    .a(1'b1),
    .b(\u2_Display/i [9]),
    .c(\u2_Display/sub0_2/c9 ),
    .o({\u2_Display/sub0_2/c10 ,\u2_Display/n96 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u2_Display/sub0_2/ucin  (
    .a(1'b0),
    .o({\u2_Display/sub0_2/c0 ,open_n5695}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub0_2/ucout  (
    .c(\u2_Display/sub0_2/c11 ),
    .o({open_n5698,\u2_Display/n96 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub1_2/u0  (
    .a(1'b0),
    .b(\u2_Display/j [0]),
    .c(\u2_Display/sub1_2/c0 ),
    .o({\u2_Display/sub1_2/c1 ,\u2_Display/n102 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub1_2/u1  (
    .a(1'b0),
    .b(\u2_Display/j [1]),
    .c(\u2_Display/sub1_2/c1 ),
    .o({\u2_Display/sub1_2/c2 ,\u2_Display/n102 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub1_2/u2  (
    .a(1'b0),
    .b(\u2_Display/j [2]),
    .c(\u2_Display/sub1_2/c2 ),
    .o({\u2_Display/sub1_2/c3 ,\u2_Display/n102 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub1_2/u3  (
    .a(1'b0),
    .b(\u2_Display/j [3]),
    .c(\u2_Display/sub1_2/c3 ),
    .o({\u2_Display/sub1_2/c4 ,\u2_Display/n102 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub1_2/u4  (
    .a(1'b0),
    .b(\u2_Display/j [4]),
    .c(\u2_Display/sub1_2/c4 ),
    .o({\u2_Display/sub1_2/c5 ,\u2_Display/n102 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub1_2/u5  (
    .a(1'b0),
    .b(\u2_Display/j [5]),
    .c(\u2_Display/sub1_2/c5 ),
    .o({\u2_Display/sub1_2/c6 ,\u2_Display/n102 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub1_2/u6  (
    .a(1'b0),
    .b(\u2_Display/j [6]),
    .c(\u2_Display/sub1_2/c6 ),
    .o({\u2_Display/sub1_2/c7 ,\u2_Display/n102 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub1_2/u7  (
    .a(1'b0),
    .b(\u2_Display/j [7]),
    .c(\u2_Display/sub1_2/c7 ),
    .o({\u2_Display/sub1_2/c8 ,\u2_Display/n102 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub1_2/u8  (
    .a(1'b0),
    .b(\u2_Display/j [8]),
    .c(\u2_Display/sub1_2/c8 ),
    .o({\u2_Display/sub1_2/c9 ,\u2_Display/n102 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub1_2/u9  (
    .a(1'b1),
    .b(\u2_Display/j [9]),
    .c(\u2_Display/sub1_2/c9 ),
    .o({\u2_Display/sub1_2/c10 ,\u2_Display/n102 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u2_Display/sub1_2/ucin  (
    .a(1'b0),
    .o({\u2_Display/sub1_2/c0 ,open_n5701}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub1_2/ucout  (
    .c(\u2_Display/sub1_2/c10 ),
    .o({open_n5704,\u2_Display/n102 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub2_2/u0  (
    .a(1'b0),
    .b(\u2_Display/j [0]),
    .c(\u2_Display/sub2_2/c0 ),
    .o({\u2_Display/sub2_2/c1 ,\u2_Display/n137 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub2_2/u1  (
    .a(1'b0),
    .b(\u2_Display/j [1]),
    .c(\u2_Display/sub2_2/c1 ),
    .o({\u2_Display/sub2_2/c2 ,\u2_Display/n137 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub2_2/u2  (
    .a(1'b0),
    .b(\u2_Display/j [2]),
    .c(\u2_Display/sub2_2/c2 ),
    .o({\u2_Display/sub2_2/c3 ,\u2_Display/n137 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub2_2/u3  (
    .a(1'b0),
    .b(\u2_Display/j [3]),
    .c(\u2_Display/sub2_2/c3 ),
    .o({\u2_Display/sub2_2/c4 ,\u2_Display/n137 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub2_2/u4  (
    .a(1'b0),
    .b(\u2_Display/j [4]),
    .c(\u2_Display/sub2_2/c4 ),
    .o({\u2_Display/sub2_2/c5 ,\u2_Display/n137 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub2_2/u5  (
    .a(1'b0),
    .b(\u2_Display/j [5]),
    .c(\u2_Display/sub2_2/c5 ),
    .o({\u2_Display/sub2_2/c6 ,\u2_Display/n137 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub2_2/u6  (
    .a(1'b0),
    .b(\u2_Display/j [6]),
    .c(\u2_Display/sub2_2/c6 ),
    .o({\u2_Display/sub2_2/c7 ,\u2_Display/n137 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub2_2/u7  (
    .a(1'b1),
    .b(\u2_Display/j [7]),
    .c(\u2_Display/sub2_2/c7 ),
    .o({\u2_Display/sub2_2/c8 ,\u2_Display/n137 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub2_2/u8  (
    .a(1'b0),
    .b(\u2_Display/j [8]),
    .c(\u2_Display/sub2_2/c8 ),
    .o({\u2_Display/sub2_2/c9 ,\u2_Display/n137 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub2_2/u9  (
    .a(1'b1),
    .b(\u2_Display/j [9]),
    .c(\u2_Display/sub2_2/c9 ),
    .o({\u2_Display/sub2_2/c10 ,\u2_Display/n137 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u2_Display/sub2_2/ucin  (
    .a(1'b0),
    .o({\u2_Display/sub2_2/c0 ,open_n5707}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub2_2/ucout  (
    .c(\u2_Display/sub2_2/c10 ),
    .o({open_n5710,\u2_Display/n137 [31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub3_2/u0  (
    .a(1'b0),
    .b(\u2_Display/i [0]),
    .c(\u2_Display/sub3_2/c0 ),
    .o({\u2_Display/sub3_2/c1 ,\u2_Display/n143 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub3_2/u1  (
    .a(1'b0),
    .b(\u2_Display/i [1]),
    .c(\u2_Display/sub3_2/c1 ),
    .o({\u2_Display/sub3_2/c2 ,\u2_Display/n143 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub3_2/u10  (
    .a(1'b0),
    .b(\u2_Display/i [10]),
    .c(\u2_Display/sub3_2/c10 ),
    .o({\u2_Display/sub3_2/c11 ,\u2_Display/n143 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub3_2/u2  (
    .a(1'b0),
    .b(\u2_Display/i [2]),
    .c(\u2_Display/sub3_2/c2 ),
    .o({\u2_Display/sub3_2/c3 ,\u2_Display/n143 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub3_2/u3  (
    .a(1'b0),
    .b(\u2_Display/i [3]),
    .c(\u2_Display/sub3_2/c3 ),
    .o({\u2_Display/sub3_2/c4 ,\u2_Display/n143 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub3_2/u4  (
    .a(1'b0),
    .b(\u2_Display/i [4]),
    .c(\u2_Display/sub3_2/c4 ),
    .o({\u2_Display/sub3_2/c5 ,\u2_Display/n143 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub3_2/u5  (
    .a(1'b0),
    .b(\u2_Display/i [5]),
    .c(\u2_Display/sub3_2/c5 ),
    .o({\u2_Display/sub3_2/c6 ,\u2_Display/n143 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub3_2/u6  (
    .a(1'b0),
    .b(\u2_Display/i [6]),
    .c(\u2_Display/sub3_2/c6 ),
    .o({\u2_Display/sub3_2/c7 ,\u2_Display/n143 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub3_2/u7  (
    .a(1'b0),
    .b(\u2_Display/i [7]),
    .c(\u2_Display/sub3_2/c7 ),
    .o({\u2_Display/sub3_2/c8 ,\u2_Display/n143 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub3_2/u8  (
    .a(1'b0),
    .b(\u2_Display/i [8]),
    .c(\u2_Display/sub3_2/c8 ),
    .o({\u2_Display/sub3_2/c9 ,\u2_Display/n143 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub3_2/u9  (
    .a(1'b1),
    .b(\u2_Display/i [9]),
    .c(\u2_Display/sub3_2/c9 ),
    .o({\u2_Display/sub3_2/c10 ,\u2_Display/n143 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u2_Display/sub3_2/ucin  (
    .a(1'b0),
    .o({\u2_Display/sub3_2/c0 ,open_n5713}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u2_Display/sub3_2/ucout  (
    .c(\u2_Display/sub3_2/c11 ),
    .o({open_n5716,\u2_Display/n143 [31]}));

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  // synthesis translate_off
  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end
  // synthesis translate_on

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

