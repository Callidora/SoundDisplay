// Verilog netlist created by TD v5.0.19080
// Sun May 31 12:05:43 2020

`timescale 1ns / 1ps
module VGA_Demo  // source/rtl/VGA_Demo.v(2)
  (
  clk_24m,
  on_off,
  rst_n,
  vga_b,
  vga_clk,
  vga_de,
  vga_g,
  vga_hs,
  vga_r,
  vga_vs
  );

  input clk_24m;  // source/rtl/VGA_Demo.v(4)
  input [7:0] on_off;  // source/rtl/VGA_Demo.v(6)
  input rst_n;  // source/rtl/VGA_Demo.v(5)
  output [7:0] vga_b;  // source/rtl/VGA_Demo.v(17)
  output vga_clk;  // source/rtl/VGA_Demo.v(9)
  output vga_de;  // source/rtl/VGA_Demo.v(13)
  output [7:0] vga_g;  // source/rtl/VGA_Demo.v(16)
  output vga_hs;  // source/rtl/VGA_Demo.v(10)
  output [7:0] vga_r;  // source/rtl/VGA_Demo.v(15)
  output vga_vs;  // source/rtl/VGA_Demo.v(11)

  wire [23:0] lcd_data;  // source/rtl/VGA_Demo.v(23)
  wire [11:0] lcd_xpos;  // source/rtl/VGA_Demo.v(21)
  wire [11:0] lcd_ypos;  // source/rtl/VGA_Demo.v(22)
  wire [7:0] on_off_pad;  // source/rtl/VGA_Demo.v(6)
  wire [11:0] \u1_Driver/hcnt ;  // source/rtl/Driver.v(44)
  wire [11:0] \u1_Driver/n2 ;
  wire [12:0] \u1_Driver/n20 ;
  wire [12:0] \u1_Driver/n21 ;
  wire [11:0] \u1_Driver/n7 ;
  wire [11:0] \u1_Driver/vcnt ;  // source/rtl/Driver.v(45)
  wire [31:0] \u2_Display/counta ;  // source/rtl/Display.v(39)
  wire [31:0] \u2_Display/i ;  // source/rtl/Display.v(41)
  wire [31:0] \u2_Display/j ;  // source/rtl/Display.v(42)
  wire [30:0] \u2_Display/n ;  // source/rtl/Display.v(48)
  wire [31:0] \u2_Display/n1014 ;
  wire [31:0] \u2_Display/n102 ;
  wire [31:0] \u2_Display/n1049 ;
  wire [31:0] \u2_Display/n1084 ;
  wire [31:0] \u2_Display/n1119 ;
  wire [31:0] \u2_Display/n1154 ;
  wire [31:0] \u2_Display/n1189 ;
  wire [24:0] \u2_Display/n135 ;
  wire [31:0] \u2_Display/n137 ;
  wire [22:0] \u2_Display/n140 ;
  wire [31:0] \u2_Display/n143 ;
  wire [31:0] \u2_Display/n1542 ;
  wire [31:0] \u2_Display/n1577 ;
  wire [31:0] \u2_Display/n1612 ;
  wire [31:0] \u2_Display/n1647 ;
  wire [31:0] \u2_Display/n1682 ;
  wire [31:0] \u2_Display/n1717 ;
  wire [31:0] \u2_Display/n1752 ;
  wire [31:0] \u2_Display/n1787 ;
  wire [31:0] \u2_Display/n1822 ;
  wire [31:0] \u2_Display/n1857 ;
  wire [31:0] \u2_Display/n1892 ;
  wire [31:0] \u2_Display/n1927 ;
  wire [31:0] \u2_Display/n1962 ;
  wire [31:0] \u2_Display/n1997 ;
  wire [31:0] \u2_Display/n2032 ;
  wire [31:0] \u2_Display/n2067 ;
  wire [31:0] \u2_Display/n2102 ;
  wire [31:0] \u2_Display/n2137 ;
  wire [31:0] \u2_Display/n2172 ;
  wire [31:0] \u2_Display/n2207 ;
  wire [31:0] \u2_Display/n2242 ;
  wire [31:0] \u2_Display/n2277 ;
  wire [31:0] \u2_Display/n2312 ;
  wire [23:0] \u2_Display/n236 ;
  wire [31:0] \u2_Display/n2665 ;
  wire [31:0] \u2_Display/n2700 ;
  wire [31:0] \u2_Display/n2735 ;
  wire [31:0] \u2_Display/n2770 ;
  wire [31:0] \u2_Display/n2805 ;
  wire [31:0] \u2_Display/n2840 ;
  wire [31:0] \u2_Display/n2875 ;
  wire [31:0] \u2_Display/n2910 ;
  wire [31:0] \u2_Display/n2945 ;
  wire [31:0] \u2_Display/n2980 ;
  wire [31:0] \u2_Display/n3015 ;
  wire [31:0] \u2_Display/n3050 ;
  wire [31:0] \u2_Display/n3085 ;
  wire [31:0] \u2_Display/n3120 ;
  wire [31:0] \u2_Display/n3155 ;
  wire [31:0] \u2_Display/n3190 ;
  wire [31:0] \u2_Display/n3225 ;
  wire [31:0] \u2_Display/n3260 ;
  wire [31:0] \u2_Display/n3295 ;
  wire [31:0] \u2_Display/n3330 ;
  wire [31:0] \u2_Display/n3365 ;
  wire [31:0] \u2_Display/n3400 ;
  wire [31:0] \u2_Display/n3435 ;
  wire [30:0] \u2_Display/n37 ;
  wire [31:0] \u2_Display/n3788 ;
  wire [31:0] \u2_Display/n3823 ;
  wire [31:0] \u2_Display/n3858 ;
  wire [31:0] \u2_Display/n3893 ;
  wire [31:0] \u2_Display/n3928 ;
  wire [31:0] \u2_Display/n3963 ;
  wire [31:0] \u2_Display/n3998 ;
  wire [31:0] \u2_Display/n4033 ;
  wire [31:0] \u2_Display/n4068 ;
  wire [31:0] \u2_Display/n41 ;
  wire [31:0] \u2_Display/n4103 ;
  wire [31:0] \u2_Display/n4138 ;
  wire [31:0] \u2_Display/n4173 ;
  wire [31:0] \u2_Display/n419 ;
  wire [31:0] \u2_Display/n4208 ;
  wire [31:0] \u2_Display/n4243 ;
  wire [31:0] \u2_Display/n4278 ;
  wire [23:0] \u2_Display/n43 ;
  wire [31:0] \u2_Display/n4313 ;
  wire [31:0] \u2_Display/n4348 ;
  wire [31:0] \u2_Display/n4383 ;
  wire [31:0] \u2_Display/n4418 ;
  wire [31:0] \u2_Display/n4453 ;
  wire [31:0] \u2_Display/n4488 ;
  wire [31:0] \u2_Display/n4523 ;
  wire [31:0] \u2_Display/n454 ;
  wire [31:0] \u2_Display/n4558 ;
  wire [31:0] \u2_Display/n489 ;
  wire [31:0] \u2_Display/n4911 ;
  wire [31:0] \u2_Display/n4946 ;
  wire [31:0] \u2_Display/n4981 ;
  wire [31:0] \u2_Display/n5016 ;
  wire [31:0] \u2_Display/n5051 ;
  wire [31:0] \u2_Display/n5086 ;
  wire [31:0] \u2_Display/n5121 ;
  wire [31:0] \u2_Display/n5156 ;
  wire [31:0] \u2_Display/n5191 ;
  wire [31:0] \u2_Display/n5226 ;
  wire [31:0] \u2_Display/n524 ;
  wire [31:0] \u2_Display/n5261 ;
  wire [31:0] \u2_Display/n5296 ;
  wire [31:0] \u2_Display/n5331 ;
  wire [31:0] \u2_Display/n5366 ;
  wire [31:0] \u2_Display/n5401 ;
  wire [31:0] \u2_Display/n5436 ;
  wire [31:0] \u2_Display/n5471 ;
  wire [31:0] \u2_Display/n5506 ;
  wire [31:0] \u2_Display/n5541 ;
  wire [31:0] \u2_Display/n5576 ;
  wire [31:0] \u2_Display/n559 ;
  wire [31:0] \u2_Display/n5611 ;
  wire [31:0] \u2_Display/n5646 ;
  wire [31:0] \u2_Display/n5681 ;
  wire [31:0] \u2_Display/n594 ;
  wire [31:0] \u2_Display/n629 ;
  wire [31:0] \u2_Display/n664 ;
  wire [31:0] \u2_Display/n699 ;
  wire [31:0] \u2_Display/n734 ;
  wire [31:0] \u2_Display/n769 ;
  wire [31:0] \u2_Display/n804 ;
  wire [31:0] \u2_Display/n839 ;
  wire [31:0] \u2_Display/n874 ;
  wire [31:0] \u2_Display/n909 ;
  wire [24:0] \u2_Display/n94 ;
  wire [31:0] \u2_Display/n944 ;
  wire [31:0] \u2_Display/n96 ;
  wire [31:0] \u2_Display/n979 ;
  wire [22:0] \u2_Display/n99 ;
  wire [7:0] vga_b_pad;  // source/rtl/VGA_Demo.v(17)
  wire _al_u1168_o;
  wire _al_u1170_o;
  wire _al_u1171_o;
  wire _al_u1345_o;
  wire _al_u1346_o;
  wire _al_u1347_o;
  wire _al_u1348_o;
  wire _al_u1349_o;
  wire _al_u1350_o;
  wire _al_u1351_o;
  wire _al_u1352_o;
  wire _al_u1353_o;
  wire _al_u3916_o;
  wire _al_u3917_o;
  wire _al_u3918_o;
  wire _al_u3920_o;
  wire _al_u3921_o;
  wire _al_u3922_o;
  wire _al_u3924_o;
  wire _al_u3925_o;
  wire _al_u3926_o;
  wire _al_u3928_o;
  wire _al_u3929_o;
  wire _al_u3930_o;
  wire _al_u3932_o;
  wire _al_u3933_o;
  wire _al_u3934_o;
  wire _al_u3936_o;
  wire _al_u3937_o;
  wire _al_u3938_o;
  wire _al_u3940_o;
  wire _al_u3941_o;
  wire _al_u3942_o;
  wire _al_u3944_o;
  wire _al_u3945_o;
  wire _al_u3946_o;
  wire _al_u3948_o;
  wire _al_u3949_o;
  wire _al_u3950_o;
  wire _al_u3952_o;
  wire _al_u3953_o;
  wire _al_u3954_o;
  wire _al_u3956_o;
  wire _al_u3957_o;
  wire _al_u3958_o;
  wire _al_u3960_o;
  wire _al_u3961_o;
  wire _al_u3962_o;
  wire _al_u3963_o;
  wire _al_u3965_o;
  wire _al_u3966_o;
  wire _al_u3967_o;
  wire _al_u3969_o;
  wire _al_u3970_o;
  wire _al_u3971_o;
  wire _al_u3972_o;
  wire _al_u3974_o;
  wire _al_u3975_o;
  wire _al_u3976_o;
  wire _al_u3978_o;
  wire _al_u3979_o;
  wire _al_u3980_o;
  wire _al_u3981_o;
  wire _al_u3983_o;
  wire _al_u3984_o;
  wire _al_u3985_o;
  wire _al_u3987_o;
  wire _al_u3988_o;
  wire _al_u3989_o;
  wire _al_u3991_o;
  wire _al_u3992_o;
  wire _al_u3993_o;
  wire _al_u3995_o;
  wire _al_u3996_o;
  wire _al_u3997_o;
  wire _al_u997_o;
  wire _al_u998_o;
  wire clk_24m_pad;  // source/rtl/VGA_Demo.v(4)
  wire clk_vga;  // source/rtl/VGA_Demo.v(20)
  wire rst_n_pad;  // source/rtl/VGA_Demo.v(5)
  wire \u0_PLL/n0 ;
  wire \u0_PLL/uut/clk0_buf ;  // al_ip/PLL.v(32)
  wire \u1_Driver/add0/c11 ;
  wire \u1_Driver/add0/c3 ;
  wire \u1_Driver/add0/c7 ;
  wire \u1_Driver/add1/c11 ;
  wire \u1_Driver/add1/c3 ;
  wire \u1_Driver/add1/c7 ;
  wire \u1_Driver/lcd_request ;  // source/rtl/Driver.v(46)
  wire \u1_Driver/lt0_c1 ;
  wire \u1_Driver/lt0_c11 ;
  wire \u1_Driver/lt0_c3 ;
  wire \u1_Driver/lt0_c5 ;
  wire \u1_Driver/lt0_c7 ;
  wire \u1_Driver/lt0_c9 ;
  wire \u1_Driver/lt1_c1 ;
  wire \u1_Driver/lt1_c11 ;
  wire \u1_Driver/lt1_c3 ;
  wire \u1_Driver/lt1_c5 ;
  wire \u1_Driver/lt1_c7 ;
  wire \u1_Driver/lt1_c9 ;
  wire \u1_Driver/lt2_c1 ;
  wire \u1_Driver/lt2_c11 ;
  wire \u1_Driver/lt2_c3 ;
  wire \u1_Driver/lt2_c5 ;
  wire \u1_Driver/lt2_c7 ;
  wire \u1_Driver/lt2_c9 ;
  wire \u1_Driver/lt3_c1 ;
  wire \u1_Driver/lt3_c11 ;
  wire \u1_Driver/lt3_c3 ;
  wire \u1_Driver/lt3_c5 ;
  wire \u1_Driver/lt3_c7 ;
  wire \u1_Driver/lt3_c9 ;
  wire \u1_Driver/lt4_c1 ;
  wire \u1_Driver/lt4_c11 ;
  wire \u1_Driver/lt4_c3 ;
  wire \u1_Driver/lt4_c5 ;
  wire \u1_Driver/lt4_c7 ;
  wire \u1_Driver/lt4_c9 ;
  wire \u1_Driver/lt5_c1 ;
  wire \u1_Driver/lt5_c11 ;
  wire \u1_Driver/lt5_c3 ;
  wire \u1_Driver/lt5_c5 ;
  wire \u1_Driver/lt5_c7 ;
  wire \u1_Driver/lt5_c9 ;
  wire \u1_Driver/lt6_c1 ;
  wire \u1_Driver/lt6_c11 ;
  wire \u1_Driver/lt6_c3 ;
  wire \u1_Driver/lt6_c5 ;
  wire \u1_Driver/lt6_c7 ;
  wire \u1_Driver/lt6_c9 ;
  wire \u1_Driver/lt7_c1 ;
  wire \u1_Driver/lt7_c11 ;
  wire \u1_Driver/lt7_c3 ;
  wire \u1_Driver/lt7_c5 ;
  wire \u1_Driver/lt7_c7 ;
  wire \u1_Driver/lt7_c9 ;
  wire \u1_Driver/lt8_c1 ;
  wire \u1_Driver/lt8_c11 ;
  wire \u1_Driver/lt8_c3 ;
  wire \u1_Driver/lt8_c5 ;
  wire \u1_Driver/lt8_c7 ;
  wire \u1_Driver/lt8_c9 ;
  wire \u1_Driver/n1 ;
  wire \u1_Driver/n10 ;
  wire \u1_Driver/n11 ;
  wire \u1_Driver/n12 ;
  wire \u1_Driver/n14 ;
  wire \u1_Driver/n15 ;
  wire \u1_Driver/n17 ;
  wire \u1_Driver/n18 ;
  wire \u1_Driver/n4 ;
  wire \u1_Driver/n5 ;
  wire \u1_Driver/n6_lutinv ;
  wire \u1_Driver/sub0/c11 ;
  wire \u1_Driver/sub0/c3 ;
  wire \u1_Driver/sub0/c7 ;
  wire \u1_Driver/sub1/c11 ;
  wire \u1_Driver/sub1/c3 ;
  wire \u1_Driver/sub1/c7 ;
  wire \u2_Display/add0/c11 ;
  wire \u2_Display/add0/c15 ;
  wire \u2_Display/add0/c19 ;
  wire \u2_Display/add0/c23 ;
  wire \u2_Display/add0/c27 ;
  wire \u2_Display/add0/c3 ;
  wire \u2_Display/add0/c7 ;
  wire \u2_Display/add1/c11 ;
  wire \u2_Display/add1/c15 ;
  wire \u2_Display/add1/c19 ;
  wire \u2_Display/add1/c23 ;
  wire \u2_Display/add1/c27 ;
  wire \u2_Display/add1/c3 ;
  wire \u2_Display/add1/c31 ;
  wire \u2_Display/add1/c7 ;
  wire \u2_Display/add100/c11 ;
  wire \u2_Display/add100/c15 ;
  wire \u2_Display/add100/c19 ;
  wire \u2_Display/add100/c23 ;
  wire \u2_Display/add100/c27 ;
  wire \u2_Display/add100/c3 ;
  wire \u2_Display/add100/c31 ;
  wire \u2_Display/add100/c7 ;
  wire \u2_Display/add101/c11 ;
  wire \u2_Display/add101/c15 ;
  wire \u2_Display/add101/c19 ;
  wire \u2_Display/add101/c23 ;
  wire \u2_Display/add101/c27 ;
  wire \u2_Display/add101/c3 ;
  wire \u2_Display/add101/c31 ;
  wire \u2_Display/add101/c7 ;
  wire \u2_Display/add102/c11 ;
  wire \u2_Display/add102/c15 ;
  wire \u2_Display/add102/c19 ;
  wire \u2_Display/add102/c23 ;
  wire \u2_Display/add102/c27 ;
  wire \u2_Display/add102/c3 ;
  wire \u2_Display/add102/c31 ;
  wire \u2_Display/add102/c7 ;
  wire \u2_Display/add103/c11 ;
  wire \u2_Display/add103/c15 ;
  wire \u2_Display/add103/c19 ;
  wire \u2_Display/add103/c23 ;
  wire \u2_Display/add103/c27 ;
  wire \u2_Display/add103/c3 ;
  wire \u2_Display/add103/c31 ;
  wire \u2_Display/add103/c7 ;
  wire \u2_Display/add104/c11 ;
  wire \u2_Display/add104/c15 ;
  wire \u2_Display/add104/c19 ;
  wire \u2_Display/add104/c23 ;
  wire \u2_Display/add104/c27 ;
  wire \u2_Display/add104/c3 ;
  wire \u2_Display/add104/c31 ;
  wire \u2_Display/add104/c7 ;
  wire \u2_Display/add105/c11 ;
  wire \u2_Display/add105/c15 ;
  wire \u2_Display/add105/c19 ;
  wire \u2_Display/add105/c23 ;
  wire \u2_Display/add105/c27 ;
  wire \u2_Display/add105/c3 ;
  wire \u2_Display/add105/c31 ;
  wire \u2_Display/add105/c7 ;
  wire \u2_Display/add106/c3 ;
  wire \u2_Display/add106/c7 ;
  wire \u2_Display/add117/c11 ;
  wire \u2_Display/add117/c15 ;
  wire \u2_Display/add117/c19 ;
  wire \u2_Display/add117/c23 ;
  wire \u2_Display/add117/c27 ;
  wire \u2_Display/add117/c3 ;
  wire \u2_Display/add117/c31 ;
  wire \u2_Display/add117/c7 ;
  wire \u2_Display/add118/c11 ;
  wire \u2_Display/add118/c15 ;
  wire \u2_Display/add118/c19 ;
  wire \u2_Display/add118/c23 ;
  wire \u2_Display/add118/c27 ;
  wire \u2_Display/add118/c3 ;
  wire \u2_Display/add118/c31 ;
  wire \u2_Display/add118/c7 ;
  wire \u2_Display/add119/c11 ;
  wire \u2_Display/add119/c15 ;
  wire \u2_Display/add119/c19 ;
  wire \u2_Display/add119/c23 ;
  wire \u2_Display/add119/c27 ;
  wire \u2_Display/add119/c3 ;
  wire \u2_Display/add119/c31 ;
  wire \u2_Display/add119/c7 ;
  wire \u2_Display/add120/c11 ;
  wire \u2_Display/add120/c15 ;
  wire \u2_Display/add120/c19 ;
  wire \u2_Display/add120/c23 ;
  wire \u2_Display/add120/c27 ;
  wire \u2_Display/add120/c3 ;
  wire \u2_Display/add120/c31 ;
  wire \u2_Display/add120/c7 ;
  wire \u2_Display/add121/c11 ;
  wire \u2_Display/add121/c15 ;
  wire \u2_Display/add121/c19 ;
  wire \u2_Display/add121/c23 ;
  wire \u2_Display/add121/c27 ;
  wire \u2_Display/add121/c3 ;
  wire \u2_Display/add121/c31 ;
  wire \u2_Display/add121/c7 ;
  wire \u2_Display/add122/c11 ;
  wire \u2_Display/add122/c15 ;
  wire \u2_Display/add122/c19 ;
  wire \u2_Display/add122/c23 ;
  wire \u2_Display/add122/c27 ;
  wire \u2_Display/add122/c3 ;
  wire \u2_Display/add122/c31 ;
  wire \u2_Display/add122/c7 ;
  wire \u2_Display/add123/c11 ;
  wire \u2_Display/add123/c15 ;
  wire \u2_Display/add123/c19 ;
  wire \u2_Display/add123/c23 ;
  wire \u2_Display/add123/c27 ;
  wire \u2_Display/add123/c3 ;
  wire \u2_Display/add123/c31 ;
  wire \u2_Display/add123/c7 ;
  wire \u2_Display/add124/c11 ;
  wire \u2_Display/add124/c15 ;
  wire \u2_Display/add124/c19 ;
  wire \u2_Display/add124/c23 ;
  wire \u2_Display/add124/c27 ;
  wire \u2_Display/add124/c3 ;
  wire \u2_Display/add124/c31 ;
  wire \u2_Display/add124/c7 ;
  wire \u2_Display/add125/c11 ;
  wire \u2_Display/add125/c15 ;
  wire \u2_Display/add125/c19 ;
  wire \u2_Display/add125/c23 ;
  wire \u2_Display/add125/c27 ;
  wire \u2_Display/add125/c3 ;
  wire \u2_Display/add125/c31 ;
  wire \u2_Display/add125/c7 ;
  wire \u2_Display/add126/c11 ;
  wire \u2_Display/add126/c15 ;
  wire \u2_Display/add126/c19 ;
  wire \u2_Display/add126/c23 ;
  wire \u2_Display/add126/c27 ;
  wire \u2_Display/add126/c3 ;
  wire \u2_Display/add126/c31 ;
  wire \u2_Display/add126/c7 ;
  wire \u2_Display/add127/c11 ;
  wire \u2_Display/add127/c15 ;
  wire \u2_Display/add127/c19 ;
  wire \u2_Display/add127/c23 ;
  wire \u2_Display/add127/c27 ;
  wire \u2_Display/add127/c3 ;
  wire \u2_Display/add127/c31 ;
  wire \u2_Display/add127/c7 ;
  wire \u2_Display/add128/c11 ;
  wire \u2_Display/add128/c15 ;
  wire \u2_Display/add128/c19 ;
  wire \u2_Display/add128/c23 ;
  wire \u2_Display/add128/c27 ;
  wire \u2_Display/add128/c3 ;
  wire \u2_Display/add128/c31 ;
  wire \u2_Display/add128/c7 ;
  wire \u2_Display/add129/c11 ;
  wire \u2_Display/add129/c15 ;
  wire \u2_Display/add129/c19 ;
  wire \u2_Display/add129/c23 ;
  wire \u2_Display/add129/c27 ;
  wire \u2_Display/add129/c3 ;
  wire \u2_Display/add129/c31 ;
  wire \u2_Display/add129/c7 ;
  wire \u2_Display/add130/c11 ;
  wire \u2_Display/add130/c15 ;
  wire \u2_Display/add130/c19 ;
  wire \u2_Display/add130/c23 ;
  wire \u2_Display/add130/c27 ;
  wire \u2_Display/add130/c3 ;
  wire \u2_Display/add130/c31 ;
  wire \u2_Display/add130/c7 ;
  wire \u2_Display/add131/c11 ;
  wire \u2_Display/add131/c15 ;
  wire \u2_Display/add131/c19 ;
  wire \u2_Display/add131/c23 ;
  wire \u2_Display/add131/c27 ;
  wire \u2_Display/add131/c3 ;
  wire \u2_Display/add131/c31 ;
  wire \u2_Display/add131/c7 ;
  wire \u2_Display/add132/c11 ;
  wire \u2_Display/add132/c15 ;
  wire \u2_Display/add132/c19 ;
  wire \u2_Display/add132/c23 ;
  wire \u2_Display/add132/c27 ;
  wire \u2_Display/add132/c3 ;
  wire \u2_Display/add132/c31 ;
  wire \u2_Display/add132/c7 ;
  wire \u2_Display/add133/c11 ;
  wire \u2_Display/add133/c15 ;
  wire \u2_Display/add133/c19 ;
  wire \u2_Display/add133/c23 ;
  wire \u2_Display/add133/c27 ;
  wire \u2_Display/add133/c3 ;
  wire \u2_Display/add133/c31 ;
  wire \u2_Display/add133/c7 ;
  wire \u2_Display/add134/c11 ;
  wire \u2_Display/add134/c15 ;
  wire \u2_Display/add134/c19 ;
  wire \u2_Display/add134/c23 ;
  wire \u2_Display/add134/c27 ;
  wire \u2_Display/add134/c3 ;
  wire \u2_Display/add134/c31 ;
  wire \u2_Display/add134/c7 ;
  wire \u2_Display/add135/c11 ;
  wire \u2_Display/add135/c15 ;
  wire \u2_Display/add135/c19 ;
  wire \u2_Display/add135/c23 ;
  wire \u2_Display/add135/c27 ;
  wire \u2_Display/add135/c3 ;
  wire \u2_Display/add135/c31 ;
  wire \u2_Display/add135/c7 ;
  wire \u2_Display/add136/c11 ;
  wire \u2_Display/add136/c15 ;
  wire \u2_Display/add136/c19 ;
  wire \u2_Display/add136/c23 ;
  wire \u2_Display/add136/c27 ;
  wire \u2_Display/add136/c3 ;
  wire \u2_Display/add136/c31 ;
  wire \u2_Display/add136/c7 ;
  wire \u2_Display/add137/c11 ;
  wire \u2_Display/add137/c15 ;
  wire \u2_Display/add137/c19 ;
  wire \u2_Display/add137/c23 ;
  wire \u2_Display/add137/c27 ;
  wire \u2_Display/add137/c3 ;
  wire \u2_Display/add137/c31 ;
  wire \u2_Display/add137/c7 ;
  wire \u2_Display/add138/c11 ;
  wire \u2_Display/add138/c15 ;
  wire \u2_Display/add138/c19 ;
  wire \u2_Display/add138/c23 ;
  wire \u2_Display/add138/c27 ;
  wire \u2_Display/add138/c3 ;
  wire \u2_Display/add138/c31 ;
  wire \u2_Display/add138/c7 ;
  wire \u2_Display/add139/c3 ;
  wire \u2_Display/add139/c7 ;
  wire \u2_Display/add14/c11 ;
  wire \u2_Display/add14/c15 ;
  wire \u2_Display/add14/c19 ;
  wire \u2_Display/add14/c23 ;
  wire \u2_Display/add14/c27 ;
  wire \u2_Display/add14/c3 ;
  wire \u2_Display/add14/c31 ;
  wire \u2_Display/add14/c7 ;
  wire \u2_Display/add151/c11 ;
  wire \u2_Display/add151/c15 ;
  wire \u2_Display/add151/c19 ;
  wire \u2_Display/add151/c23 ;
  wire \u2_Display/add151/c27 ;
  wire \u2_Display/add151/c3 ;
  wire \u2_Display/add151/c31 ;
  wire \u2_Display/add151/c7 ;
  wire \u2_Display/add152/c11 ;
  wire \u2_Display/add152/c15 ;
  wire \u2_Display/add152/c19 ;
  wire \u2_Display/add152/c23 ;
  wire \u2_Display/add152/c27 ;
  wire \u2_Display/add152/c3 ;
  wire \u2_Display/add152/c31 ;
  wire \u2_Display/add152/c7 ;
  wire \u2_Display/add153/c11 ;
  wire \u2_Display/add153/c15 ;
  wire \u2_Display/add153/c19 ;
  wire \u2_Display/add153/c23 ;
  wire \u2_Display/add153/c27 ;
  wire \u2_Display/add153/c3 ;
  wire \u2_Display/add153/c31 ;
  wire \u2_Display/add153/c7 ;
  wire \u2_Display/add154/c11 ;
  wire \u2_Display/add154/c15 ;
  wire \u2_Display/add154/c19 ;
  wire \u2_Display/add154/c23 ;
  wire \u2_Display/add154/c27 ;
  wire \u2_Display/add154/c3 ;
  wire \u2_Display/add154/c31 ;
  wire \u2_Display/add154/c7 ;
  wire \u2_Display/add155/c11 ;
  wire \u2_Display/add155/c15 ;
  wire \u2_Display/add155/c19 ;
  wire \u2_Display/add155/c23 ;
  wire \u2_Display/add155/c27 ;
  wire \u2_Display/add155/c3 ;
  wire \u2_Display/add155/c31 ;
  wire \u2_Display/add155/c7 ;
  wire \u2_Display/add156/c11 ;
  wire \u2_Display/add156/c15 ;
  wire \u2_Display/add156/c19 ;
  wire \u2_Display/add156/c23 ;
  wire \u2_Display/add156/c27 ;
  wire \u2_Display/add156/c3 ;
  wire \u2_Display/add156/c31 ;
  wire \u2_Display/add156/c7 ;
  wire \u2_Display/add157/c11 ;
  wire \u2_Display/add157/c15 ;
  wire \u2_Display/add157/c19 ;
  wire \u2_Display/add157/c23 ;
  wire \u2_Display/add157/c27 ;
  wire \u2_Display/add157/c3 ;
  wire \u2_Display/add157/c31 ;
  wire \u2_Display/add157/c7 ;
  wire \u2_Display/add158/c11 ;
  wire \u2_Display/add158/c15 ;
  wire \u2_Display/add158/c19 ;
  wire \u2_Display/add158/c23 ;
  wire \u2_Display/add158/c27 ;
  wire \u2_Display/add158/c3 ;
  wire \u2_Display/add158/c31 ;
  wire \u2_Display/add158/c7 ;
  wire \u2_Display/add159/c11 ;
  wire \u2_Display/add159/c15 ;
  wire \u2_Display/add159/c19 ;
  wire \u2_Display/add159/c23 ;
  wire \u2_Display/add159/c27 ;
  wire \u2_Display/add159/c3 ;
  wire \u2_Display/add159/c31 ;
  wire \u2_Display/add159/c7 ;
  wire \u2_Display/add160/c11 ;
  wire \u2_Display/add160/c15 ;
  wire \u2_Display/add160/c19 ;
  wire \u2_Display/add160/c23 ;
  wire \u2_Display/add160/c27 ;
  wire \u2_Display/add160/c3 ;
  wire \u2_Display/add160/c31 ;
  wire \u2_Display/add160/c7 ;
  wire \u2_Display/add161/c11 ;
  wire \u2_Display/add161/c15 ;
  wire \u2_Display/add161/c19 ;
  wire \u2_Display/add161/c23 ;
  wire \u2_Display/add161/c27 ;
  wire \u2_Display/add161/c3 ;
  wire \u2_Display/add161/c31 ;
  wire \u2_Display/add161/c7 ;
  wire \u2_Display/add162/c11 ;
  wire \u2_Display/add162/c15 ;
  wire \u2_Display/add162/c19 ;
  wire \u2_Display/add162/c23 ;
  wire \u2_Display/add162/c27 ;
  wire \u2_Display/add162/c3 ;
  wire \u2_Display/add162/c31 ;
  wire \u2_Display/add162/c7 ;
  wire \u2_Display/add163/c11 ;
  wire \u2_Display/add163/c15 ;
  wire \u2_Display/add163/c19 ;
  wire \u2_Display/add163/c23 ;
  wire \u2_Display/add163/c27 ;
  wire \u2_Display/add163/c3 ;
  wire \u2_Display/add163/c31 ;
  wire \u2_Display/add163/c7 ;
  wire \u2_Display/add164/c11 ;
  wire \u2_Display/add164/c15 ;
  wire \u2_Display/add164/c19 ;
  wire \u2_Display/add164/c23 ;
  wire \u2_Display/add164/c27 ;
  wire \u2_Display/add164/c3 ;
  wire \u2_Display/add164/c31 ;
  wire \u2_Display/add164/c7 ;
  wire \u2_Display/add165/c11 ;
  wire \u2_Display/add165/c15 ;
  wire \u2_Display/add165/c19 ;
  wire \u2_Display/add165/c23 ;
  wire \u2_Display/add165/c27 ;
  wire \u2_Display/add165/c3 ;
  wire \u2_Display/add165/c31 ;
  wire \u2_Display/add165/c7 ;
  wire \u2_Display/add166/c11 ;
  wire \u2_Display/add166/c15 ;
  wire \u2_Display/add166/c19 ;
  wire \u2_Display/add166/c23 ;
  wire \u2_Display/add166/c27 ;
  wire \u2_Display/add166/c3 ;
  wire \u2_Display/add166/c31 ;
  wire \u2_Display/add166/c7 ;
  wire \u2_Display/add167/c11 ;
  wire \u2_Display/add167/c15 ;
  wire \u2_Display/add167/c19 ;
  wire \u2_Display/add167/c23 ;
  wire \u2_Display/add167/c27 ;
  wire \u2_Display/add167/c3 ;
  wire \u2_Display/add167/c31 ;
  wire \u2_Display/add167/c7 ;
  wire \u2_Display/add168/c11 ;
  wire \u2_Display/add168/c15 ;
  wire \u2_Display/add168/c19 ;
  wire \u2_Display/add168/c23 ;
  wire \u2_Display/add168/c27 ;
  wire \u2_Display/add168/c3 ;
  wire \u2_Display/add168/c31 ;
  wire \u2_Display/add168/c7 ;
  wire \u2_Display/add169/c11 ;
  wire \u2_Display/add169/c15 ;
  wire \u2_Display/add169/c19 ;
  wire \u2_Display/add169/c23 ;
  wire \u2_Display/add169/c27 ;
  wire \u2_Display/add169/c3 ;
  wire \u2_Display/add169/c31 ;
  wire \u2_Display/add169/c7 ;
  wire \u2_Display/add170/c11 ;
  wire \u2_Display/add170/c15 ;
  wire \u2_Display/add170/c19 ;
  wire \u2_Display/add170/c23 ;
  wire \u2_Display/add170/c27 ;
  wire \u2_Display/add170/c3 ;
  wire \u2_Display/add170/c31 ;
  wire \u2_Display/add170/c7 ;
  wire \u2_Display/add171/c11 ;
  wire \u2_Display/add171/c15 ;
  wire \u2_Display/add171/c19 ;
  wire \u2_Display/add171/c23 ;
  wire \u2_Display/add171/c27 ;
  wire \u2_Display/add171/c3 ;
  wire \u2_Display/add171/c31 ;
  wire \u2_Display/add171/c7 ;
  wire \u2_Display/add172/c3 ;
  wire \u2_Display/add172/c7 ;
  wire \u2_Display/add18/c11 ;
  wire \u2_Display/add18/c15 ;
  wire \u2_Display/add18/c19 ;
  wire \u2_Display/add18/c23 ;
  wire \u2_Display/add18/c27 ;
  wire \u2_Display/add18/c3 ;
  wire \u2_Display/add18/c31 ;
  wire \u2_Display/add18/c7 ;
  wire \u2_Display/add19/c11 ;
  wire \u2_Display/add19/c15 ;
  wire \u2_Display/add19/c19 ;
  wire \u2_Display/add19/c23 ;
  wire \u2_Display/add19/c27 ;
  wire \u2_Display/add19/c3 ;
  wire \u2_Display/add19/c31 ;
  wire \u2_Display/add19/c7 ;
  wire \u2_Display/add20/c11 ;
  wire \u2_Display/add20/c15 ;
  wire \u2_Display/add20/c19 ;
  wire \u2_Display/add20/c23 ;
  wire \u2_Display/add20/c27 ;
  wire \u2_Display/add20/c3 ;
  wire \u2_Display/add20/c31 ;
  wire \u2_Display/add20/c7 ;
  wire \u2_Display/add21/c11 ;
  wire \u2_Display/add21/c15 ;
  wire \u2_Display/add21/c19 ;
  wire \u2_Display/add21/c23 ;
  wire \u2_Display/add21/c27 ;
  wire \u2_Display/add21/c3 ;
  wire \u2_Display/add21/c31 ;
  wire \u2_Display/add21/c7 ;
  wire \u2_Display/add22/c11 ;
  wire \u2_Display/add22/c15 ;
  wire \u2_Display/add22/c19 ;
  wire \u2_Display/add22/c23 ;
  wire \u2_Display/add22/c27 ;
  wire \u2_Display/add22/c3 ;
  wire \u2_Display/add22/c31 ;
  wire \u2_Display/add22/c7 ;
  wire \u2_Display/add23/c11 ;
  wire \u2_Display/add23/c15 ;
  wire \u2_Display/add23/c19 ;
  wire \u2_Display/add23/c23 ;
  wire \u2_Display/add23/c27 ;
  wire \u2_Display/add23/c3 ;
  wire \u2_Display/add23/c31 ;
  wire \u2_Display/add23/c7 ;
  wire \u2_Display/add24/c11 ;
  wire \u2_Display/add24/c15 ;
  wire \u2_Display/add24/c19 ;
  wire \u2_Display/add24/c23 ;
  wire \u2_Display/add24/c27 ;
  wire \u2_Display/add24/c3 ;
  wire \u2_Display/add24/c31 ;
  wire \u2_Display/add24/c7 ;
  wire \u2_Display/add25/c11 ;
  wire \u2_Display/add25/c15 ;
  wire \u2_Display/add25/c19 ;
  wire \u2_Display/add25/c23 ;
  wire \u2_Display/add25/c27 ;
  wire \u2_Display/add25/c3 ;
  wire \u2_Display/add25/c31 ;
  wire \u2_Display/add25/c7 ;
  wire \u2_Display/add26/c11 ;
  wire \u2_Display/add26/c15 ;
  wire \u2_Display/add26/c19 ;
  wire \u2_Display/add26/c23 ;
  wire \u2_Display/add26/c27 ;
  wire \u2_Display/add26/c3 ;
  wire \u2_Display/add26/c31 ;
  wire \u2_Display/add26/c7 ;
  wire \u2_Display/add27/c11 ;
  wire \u2_Display/add27/c15 ;
  wire \u2_Display/add27/c19 ;
  wire \u2_Display/add27/c23 ;
  wire \u2_Display/add27/c27 ;
  wire \u2_Display/add27/c3 ;
  wire \u2_Display/add27/c31 ;
  wire \u2_Display/add27/c7 ;
  wire \u2_Display/add28/c11 ;
  wire \u2_Display/add28/c15 ;
  wire \u2_Display/add28/c19 ;
  wire \u2_Display/add28/c23 ;
  wire \u2_Display/add28/c27 ;
  wire \u2_Display/add28/c3 ;
  wire \u2_Display/add28/c31 ;
  wire \u2_Display/add28/c7 ;
  wire \u2_Display/add29/c11 ;
  wire \u2_Display/add29/c15 ;
  wire \u2_Display/add29/c19 ;
  wire \u2_Display/add29/c23 ;
  wire \u2_Display/add29/c27 ;
  wire \u2_Display/add29/c3 ;
  wire \u2_Display/add29/c31 ;
  wire \u2_Display/add29/c7 ;
  wire \u2_Display/add2_2/c1 ;
  wire \u2_Display/add2_2/c3 ;
  wire \u2_Display/add2_2_co ;
  wire \u2_Display/add30/c11 ;
  wire \u2_Display/add30/c15 ;
  wire \u2_Display/add30/c19 ;
  wire \u2_Display/add30/c23 ;
  wire \u2_Display/add30/c27 ;
  wire \u2_Display/add30/c3 ;
  wire \u2_Display/add30/c31 ;
  wire \u2_Display/add30/c7 ;
  wire \u2_Display/add31/c11 ;
  wire \u2_Display/add31/c15 ;
  wire \u2_Display/add31/c19 ;
  wire \u2_Display/add31/c23 ;
  wire \u2_Display/add31/c27 ;
  wire \u2_Display/add31/c3 ;
  wire \u2_Display/add31/c31 ;
  wire \u2_Display/add31/c7 ;
  wire \u2_Display/add32/c11 ;
  wire \u2_Display/add32/c15 ;
  wire \u2_Display/add32/c19 ;
  wire \u2_Display/add32/c23 ;
  wire \u2_Display/add32/c27 ;
  wire \u2_Display/add32/c3 ;
  wire \u2_Display/add32/c31 ;
  wire \u2_Display/add32/c7 ;
  wire \u2_Display/add33/c11 ;
  wire \u2_Display/add33/c15 ;
  wire \u2_Display/add33/c19 ;
  wire \u2_Display/add33/c23 ;
  wire \u2_Display/add33/c27 ;
  wire \u2_Display/add33/c3 ;
  wire \u2_Display/add33/c31 ;
  wire \u2_Display/add33/c7 ;
  wire \u2_Display/add34/c11 ;
  wire \u2_Display/add34/c15 ;
  wire \u2_Display/add34/c19 ;
  wire \u2_Display/add34/c23 ;
  wire \u2_Display/add34/c27 ;
  wire \u2_Display/add34/c3 ;
  wire \u2_Display/add34/c31 ;
  wire \u2_Display/add34/c7 ;
  wire \u2_Display/add35/c11 ;
  wire \u2_Display/add35/c15 ;
  wire \u2_Display/add35/c19 ;
  wire \u2_Display/add35/c23 ;
  wire \u2_Display/add35/c27 ;
  wire \u2_Display/add35/c3 ;
  wire \u2_Display/add35/c31 ;
  wire \u2_Display/add35/c7 ;
  wire \u2_Display/add36/c11 ;
  wire \u2_Display/add36/c15 ;
  wire \u2_Display/add36/c19 ;
  wire \u2_Display/add36/c23 ;
  wire \u2_Display/add36/c27 ;
  wire \u2_Display/add36/c3 ;
  wire \u2_Display/add36/c31 ;
  wire \u2_Display/add36/c7 ;
  wire \u2_Display/add37/c11 ;
  wire \u2_Display/add37/c15 ;
  wire \u2_Display/add37/c19 ;
  wire \u2_Display/add37/c23 ;
  wire \u2_Display/add37/c27 ;
  wire \u2_Display/add37/c3 ;
  wire \u2_Display/add37/c31 ;
  wire \u2_Display/add37/c7 ;
  wire \u2_Display/add38/c11 ;
  wire \u2_Display/add38/c15 ;
  wire \u2_Display/add38/c19 ;
  wire \u2_Display/add38/c23 ;
  wire \u2_Display/add38/c27 ;
  wire \u2_Display/add38/c3 ;
  wire \u2_Display/add38/c31 ;
  wire \u2_Display/add38/c7 ;
  wire \u2_Display/add39/c11 ;
  wire \u2_Display/add39/c15 ;
  wire \u2_Display/add39/c19 ;
  wire \u2_Display/add39/c23 ;
  wire \u2_Display/add39/c27 ;
  wire \u2_Display/add39/c3 ;
  wire \u2_Display/add39/c31 ;
  wire \u2_Display/add39/c7 ;
  wire \u2_Display/add40/c3 ;
  wire \u2_Display/add40/c7 ;
  wire \u2_Display/add4_2/c1 ;
  wire \u2_Display/add4_2/c3 ;
  wire \u2_Display/add4_2_co ;
  wire \u2_Display/add51/c11 ;
  wire \u2_Display/add51/c15 ;
  wire \u2_Display/add51/c19 ;
  wire \u2_Display/add51/c23 ;
  wire \u2_Display/add51/c27 ;
  wire \u2_Display/add51/c3 ;
  wire \u2_Display/add51/c31 ;
  wire \u2_Display/add51/c7 ;
  wire \u2_Display/add52/c11 ;
  wire \u2_Display/add52/c15 ;
  wire \u2_Display/add52/c19 ;
  wire \u2_Display/add52/c23 ;
  wire \u2_Display/add52/c27 ;
  wire \u2_Display/add52/c3 ;
  wire \u2_Display/add52/c31 ;
  wire \u2_Display/add52/c7 ;
  wire \u2_Display/add53/c11 ;
  wire \u2_Display/add53/c15 ;
  wire \u2_Display/add53/c19 ;
  wire \u2_Display/add53/c23 ;
  wire \u2_Display/add53/c27 ;
  wire \u2_Display/add53/c3 ;
  wire \u2_Display/add53/c31 ;
  wire \u2_Display/add53/c7 ;
  wire \u2_Display/add54/c11 ;
  wire \u2_Display/add54/c15 ;
  wire \u2_Display/add54/c19 ;
  wire \u2_Display/add54/c23 ;
  wire \u2_Display/add54/c27 ;
  wire \u2_Display/add54/c3 ;
  wire \u2_Display/add54/c31 ;
  wire \u2_Display/add54/c7 ;
  wire \u2_Display/add55/c11 ;
  wire \u2_Display/add55/c15 ;
  wire \u2_Display/add55/c19 ;
  wire \u2_Display/add55/c23 ;
  wire \u2_Display/add55/c27 ;
  wire \u2_Display/add55/c3 ;
  wire \u2_Display/add55/c31 ;
  wire \u2_Display/add55/c7 ;
  wire \u2_Display/add56/c11 ;
  wire \u2_Display/add56/c15 ;
  wire \u2_Display/add56/c19 ;
  wire \u2_Display/add56/c23 ;
  wire \u2_Display/add56/c27 ;
  wire \u2_Display/add56/c3 ;
  wire \u2_Display/add56/c31 ;
  wire \u2_Display/add56/c7 ;
  wire \u2_Display/add57/c11 ;
  wire \u2_Display/add57/c15 ;
  wire \u2_Display/add57/c19 ;
  wire \u2_Display/add57/c23 ;
  wire \u2_Display/add57/c27 ;
  wire \u2_Display/add57/c3 ;
  wire \u2_Display/add57/c31 ;
  wire \u2_Display/add57/c7 ;
  wire \u2_Display/add58/c11 ;
  wire \u2_Display/add58/c15 ;
  wire \u2_Display/add58/c19 ;
  wire \u2_Display/add58/c23 ;
  wire \u2_Display/add58/c27 ;
  wire \u2_Display/add58/c3 ;
  wire \u2_Display/add58/c31 ;
  wire \u2_Display/add58/c7 ;
  wire \u2_Display/add59/c11 ;
  wire \u2_Display/add59/c15 ;
  wire \u2_Display/add59/c19 ;
  wire \u2_Display/add59/c23 ;
  wire \u2_Display/add59/c27 ;
  wire \u2_Display/add59/c3 ;
  wire \u2_Display/add59/c31 ;
  wire \u2_Display/add59/c7 ;
  wire \u2_Display/add60/c11 ;
  wire \u2_Display/add60/c15 ;
  wire \u2_Display/add60/c19 ;
  wire \u2_Display/add60/c23 ;
  wire \u2_Display/add60/c27 ;
  wire \u2_Display/add60/c3 ;
  wire \u2_Display/add60/c31 ;
  wire \u2_Display/add60/c7 ;
  wire \u2_Display/add61/c11 ;
  wire \u2_Display/add61/c15 ;
  wire \u2_Display/add61/c19 ;
  wire \u2_Display/add61/c23 ;
  wire \u2_Display/add61/c27 ;
  wire \u2_Display/add61/c3 ;
  wire \u2_Display/add61/c31 ;
  wire \u2_Display/add61/c7 ;
  wire \u2_Display/add62/c11 ;
  wire \u2_Display/add62/c15 ;
  wire \u2_Display/add62/c19 ;
  wire \u2_Display/add62/c23 ;
  wire \u2_Display/add62/c27 ;
  wire \u2_Display/add62/c3 ;
  wire \u2_Display/add62/c31 ;
  wire \u2_Display/add62/c7 ;
  wire \u2_Display/add63/c11 ;
  wire \u2_Display/add63/c15 ;
  wire \u2_Display/add63/c19 ;
  wire \u2_Display/add63/c23 ;
  wire \u2_Display/add63/c27 ;
  wire \u2_Display/add63/c3 ;
  wire \u2_Display/add63/c31 ;
  wire \u2_Display/add63/c7 ;
  wire \u2_Display/add64/c11 ;
  wire \u2_Display/add64/c15 ;
  wire \u2_Display/add64/c19 ;
  wire \u2_Display/add64/c23 ;
  wire \u2_Display/add64/c27 ;
  wire \u2_Display/add64/c3 ;
  wire \u2_Display/add64/c31 ;
  wire \u2_Display/add64/c7 ;
  wire \u2_Display/add65/c11 ;
  wire \u2_Display/add65/c15 ;
  wire \u2_Display/add65/c19 ;
  wire \u2_Display/add65/c23 ;
  wire \u2_Display/add65/c27 ;
  wire \u2_Display/add65/c3 ;
  wire \u2_Display/add65/c31 ;
  wire \u2_Display/add65/c7 ;
  wire \u2_Display/add66/c11 ;
  wire \u2_Display/add66/c15 ;
  wire \u2_Display/add66/c19 ;
  wire \u2_Display/add66/c23 ;
  wire \u2_Display/add66/c27 ;
  wire \u2_Display/add66/c3 ;
  wire \u2_Display/add66/c31 ;
  wire \u2_Display/add66/c7 ;
  wire \u2_Display/add67/c11 ;
  wire \u2_Display/add67/c15 ;
  wire \u2_Display/add67/c19 ;
  wire \u2_Display/add67/c23 ;
  wire \u2_Display/add67/c27 ;
  wire \u2_Display/add67/c3 ;
  wire \u2_Display/add67/c31 ;
  wire \u2_Display/add67/c7 ;
  wire \u2_Display/add68/c11 ;
  wire \u2_Display/add68/c15 ;
  wire \u2_Display/add68/c19 ;
  wire \u2_Display/add68/c23 ;
  wire \u2_Display/add68/c27 ;
  wire \u2_Display/add68/c3 ;
  wire \u2_Display/add68/c31 ;
  wire \u2_Display/add68/c7 ;
  wire \u2_Display/add69/c11 ;
  wire \u2_Display/add69/c15 ;
  wire \u2_Display/add69/c19 ;
  wire \u2_Display/add69/c23 ;
  wire \u2_Display/add69/c27 ;
  wire \u2_Display/add69/c3 ;
  wire \u2_Display/add69/c31 ;
  wire \u2_Display/add69/c7 ;
  wire \u2_Display/add6_2/c1 ;
  wire \u2_Display/add6_2/c3 ;
  wire \u2_Display/add6_2_co ;
  wire \u2_Display/add70/c11 ;
  wire \u2_Display/add70/c15 ;
  wire \u2_Display/add70/c19 ;
  wire \u2_Display/add70/c23 ;
  wire \u2_Display/add70/c27 ;
  wire \u2_Display/add70/c3 ;
  wire \u2_Display/add70/c31 ;
  wire \u2_Display/add70/c7 ;
  wire \u2_Display/add71/c11 ;
  wire \u2_Display/add71/c15 ;
  wire \u2_Display/add71/c19 ;
  wire \u2_Display/add71/c23 ;
  wire \u2_Display/add71/c27 ;
  wire \u2_Display/add71/c3 ;
  wire \u2_Display/add71/c31 ;
  wire \u2_Display/add71/c7 ;
  wire \u2_Display/add72/c11 ;
  wire \u2_Display/add72/c15 ;
  wire \u2_Display/add72/c19 ;
  wire \u2_Display/add72/c23 ;
  wire \u2_Display/add72/c27 ;
  wire \u2_Display/add72/c3 ;
  wire \u2_Display/add72/c31 ;
  wire \u2_Display/add72/c7 ;
  wire \u2_Display/add73/c3 ;
  wire \u2_Display/add73/c7 ;
  wire \u2_Display/add7_2_co ;
  wire \u2_Display/add84/c11 ;
  wire \u2_Display/add84/c15 ;
  wire \u2_Display/add84/c19 ;
  wire \u2_Display/add84/c23 ;
  wire \u2_Display/add84/c27 ;
  wire \u2_Display/add84/c3 ;
  wire \u2_Display/add84/c31 ;
  wire \u2_Display/add84/c7 ;
  wire \u2_Display/add85/c11 ;
  wire \u2_Display/add85/c15 ;
  wire \u2_Display/add85/c19 ;
  wire \u2_Display/add85/c23 ;
  wire \u2_Display/add85/c27 ;
  wire \u2_Display/add85/c3 ;
  wire \u2_Display/add85/c31 ;
  wire \u2_Display/add85/c7 ;
  wire \u2_Display/add86/c11 ;
  wire \u2_Display/add86/c15 ;
  wire \u2_Display/add86/c19 ;
  wire \u2_Display/add86/c23 ;
  wire \u2_Display/add86/c27 ;
  wire \u2_Display/add86/c3 ;
  wire \u2_Display/add86/c31 ;
  wire \u2_Display/add86/c7 ;
  wire \u2_Display/add87/c11 ;
  wire \u2_Display/add87/c15 ;
  wire \u2_Display/add87/c19 ;
  wire \u2_Display/add87/c23 ;
  wire \u2_Display/add87/c27 ;
  wire \u2_Display/add87/c3 ;
  wire \u2_Display/add87/c31 ;
  wire \u2_Display/add87/c7 ;
  wire \u2_Display/add88/c11 ;
  wire \u2_Display/add88/c15 ;
  wire \u2_Display/add88/c19 ;
  wire \u2_Display/add88/c23 ;
  wire \u2_Display/add88/c27 ;
  wire \u2_Display/add88/c3 ;
  wire \u2_Display/add88/c31 ;
  wire \u2_Display/add88/c7 ;
  wire \u2_Display/add89/c11 ;
  wire \u2_Display/add89/c15 ;
  wire \u2_Display/add89/c19 ;
  wire \u2_Display/add89/c23 ;
  wire \u2_Display/add89/c27 ;
  wire \u2_Display/add89/c3 ;
  wire \u2_Display/add89/c31 ;
  wire \u2_Display/add89/c7 ;
  wire \u2_Display/add90/c11 ;
  wire \u2_Display/add90/c15 ;
  wire \u2_Display/add90/c19 ;
  wire \u2_Display/add90/c23 ;
  wire \u2_Display/add90/c27 ;
  wire \u2_Display/add90/c3 ;
  wire \u2_Display/add90/c31 ;
  wire \u2_Display/add90/c7 ;
  wire \u2_Display/add91/c11 ;
  wire \u2_Display/add91/c15 ;
  wire \u2_Display/add91/c19 ;
  wire \u2_Display/add91/c23 ;
  wire \u2_Display/add91/c27 ;
  wire \u2_Display/add91/c3 ;
  wire \u2_Display/add91/c31 ;
  wire \u2_Display/add91/c7 ;
  wire \u2_Display/add92/c11 ;
  wire \u2_Display/add92/c15 ;
  wire \u2_Display/add92/c19 ;
  wire \u2_Display/add92/c23 ;
  wire \u2_Display/add92/c27 ;
  wire \u2_Display/add92/c3 ;
  wire \u2_Display/add92/c31 ;
  wire \u2_Display/add92/c7 ;
  wire \u2_Display/add93/c11 ;
  wire \u2_Display/add93/c15 ;
  wire \u2_Display/add93/c19 ;
  wire \u2_Display/add93/c23 ;
  wire \u2_Display/add93/c27 ;
  wire \u2_Display/add93/c3 ;
  wire \u2_Display/add93/c31 ;
  wire \u2_Display/add93/c7 ;
  wire \u2_Display/add94/c11 ;
  wire \u2_Display/add94/c15 ;
  wire \u2_Display/add94/c19 ;
  wire \u2_Display/add94/c23 ;
  wire \u2_Display/add94/c27 ;
  wire \u2_Display/add94/c3 ;
  wire \u2_Display/add94/c31 ;
  wire \u2_Display/add94/c7 ;
  wire \u2_Display/add95/c11 ;
  wire \u2_Display/add95/c15 ;
  wire \u2_Display/add95/c19 ;
  wire \u2_Display/add95/c23 ;
  wire \u2_Display/add95/c27 ;
  wire \u2_Display/add95/c3 ;
  wire \u2_Display/add95/c31 ;
  wire \u2_Display/add95/c7 ;
  wire \u2_Display/add96/c11 ;
  wire \u2_Display/add96/c15 ;
  wire \u2_Display/add96/c19 ;
  wire \u2_Display/add96/c23 ;
  wire \u2_Display/add96/c27 ;
  wire \u2_Display/add96/c3 ;
  wire \u2_Display/add96/c31 ;
  wire \u2_Display/add96/c7 ;
  wire \u2_Display/add97/c11 ;
  wire \u2_Display/add97/c15 ;
  wire \u2_Display/add97/c19 ;
  wire \u2_Display/add97/c23 ;
  wire \u2_Display/add97/c27 ;
  wire \u2_Display/add97/c3 ;
  wire \u2_Display/add97/c31 ;
  wire \u2_Display/add97/c7 ;
  wire \u2_Display/add98/c11 ;
  wire \u2_Display/add98/c15 ;
  wire \u2_Display/add98/c19 ;
  wire \u2_Display/add98/c23 ;
  wire \u2_Display/add98/c27 ;
  wire \u2_Display/add98/c3 ;
  wire \u2_Display/add98/c31 ;
  wire \u2_Display/add98/c7 ;
  wire \u2_Display/add99/c11 ;
  wire \u2_Display/add99/c15 ;
  wire \u2_Display/add99/c19 ;
  wire \u2_Display/add99/c23 ;
  wire \u2_Display/add99/c27 ;
  wire \u2_Display/add99/c3 ;
  wire \u2_Display/add99/c31 ;
  wire \u2_Display/add99/c7 ;
  wire \u2_Display/clk1s ;  // source/rtl/Display.v(46)
  wire \u2_Display/clk1s_gclk_net ;
  wire \u2_Display/lt0_2_c1 ;
  wire \u2_Display/lt0_2_c11 ;
  wire \u2_Display/lt0_2_c3 ;
  wire \u2_Display/lt0_2_c5 ;
  wire \u2_Display/lt0_2_c7 ;
  wire \u2_Display/lt0_2_c9 ;
  wire \u2_Display/lt100_c1 ;
  wire \u2_Display/lt100_c11 ;
  wire \u2_Display/lt100_c13 ;
  wire \u2_Display/lt100_c15 ;
  wire \u2_Display/lt100_c17 ;
  wire \u2_Display/lt100_c19 ;
  wire \u2_Display/lt100_c21 ;
  wire \u2_Display/lt100_c23 ;
  wire \u2_Display/lt100_c25 ;
  wire \u2_Display/lt100_c27 ;
  wire \u2_Display/lt100_c29 ;
  wire \u2_Display/lt100_c3 ;
  wire \u2_Display/lt100_c31 ;
  wire \u2_Display/lt100_c5 ;
  wire \u2_Display/lt100_c7 ;
  wire \u2_Display/lt100_c9 ;
  wire \u2_Display/lt101_c1 ;
  wire \u2_Display/lt101_c11 ;
  wire \u2_Display/lt101_c13 ;
  wire \u2_Display/lt101_c15 ;
  wire \u2_Display/lt101_c17 ;
  wire \u2_Display/lt101_c19 ;
  wire \u2_Display/lt101_c21 ;
  wire \u2_Display/lt101_c23 ;
  wire \u2_Display/lt101_c25 ;
  wire \u2_Display/lt101_c27 ;
  wire \u2_Display/lt101_c29 ;
  wire \u2_Display/lt101_c3 ;
  wire \u2_Display/lt101_c31 ;
  wire \u2_Display/lt101_c5 ;
  wire \u2_Display/lt101_c7 ;
  wire \u2_Display/lt101_c9 ;
  wire \u2_Display/lt102_c1 ;
  wire \u2_Display/lt102_c11 ;
  wire \u2_Display/lt102_c13 ;
  wire \u2_Display/lt102_c15 ;
  wire \u2_Display/lt102_c17 ;
  wire \u2_Display/lt102_c19 ;
  wire \u2_Display/lt102_c21 ;
  wire \u2_Display/lt102_c23 ;
  wire \u2_Display/lt102_c25 ;
  wire \u2_Display/lt102_c27 ;
  wire \u2_Display/lt102_c29 ;
  wire \u2_Display/lt102_c3 ;
  wire \u2_Display/lt102_c31 ;
  wire \u2_Display/lt102_c5 ;
  wire \u2_Display/lt102_c7 ;
  wire \u2_Display/lt102_c9 ;
  wire \u2_Display/lt103_c1 ;
  wire \u2_Display/lt103_c11 ;
  wire \u2_Display/lt103_c13 ;
  wire \u2_Display/lt103_c15 ;
  wire \u2_Display/lt103_c17 ;
  wire \u2_Display/lt103_c19 ;
  wire \u2_Display/lt103_c21 ;
  wire \u2_Display/lt103_c23 ;
  wire \u2_Display/lt103_c25 ;
  wire \u2_Display/lt103_c27 ;
  wire \u2_Display/lt103_c29 ;
  wire \u2_Display/lt103_c3 ;
  wire \u2_Display/lt103_c31 ;
  wire \u2_Display/lt103_c5 ;
  wire \u2_Display/lt103_c7 ;
  wire \u2_Display/lt103_c9 ;
  wire \u2_Display/lt104_c1 ;
  wire \u2_Display/lt104_c11 ;
  wire \u2_Display/lt104_c13 ;
  wire \u2_Display/lt104_c15 ;
  wire \u2_Display/lt104_c17 ;
  wire \u2_Display/lt104_c19 ;
  wire \u2_Display/lt104_c21 ;
  wire \u2_Display/lt104_c23 ;
  wire \u2_Display/lt104_c25 ;
  wire \u2_Display/lt104_c27 ;
  wire \u2_Display/lt104_c29 ;
  wire \u2_Display/lt104_c3 ;
  wire \u2_Display/lt104_c31 ;
  wire \u2_Display/lt104_c5 ;
  wire \u2_Display/lt104_c7 ;
  wire \u2_Display/lt104_c9 ;
  wire \u2_Display/lt105_c1 ;
  wire \u2_Display/lt105_c11 ;
  wire \u2_Display/lt105_c13 ;
  wire \u2_Display/lt105_c15 ;
  wire \u2_Display/lt105_c17 ;
  wire \u2_Display/lt105_c19 ;
  wire \u2_Display/lt105_c21 ;
  wire \u2_Display/lt105_c23 ;
  wire \u2_Display/lt105_c25 ;
  wire \u2_Display/lt105_c27 ;
  wire \u2_Display/lt105_c29 ;
  wire \u2_Display/lt105_c3 ;
  wire \u2_Display/lt105_c31 ;
  wire \u2_Display/lt105_c5 ;
  wire \u2_Display/lt105_c7 ;
  wire \u2_Display/lt105_c9 ;
  wire \u2_Display/lt106_c1 ;
  wire \u2_Display/lt106_c11 ;
  wire \u2_Display/lt106_c13 ;
  wire \u2_Display/lt106_c15 ;
  wire \u2_Display/lt106_c17 ;
  wire \u2_Display/lt106_c19 ;
  wire \u2_Display/lt106_c21 ;
  wire \u2_Display/lt106_c23 ;
  wire \u2_Display/lt106_c25 ;
  wire \u2_Display/lt106_c27 ;
  wire \u2_Display/lt106_c29 ;
  wire \u2_Display/lt106_c3 ;
  wire \u2_Display/lt106_c31 ;
  wire \u2_Display/lt106_c5 ;
  wire \u2_Display/lt106_c7 ;
  wire \u2_Display/lt106_c9 ;
  wire \u2_Display/lt107_c1 ;
  wire \u2_Display/lt107_c11 ;
  wire \u2_Display/lt107_c13 ;
  wire \u2_Display/lt107_c15 ;
  wire \u2_Display/lt107_c17 ;
  wire \u2_Display/lt107_c19 ;
  wire \u2_Display/lt107_c21 ;
  wire \u2_Display/lt107_c23 ;
  wire \u2_Display/lt107_c25 ;
  wire \u2_Display/lt107_c27 ;
  wire \u2_Display/lt107_c29 ;
  wire \u2_Display/lt107_c3 ;
  wire \u2_Display/lt107_c31 ;
  wire \u2_Display/lt107_c5 ;
  wire \u2_Display/lt107_c7 ;
  wire \u2_Display/lt107_c9 ;
  wire \u2_Display/lt108_c1 ;
  wire \u2_Display/lt108_c11 ;
  wire \u2_Display/lt108_c13 ;
  wire \u2_Display/lt108_c15 ;
  wire \u2_Display/lt108_c17 ;
  wire \u2_Display/lt108_c19 ;
  wire \u2_Display/lt108_c21 ;
  wire \u2_Display/lt108_c23 ;
  wire \u2_Display/lt108_c25 ;
  wire \u2_Display/lt108_c27 ;
  wire \u2_Display/lt108_c29 ;
  wire \u2_Display/lt108_c3 ;
  wire \u2_Display/lt108_c31 ;
  wire \u2_Display/lt108_c5 ;
  wire \u2_Display/lt108_c7 ;
  wire \u2_Display/lt108_c9 ;
  wire \u2_Display/lt109_c1 ;
  wire \u2_Display/lt109_c11 ;
  wire \u2_Display/lt109_c13 ;
  wire \u2_Display/lt109_c15 ;
  wire \u2_Display/lt109_c17 ;
  wire \u2_Display/lt109_c19 ;
  wire \u2_Display/lt109_c21 ;
  wire \u2_Display/lt109_c23 ;
  wire \u2_Display/lt109_c25 ;
  wire \u2_Display/lt109_c27 ;
  wire \u2_Display/lt109_c29 ;
  wire \u2_Display/lt109_c3 ;
  wire \u2_Display/lt109_c31 ;
  wire \u2_Display/lt109_c5 ;
  wire \u2_Display/lt109_c7 ;
  wire \u2_Display/lt109_c9 ;
  wire \u2_Display/lt10_2_c1 ;
  wire \u2_Display/lt10_2_c11 ;
  wire \u2_Display/lt10_2_c3 ;
  wire \u2_Display/lt10_2_c5 ;
  wire \u2_Display/lt10_2_c7 ;
  wire \u2_Display/lt10_2_c9 ;
  wire \u2_Display/lt110_c1 ;
  wire \u2_Display/lt110_c11 ;
  wire \u2_Display/lt110_c13 ;
  wire \u2_Display/lt110_c15 ;
  wire \u2_Display/lt110_c17 ;
  wire \u2_Display/lt110_c19 ;
  wire \u2_Display/lt110_c21 ;
  wire \u2_Display/lt110_c23 ;
  wire \u2_Display/lt110_c25 ;
  wire \u2_Display/lt110_c27 ;
  wire \u2_Display/lt110_c29 ;
  wire \u2_Display/lt110_c3 ;
  wire \u2_Display/lt110_c31 ;
  wire \u2_Display/lt110_c5 ;
  wire \u2_Display/lt110_c7 ;
  wire \u2_Display/lt110_c9 ;
  wire \u2_Display/lt11_2_c1 ;
  wire \u2_Display/lt11_2_c11 ;
  wire \u2_Display/lt11_2_c13 ;
  wire \u2_Display/lt11_2_c3 ;
  wire \u2_Display/lt11_2_c5 ;
  wire \u2_Display/lt11_2_c7 ;
  wire \u2_Display/lt11_2_c9 ;
  wire \u2_Display/lt121_c1 ;
  wire \u2_Display/lt121_c11 ;
  wire \u2_Display/lt121_c13 ;
  wire \u2_Display/lt121_c15 ;
  wire \u2_Display/lt121_c17 ;
  wire \u2_Display/lt121_c19 ;
  wire \u2_Display/lt121_c21 ;
  wire \u2_Display/lt121_c23 ;
  wire \u2_Display/lt121_c25 ;
  wire \u2_Display/lt121_c27 ;
  wire \u2_Display/lt121_c29 ;
  wire \u2_Display/lt121_c3 ;
  wire \u2_Display/lt121_c31 ;
  wire \u2_Display/lt121_c5 ;
  wire \u2_Display/lt121_c7 ;
  wire \u2_Display/lt121_c9 ;
  wire \u2_Display/lt122_c1 ;
  wire \u2_Display/lt122_c11 ;
  wire \u2_Display/lt122_c13 ;
  wire \u2_Display/lt122_c15 ;
  wire \u2_Display/lt122_c17 ;
  wire \u2_Display/lt122_c19 ;
  wire \u2_Display/lt122_c21 ;
  wire \u2_Display/lt122_c23 ;
  wire \u2_Display/lt122_c25 ;
  wire \u2_Display/lt122_c27 ;
  wire \u2_Display/lt122_c29 ;
  wire \u2_Display/lt122_c3 ;
  wire \u2_Display/lt122_c31 ;
  wire \u2_Display/lt122_c5 ;
  wire \u2_Display/lt122_c7 ;
  wire \u2_Display/lt122_c9 ;
  wire \u2_Display/lt123_c1 ;
  wire \u2_Display/lt123_c11 ;
  wire \u2_Display/lt123_c13 ;
  wire \u2_Display/lt123_c15 ;
  wire \u2_Display/lt123_c17 ;
  wire \u2_Display/lt123_c19 ;
  wire \u2_Display/lt123_c21 ;
  wire \u2_Display/lt123_c23 ;
  wire \u2_Display/lt123_c25 ;
  wire \u2_Display/lt123_c27 ;
  wire \u2_Display/lt123_c29 ;
  wire \u2_Display/lt123_c3 ;
  wire \u2_Display/lt123_c31 ;
  wire \u2_Display/lt123_c5 ;
  wire \u2_Display/lt123_c7 ;
  wire \u2_Display/lt123_c9 ;
  wire \u2_Display/lt124_c1 ;
  wire \u2_Display/lt124_c11 ;
  wire \u2_Display/lt124_c13 ;
  wire \u2_Display/lt124_c15 ;
  wire \u2_Display/lt124_c17 ;
  wire \u2_Display/lt124_c19 ;
  wire \u2_Display/lt124_c21 ;
  wire \u2_Display/lt124_c23 ;
  wire \u2_Display/lt124_c25 ;
  wire \u2_Display/lt124_c27 ;
  wire \u2_Display/lt124_c29 ;
  wire \u2_Display/lt124_c3 ;
  wire \u2_Display/lt124_c31 ;
  wire \u2_Display/lt124_c5 ;
  wire \u2_Display/lt124_c7 ;
  wire \u2_Display/lt124_c9 ;
  wire \u2_Display/lt125_c1 ;
  wire \u2_Display/lt125_c11 ;
  wire \u2_Display/lt125_c13 ;
  wire \u2_Display/lt125_c15 ;
  wire \u2_Display/lt125_c17 ;
  wire \u2_Display/lt125_c19 ;
  wire \u2_Display/lt125_c21 ;
  wire \u2_Display/lt125_c23 ;
  wire \u2_Display/lt125_c25 ;
  wire \u2_Display/lt125_c27 ;
  wire \u2_Display/lt125_c29 ;
  wire \u2_Display/lt125_c3 ;
  wire \u2_Display/lt125_c31 ;
  wire \u2_Display/lt125_c5 ;
  wire \u2_Display/lt125_c7 ;
  wire \u2_Display/lt125_c9 ;
  wire \u2_Display/lt126_c1 ;
  wire \u2_Display/lt126_c11 ;
  wire \u2_Display/lt126_c13 ;
  wire \u2_Display/lt126_c15 ;
  wire \u2_Display/lt126_c17 ;
  wire \u2_Display/lt126_c19 ;
  wire \u2_Display/lt126_c21 ;
  wire \u2_Display/lt126_c23 ;
  wire \u2_Display/lt126_c25 ;
  wire \u2_Display/lt126_c27 ;
  wire \u2_Display/lt126_c29 ;
  wire \u2_Display/lt126_c3 ;
  wire \u2_Display/lt126_c31 ;
  wire \u2_Display/lt126_c5 ;
  wire \u2_Display/lt126_c7 ;
  wire \u2_Display/lt126_c9 ;
  wire \u2_Display/lt127_c1 ;
  wire \u2_Display/lt127_c11 ;
  wire \u2_Display/lt127_c13 ;
  wire \u2_Display/lt127_c15 ;
  wire \u2_Display/lt127_c17 ;
  wire \u2_Display/lt127_c19 ;
  wire \u2_Display/lt127_c21 ;
  wire \u2_Display/lt127_c23 ;
  wire \u2_Display/lt127_c25 ;
  wire \u2_Display/lt127_c27 ;
  wire \u2_Display/lt127_c29 ;
  wire \u2_Display/lt127_c3 ;
  wire \u2_Display/lt127_c31 ;
  wire \u2_Display/lt127_c5 ;
  wire \u2_Display/lt127_c7 ;
  wire \u2_Display/lt127_c9 ;
  wire \u2_Display/lt128_c1 ;
  wire \u2_Display/lt128_c11 ;
  wire \u2_Display/lt128_c13 ;
  wire \u2_Display/lt128_c15 ;
  wire \u2_Display/lt128_c17 ;
  wire \u2_Display/lt128_c19 ;
  wire \u2_Display/lt128_c21 ;
  wire \u2_Display/lt128_c23 ;
  wire \u2_Display/lt128_c25 ;
  wire \u2_Display/lt128_c27 ;
  wire \u2_Display/lt128_c29 ;
  wire \u2_Display/lt128_c3 ;
  wire \u2_Display/lt128_c31 ;
  wire \u2_Display/lt128_c5 ;
  wire \u2_Display/lt128_c7 ;
  wire \u2_Display/lt128_c9 ;
  wire \u2_Display/lt129_c1 ;
  wire \u2_Display/lt129_c11 ;
  wire \u2_Display/lt129_c13 ;
  wire \u2_Display/lt129_c15 ;
  wire \u2_Display/lt129_c17 ;
  wire \u2_Display/lt129_c19 ;
  wire \u2_Display/lt129_c21 ;
  wire \u2_Display/lt129_c23 ;
  wire \u2_Display/lt129_c25 ;
  wire \u2_Display/lt129_c27 ;
  wire \u2_Display/lt129_c29 ;
  wire \u2_Display/lt129_c3 ;
  wire \u2_Display/lt129_c31 ;
  wire \u2_Display/lt129_c5 ;
  wire \u2_Display/lt129_c7 ;
  wire \u2_Display/lt129_c9 ;
  wire \u2_Display/lt130_c1 ;
  wire \u2_Display/lt130_c11 ;
  wire \u2_Display/lt130_c13 ;
  wire \u2_Display/lt130_c15 ;
  wire \u2_Display/lt130_c17 ;
  wire \u2_Display/lt130_c19 ;
  wire \u2_Display/lt130_c21 ;
  wire \u2_Display/lt130_c23 ;
  wire \u2_Display/lt130_c25 ;
  wire \u2_Display/lt130_c27 ;
  wire \u2_Display/lt130_c29 ;
  wire \u2_Display/lt130_c3 ;
  wire \u2_Display/lt130_c31 ;
  wire \u2_Display/lt130_c5 ;
  wire \u2_Display/lt130_c7 ;
  wire \u2_Display/lt130_c9 ;
  wire \u2_Display/lt131_c1 ;
  wire \u2_Display/lt131_c11 ;
  wire \u2_Display/lt131_c13 ;
  wire \u2_Display/lt131_c15 ;
  wire \u2_Display/lt131_c17 ;
  wire \u2_Display/lt131_c19 ;
  wire \u2_Display/lt131_c21 ;
  wire \u2_Display/lt131_c23 ;
  wire \u2_Display/lt131_c25 ;
  wire \u2_Display/lt131_c27 ;
  wire \u2_Display/lt131_c29 ;
  wire \u2_Display/lt131_c3 ;
  wire \u2_Display/lt131_c31 ;
  wire \u2_Display/lt131_c5 ;
  wire \u2_Display/lt131_c7 ;
  wire \u2_Display/lt131_c9 ;
  wire \u2_Display/lt132_c1 ;
  wire \u2_Display/lt132_c11 ;
  wire \u2_Display/lt132_c13 ;
  wire \u2_Display/lt132_c15 ;
  wire \u2_Display/lt132_c17 ;
  wire \u2_Display/lt132_c19 ;
  wire \u2_Display/lt132_c21 ;
  wire \u2_Display/lt132_c23 ;
  wire \u2_Display/lt132_c25 ;
  wire \u2_Display/lt132_c27 ;
  wire \u2_Display/lt132_c29 ;
  wire \u2_Display/lt132_c3 ;
  wire \u2_Display/lt132_c31 ;
  wire \u2_Display/lt132_c5 ;
  wire \u2_Display/lt132_c7 ;
  wire \u2_Display/lt132_c9 ;
  wire \u2_Display/lt133_c1 ;
  wire \u2_Display/lt133_c11 ;
  wire \u2_Display/lt133_c13 ;
  wire \u2_Display/lt133_c15 ;
  wire \u2_Display/lt133_c17 ;
  wire \u2_Display/lt133_c19 ;
  wire \u2_Display/lt133_c21 ;
  wire \u2_Display/lt133_c23 ;
  wire \u2_Display/lt133_c25 ;
  wire \u2_Display/lt133_c27 ;
  wire \u2_Display/lt133_c29 ;
  wire \u2_Display/lt133_c3 ;
  wire \u2_Display/lt133_c31 ;
  wire \u2_Display/lt133_c5 ;
  wire \u2_Display/lt133_c7 ;
  wire \u2_Display/lt133_c9 ;
  wire \u2_Display/lt134_c1 ;
  wire \u2_Display/lt134_c11 ;
  wire \u2_Display/lt134_c13 ;
  wire \u2_Display/lt134_c15 ;
  wire \u2_Display/lt134_c17 ;
  wire \u2_Display/lt134_c19 ;
  wire \u2_Display/lt134_c21 ;
  wire \u2_Display/lt134_c23 ;
  wire \u2_Display/lt134_c25 ;
  wire \u2_Display/lt134_c27 ;
  wire \u2_Display/lt134_c29 ;
  wire \u2_Display/lt134_c3 ;
  wire \u2_Display/lt134_c31 ;
  wire \u2_Display/lt134_c5 ;
  wire \u2_Display/lt134_c7 ;
  wire \u2_Display/lt134_c9 ;
  wire \u2_Display/lt135_c1 ;
  wire \u2_Display/lt135_c11 ;
  wire \u2_Display/lt135_c13 ;
  wire \u2_Display/lt135_c15 ;
  wire \u2_Display/lt135_c17 ;
  wire \u2_Display/lt135_c19 ;
  wire \u2_Display/lt135_c21 ;
  wire \u2_Display/lt135_c23 ;
  wire \u2_Display/lt135_c25 ;
  wire \u2_Display/lt135_c27 ;
  wire \u2_Display/lt135_c29 ;
  wire \u2_Display/lt135_c3 ;
  wire \u2_Display/lt135_c31 ;
  wire \u2_Display/lt135_c5 ;
  wire \u2_Display/lt135_c7 ;
  wire \u2_Display/lt135_c9 ;
  wire \u2_Display/lt136_c1 ;
  wire \u2_Display/lt136_c11 ;
  wire \u2_Display/lt136_c13 ;
  wire \u2_Display/lt136_c15 ;
  wire \u2_Display/lt136_c17 ;
  wire \u2_Display/lt136_c19 ;
  wire \u2_Display/lt136_c21 ;
  wire \u2_Display/lt136_c23 ;
  wire \u2_Display/lt136_c25 ;
  wire \u2_Display/lt136_c27 ;
  wire \u2_Display/lt136_c29 ;
  wire \u2_Display/lt136_c3 ;
  wire \u2_Display/lt136_c31 ;
  wire \u2_Display/lt136_c5 ;
  wire \u2_Display/lt136_c7 ;
  wire \u2_Display/lt136_c9 ;
  wire \u2_Display/lt137_c1 ;
  wire \u2_Display/lt137_c11 ;
  wire \u2_Display/lt137_c13 ;
  wire \u2_Display/lt137_c15 ;
  wire \u2_Display/lt137_c17 ;
  wire \u2_Display/lt137_c19 ;
  wire \u2_Display/lt137_c21 ;
  wire \u2_Display/lt137_c23 ;
  wire \u2_Display/lt137_c25 ;
  wire \u2_Display/lt137_c27 ;
  wire \u2_Display/lt137_c29 ;
  wire \u2_Display/lt137_c3 ;
  wire \u2_Display/lt137_c31 ;
  wire \u2_Display/lt137_c5 ;
  wire \u2_Display/lt137_c7 ;
  wire \u2_Display/lt137_c9 ;
  wire \u2_Display/lt138_c1 ;
  wire \u2_Display/lt138_c11 ;
  wire \u2_Display/lt138_c13 ;
  wire \u2_Display/lt138_c15 ;
  wire \u2_Display/lt138_c17 ;
  wire \u2_Display/lt138_c19 ;
  wire \u2_Display/lt138_c21 ;
  wire \u2_Display/lt138_c23 ;
  wire \u2_Display/lt138_c25 ;
  wire \u2_Display/lt138_c27 ;
  wire \u2_Display/lt138_c29 ;
  wire \u2_Display/lt138_c3 ;
  wire \u2_Display/lt138_c31 ;
  wire \u2_Display/lt138_c5 ;
  wire \u2_Display/lt138_c7 ;
  wire \u2_Display/lt138_c9 ;
  wire \u2_Display/lt139_c1 ;
  wire \u2_Display/lt139_c11 ;
  wire \u2_Display/lt139_c13 ;
  wire \u2_Display/lt139_c15 ;
  wire \u2_Display/lt139_c17 ;
  wire \u2_Display/lt139_c19 ;
  wire \u2_Display/lt139_c21 ;
  wire \u2_Display/lt139_c23 ;
  wire \u2_Display/lt139_c25 ;
  wire \u2_Display/lt139_c27 ;
  wire \u2_Display/lt139_c29 ;
  wire \u2_Display/lt139_c3 ;
  wire \u2_Display/lt139_c31 ;
  wire \u2_Display/lt139_c5 ;
  wire \u2_Display/lt139_c7 ;
  wire \u2_Display/lt139_c9 ;
  wire \u2_Display/lt140_c1 ;
  wire \u2_Display/lt140_c11 ;
  wire \u2_Display/lt140_c13 ;
  wire \u2_Display/lt140_c15 ;
  wire \u2_Display/lt140_c17 ;
  wire \u2_Display/lt140_c19 ;
  wire \u2_Display/lt140_c21 ;
  wire \u2_Display/lt140_c23 ;
  wire \u2_Display/lt140_c25 ;
  wire \u2_Display/lt140_c27 ;
  wire \u2_Display/lt140_c29 ;
  wire \u2_Display/lt140_c3 ;
  wire \u2_Display/lt140_c31 ;
  wire \u2_Display/lt140_c5 ;
  wire \u2_Display/lt140_c7 ;
  wire \u2_Display/lt140_c9 ;
  wire \u2_Display/lt141_c1 ;
  wire \u2_Display/lt141_c11 ;
  wire \u2_Display/lt141_c13 ;
  wire \u2_Display/lt141_c15 ;
  wire \u2_Display/lt141_c17 ;
  wire \u2_Display/lt141_c19 ;
  wire \u2_Display/lt141_c21 ;
  wire \u2_Display/lt141_c23 ;
  wire \u2_Display/lt141_c25 ;
  wire \u2_Display/lt141_c27 ;
  wire \u2_Display/lt141_c29 ;
  wire \u2_Display/lt141_c3 ;
  wire \u2_Display/lt141_c31 ;
  wire \u2_Display/lt141_c5 ;
  wire \u2_Display/lt141_c7 ;
  wire \u2_Display/lt141_c9 ;
  wire \u2_Display/lt142_c1 ;
  wire \u2_Display/lt142_c11 ;
  wire \u2_Display/lt142_c13 ;
  wire \u2_Display/lt142_c15 ;
  wire \u2_Display/lt142_c17 ;
  wire \u2_Display/lt142_c19 ;
  wire \u2_Display/lt142_c21 ;
  wire \u2_Display/lt142_c23 ;
  wire \u2_Display/lt142_c25 ;
  wire \u2_Display/lt142_c27 ;
  wire \u2_Display/lt142_c29 ;
  wire \u2_Display/lt142_c3 ;
  wire \u2_Display/lt142_c31 ;
  wire \u2_Display/lt142_c5 ;
  wire \u2_Display/lt142_c7 ;
  wire \u2_Display/lt142_c9 ;
  wire \u2_Display/lt143_c1 ;
  wire \u2_Display/lt143_c11 ;
  wire \u2_Display/lt143_c13 ;
  wire \u2_Display/lt143_c15 ;
  wire \u2_Display/lt143_c17 ;
  wire \u2_Display/lt143_c19 ;
  wire \u2_Display/lt143_c21 ;
  wire \u2_Display/lt143_c23 ;
  wire \u2_Display/lt143_c25 ;
  wire \u2_Display/lt143_c27 ;
  wire \u2_Display/lt143_c29 ;
  wire \u2_Display/lt143_c3 ;
  wire \u2_Display/lt143_c31 ;
  wire \u2_Display/lt143_c5 ;
  wire \u2_Display/lt143_c7 ;
  wire \u2_Display/lt143_c9 ;
  wire \u2_Display/lt154_c1 ;
  wire \u2_Display/lt154_c11 ;
  wire \u2_Display/lt154_c13 ;
  wire \u2_Display/lt154_c15 ;
  wire \u2_Display/lt154_c17 ;
  wire \u2_Display/lt154_c19 ;
  wire \u2_Display/lt154_c21 ;
  wire \u2_Display/lt154_c23 ;
  wire \u2_Display/lt154_c25 ;
  wire \u2_Display/lt154_c27 ;
  wire \u2_Display/lt154_c29 ;
  wire \u2_Display/lt154_c3 ;
  wire \u2_Display/lt154_c31 ;
  wire \u2_Display/lt154_c5 ;
  wire \u2_Display/lt154_c7 ;
  wire \u2_Display/lt154_c9 ;
  wire \u2_Display/lt155_c1 ;
  wire \u2_Display/lt155_c11 ;
  wire \u2_Display/lt155_c13 ;
  wire \u2_Display/lt155_c15 ;
  wire \u2_Display/lt155_c17 ;
  wire \u2_Display/lt155_c19 ;
  wire \u2_Display/lt155_c21 ;
  wire \u2_Display/lt155_c23 ;
  wire \u2_Display/lt155_c25 ;
  wire \u2_Display/lt155_c27 ;
  wire \u2_Display/lt155_c29 ;
  wire \u2_Display/lt155_c3 ;
  wire \u2_Display/lt155_c31 ;
  wire \u2_Display/lt155_c5 ;
  wire \u2_Display/lt155_c7 ;
  wire \u2_Display/lt155_c9 ;
  wire \u2_Display/lt156_c1 ;
  wire \u2_Display/lt156_c11 ;
  wire \u2_Display/lt156_c13 ;
  wire \u2_Display/lt156_c15 ;
  wire \u2_Display/lt156_c17 ;
  wire \u2_Display/lt156_c19 ;
  wire \u2_Display/lt156_c21 ;
  wire \u2_Display/lt156_c23 ;
  wire \u2_Display/lt156_c25 ;
  wire \u2_Display/lt156_c27 ;
  wire \u2_Display/lt156_c29 ;
  wire \u2_Display/lt156_c3 ;
  wire \u2_Display/lt156_c31 ;
  wire \u2_Display/lt156_c5 ;
  wire \u2_Display/lt156_c7 ;
  wire \u2_Display/lt156_c9 ;
  wire \u2_Display/lt157_c1 ;
  wire \u2_Display/lt157_c11 ;
  wire \u2_Display/lt157_c13 ;
  wire \u2_Display/lt157_c15 ;
  wire \u2_Display/lt157_c17 ;
  wire \u2_Display/lt157_c19 ;
  wire \u2_Display/lt157_c21 ;
  wire \u2_Display/lt157_c23 ;
  wire \u2_Display/lt157_c25 ;
  wire \u2_Display/lt157_c27 ;
  wire \u2_Display/lt157_c29 ;
  wire \u2_Display/lt157_c3 ;
  wire \u2_Display/lt157_c31 ;
  wire \u2_Display/lt157_c5 ;
  wire \u2_Display/lt157_c7 ;
  wire \u2_Display/lt157_c9 ;
  wire \u2_Display/lt158_c1 ;
  wire \u2_Display/lt158_c11 ;
  wire \u2_Display/lt158_c13 ;
  wire \u2_Display/lt158_c15 ;
  wire \u2_Display/lt158_c17 ;
  wire \u2_Display/lt158_c19 ;
  wire \u2_Display/lt158_c21 ;
  wire \u2_Display/lt158_c23 ;
  wire \u2_Display/lt158_c25 ;
  wire \u2_Display/lt158_c27 ;
  wire \u2_Display/lt158_c29 ;
  wire \u2_Display/lt158_c3 ;
  wire \u2_Display/lt158_c31 ;
  wire \u2_Display/lt158_c5 ;
  wire \u2_Display/lt158_c7 ;
  wire \u2_Display/lt158_c9 ;
  wire \u2_Display/lt159_c1 ;
  wire \u2_Display/lt159_c11 ;
  wire \u2_Display/lt159_c13 ;
  wire \u2_Display/lt159_c15 ;
  wire \u2_Display/lt159_c17 ;
  wire \u2_Display/lt159_c19 ;
  wire \u2_Display/lt159_c21 ;
  wire \u2_Display/lt159_c23 ;
  wire \u2_Display/lt159_c25 ;
  wire \u2_Display/lt159_c27 ;
  wire \u2_Display/lt159_c29 ;
  wire \u2_Display/lt159_c3 ;
  wire \u2_Display/lt159_c31 ;
  wire \u2_Display/lt159_c5 ;
  wire \u2_Display/lt159_c7 ;
  wire \u2_Display/lt159_c9 ;
  wire \u2_Display/lt160_c1 ;
  wire \u2_Display/lt160_c11 ;
  wire \u2_Display/lt160_c13 ;
  wire \u2_Display/lt160_c15 ;
  wire \u2_Display/lt160_c17 ;
  wire \u2_Display/lt160_c19 ;
  wire \u2_Display/lt160_c21 ;
  wire \u2_Display/lt160_c23 ;
  wire \u2_Display/lt160_c25 ;
  wire \u2_Display/lt160_c27 ;
  wire \u2_Display/lt160_c29 ;
  wire \u2_Display/lt160_c3 ;
  wire \u2_Display/lt160_c31 ;
  wire \u2_Display/lt160_c5 ;
  wire \u2_Display/lt160_c7 ;
  wire \u2_Display/lt160_c9 ;
  wire \u2_Display/lt161_c1 ;
  wire \u2_Display/lt161_c11 ;
  wire \u2_Display/lt161_c13 ;
  wire \u2_Display/lt161_c15 ;
  wire \u2_Display/lt161_c17 ;
  wire \u2_Display/lt161_c19 ;
  wire \u2_Display/lt161_c21 ;
  wire \u2_Display/lt161_c23 ;
  wire \u2_Display/lt161_c25 ;
  wire \u2_Display/lt161_c27 ;
  wire \u2_Display/lt161_c29 ;
  wire \u2_Display/lt161_c3 ;
  wire \u2_Display/lt161_c31 ;
  wire \u2_Display/lt161_c5 ;
  wire \u2_Display/lt161_c7 ;
  wire \u2_Display/lt161_c9 ;
  wire \u2_Display/lt162_c1 ;
  wire \u2_Display/lt162_c11 ;
  wire \u2_Display/lt162_c13 ;
  wire \u2_Display/lt162_c15 ;
  wire \u2_Display/lt162_c17 ;
  wire \u2_Display/lt162_c19 ;
  wire \u2_Display/lt162_c21 ;
  wire \u2_Display/lt162_c23 ;
  wire \u2_Display/lt162_c25 ;
  wire \u2_Display/lt162_c27 ;
  wire \u2_Display/lt162_c29 ;
  wire \u2_Display/lt162_c3 ;
  wire \u2_Display/lt162_c31 ;
  wire \u2_Display/lt162_c5 ;
  wire \u2_Display/lt162_c7 ;
  wire \u2_Display/lt162_c9 ;
  wire \u2_Display/lt163_c1 ;
  wire \u2_Display/lt163_c11 ;
  wire \u2_Display/lt163_c13 ;
  wire \u2_Display/lt163_c15 ;
  wire \u2_Display/lt163_c17 ;
  wire \u2_Display/lt163_c19 ;
  wire \u2_Display/lt163_c21 ;
  wire \u2_Display/lt163_c23 ;
  wire \u2_Display/lt163_c25 ;
  wire \u2_Display/lt163_c27 ;
  wire \u2_Display/lt163_c29 ;
  wire \u2_Display/lt163_c3 ;
  wire \u2_Display/lt163_c31 ;
  wire \u2_Display/lt163_c5 ;
  wire \u2_Display/lt163_c7 ;
  wire \u2_Display/lt163_c9 ;
  wire \u2_Display/lt164_c1 ;
  wire \u2_Display/lt164_c11 ;
  wire \u2_Display/lt164_c13 ;
  wire \u2_Display/lt164_c15 ;
  wire \u2_Display/lt164_c17 ;
  wire \u2_Display/lt164_c19 ;
  wire \u2_Display/lt164_c21 ;
  wire \u2_Display/lt164_c23 ;
  wire \u2_Display/lt164_c25 ;
  wire \u2_Display/lt164_c27 ;
  wire \u2_Display/lt164_c29 ;
  wire \u2_Display/lt164_c3 ;
  wire \u2_Display/lt164_c31 ;
  wire \u2_Display/lt164_c5 ;
  wire \u2_Display/lt164_c7 ;
  wire \u2_Display/lt164_c9 ;
  wire \u2_Display/lt165_c1 ;
  wire \u2_Display/lt165_c11 ;
  wire \u2_Display/lt165_c13 ;
  wire \u2_Display/lt165_c15 ;
  wire \u2_Display/lt165_c17 ;
  wire \u2_Display/lt165_c19 ;
  wire \u2_Display/lt165_c21 ;
  wire \u2_Display/lt165_c23 ;
  wire \u2_Display/lt165_c25 ;
  wire \u2_Display/lt165_c27 ;
  wire \u2_Display/lt165_c29 ;
  wire \u2_Display/lt165_c3 ;
  wire \u2_Display/lt165_c31 ;
  wire \u2_Display/lt165_c5 ;
  wire \u2_Display/lt165_c7 ;
  wire \u2_Display/lt165_c9 ;
  wire \u2_Display/lt166_c1 ;
  wire \u2_Display/lt166_c11 ;
  wire \u2_Display/lt166_c13 ;
  wire \u2_Display/lt166_c15 ;
  wire \u2_Display/lt166_c17 ;
  wire \u2_Display/lt166_c19 ;
  wire \u2_Display/lt166_c21 ;
  wire \u2_Display/lt166_c23 ;
  wire \u2_Display/lt166_c25 ;
  wire \u2_Display/lt166_c27 ;
  wire \u2_Display/lt166_c29 ;
  wire \u2_Display/lt166_c3 ;
  wire \u2_Display/lt166_c31 ;
  wire \u2_Display/lt166_c5 ;
  wire \u2_Display/lt166_c7 ;
  wire \u2_Display/lt166_c9 ;
  wire \u2_Display/lt167_c1 ;
  wire \u2_Display/lt167_c11 ;
  wire \u2_Display/lt167_c13 ;
  wire \u2_Display/lt167_c15 ;
  wire \u2_Display/lt167_c17 ;
  wire \u2_Display/lt167_c19 ;
  wire \u2_Display/lt167_c21 ;
  wire \u2_Display/lt167_c23 ;
  wire \u2_Display/lt167_c25 ;
  wire \u2_Display/lt167_c27 ;
  wire \u2_Display/lt167_c29 ;
  wire \u2_Display/lt167_c3 ;
  wire \u2_Display/lt167_c31 ;
  wire \u2_Display/lt167_c5 ;
  wire \u2_Display/lt167_c7 ;
  wire \u2_Display/lt167_c9 ;
  wire \u2_Display/lt168_c1 ;
  wire \u2_Display/lt168_c11 ;
  wire \u2_Display/lt168_c13 ;
  wire \u2_Display/lt168_c15 ;
  wire \u2_Display/lt168_c17 ;
  wire \u2_Display/lt168_c19 ;
  wire \u2_Display/lt168_c21 ;
  wire \u2_Display/lt168_c23 ;
  wire \u2_Display/lt168_c25 ;
  wire \u2_Display/lt168_c27 ;
  wire \u2_Display/lt168_c29 ;
  wire \u2_Display/lt168_c3 ;
  wire \u2_Display/lt168_c31 ;
  wire \u2_Display/lt168_c5 ;
  wire \u2_Display/lt168_c7 ;
  wire \u2_Display/lt168_c9 ;
  wire \u2_Display/lt169_c1 ;
  wire \u2_Display/lt169_c11 ;
  wire \u2_Display/lt169_c13 ;
  wire \u2_Display/lt169_c15 ;
  wire \u2_Display/lt169_c17 ;
  wire \u2_Display/lt169_c19 ;
  wire \u2_Display/lt169_c21 ;
  wire \u2_Display/lt169_c23 ;
  wire \u2_Display/lt169_c25 ;
  wire \u2_Display/lt169_c27 ;
  wire \u2_Display/lt169_c29 ;
  wire \u2_Display/lt169_c3 ;
  wire \u2_Display/lt169_c31 ;
  wire \u2_Display/lt169_c5 ;
  wire \u2_Display/lt169_c7 ;
  wire \u2_Display/lt169_c9 ;
  wire \u2_Display/lt170_c1 ;
  wire \u2_Display/lt170_c11 ;
  wire \u2_Display/lt170_c13 ;
  wire \u2_Display/lt170_c15 ;
  wire \u2_Display/lt170_c17 ;
  wire \u2_Display/lt170_c19 ;
  wire \u2_Display/lt170_c21 ;
  wire \u2_Display/lt170_c23 ;
  wire \u2_Display/lt170_c25 ;
  wire \u2_Display/lt170_c27 ;
  wire \u2_Display/lt170_c29 ;
  wire \u2_Display/lt170_c3 ;
  wire \u2_Display/lt170_c31 ;
  wire \u2_Display/lt170_c5 ;
  wire \u2_Display/lt170_c7 ;
  wire \u2_Display/lt170_c9 ;
  wire \u2_Display/lt171_c1 ;
  wire \u2_Display/lt171_c11 ;
  wire \u2_Display/lt171_c13 ;
  wire \u2_Display/lt171_c15 ;
  wire \u2_Display/lt171_c17 ;
  wire \u2_Display/lt171_c19 ;
  wire \u2_Display/lt171_c21 ;
  wire \u2_Display/lt171_c23 ;
  wire \u2_Display/lt171_c25 ;
  wire \u2_Display/lt171_c27 ;
  wire \u2_Display/lt171_c29 ;
  wire \u2_Display/lt171_c3 ;
  wire \u2_Display/lt171_c31 ;
  wire \u2_Display/lt171_c5 ;
  wire \u2_Display/lt171_c7 ;
  wire \u2_Display/lt171_c9 ;
  wire \u2_Display/lt172_c1 ;
  wire \u2_Display/lt172_c11 ;
  wire \u2_Display/lt172_c13 ;
  wire \u2_Display/lt172_c15 ;
  wire \u2_Display/lt172_c17 ;
  wire \u2_Display/lt172_c19 ;
  wire \u2_Display/lt172_c21 ;
  wire \u2_Display/lt172_c23 ;
  wire \u2_Display/lt172_c25 ;
  wire \u2_Display/lt172_c27 ;
  wire \u2_Display/lt172_c29 ;
  wire \u2_Display/lt172_c3 ;
  wire \u2_Display/lt172_c31 ;
  wire \u2_Display/lt172_c5 ;
  wire \u2_Display/lt172_c7 ;
  wire \u2_Display/lt172_c9 ;
  wire \u2_Display/lt173_c1 ;
  wire \u2_Display/lt173_c11 ;
  wire \u2_Display/lt173_c13 ;
  wire \u2_Display/lt173_c15 ;
  wire \u2_Display/lt173_c17 ;
  wire \u2_Display/lt173_c19 ;
  wire \u2_Display/lt173_c21 ;
  wire \u2_Display/lt173_c23 ;
  wire \u2_Display/lt173_c25 ;
  wire \u2_Display/lt173_c27 ;
  wire \u2_Display/lt173_c29 ;
  wire \u2_Display/lt173_c3 ;
  wire \u2_Display/lt173_c31 ;
  wire \u2_Display/lt173_c5 ;
  wire \u2_Display/lt173_c7 ;
  wire \u2_Display/lt173_c9 ;
  wire \u2_Display/lt174_c1 ;
  wire \u2_Display/lt174_c11 ;
  wire \u2_Display/lt174_c13 ;
  wire \u2_Display/lt174_c15 ;
  wire \u2_Display/lt174_c17 ;
  wire \u2_Display/lt174_c19 ;
  wire \u2_Display/lt174_c21 ;
  wire \u2_Display/lt174_c23 ;
  wire \u2_Display/lt174_c25 ;
  wire \u2_Display/lt174_c27 ;
  wire \u2_Display/lt174_c29 ;
  wire \u2_Display/lt174_c3 ;
  wire \u2_Display/lt174_c31 ;
  wire \u2_Display/lt174_c5 ;
  wire \u2_Display/lt174_c7 ;
  wire \u2_Display/lt174_c9 ;
  wire \u2_Display/lt175_c1 ;
  wire \u2_Display/lt175_c11 ;
  wire \u2_Display/lt175_c13 ;
  wire \u2_Display/lt175_c15 ;
  wire \u2_Display/lt175_c17 ;
  wire \u2_Display/lt175_c19 ;
  wire \u2_Display/lt175_c21 ;
  wire \u2_Display/lt175_c23 ;
  wire \u2_Display/lt175_c25 ;
  wire \u2_Display/lt175_c27 ;
  wire \u2_Display/lt175_c29 ;
  wire \u2_Display/lt175_c3 ;
  wire \u2_Display/lt175_c31 ;
  wire \u2_Display/lt175_c5 ;
  wire \u2_Display/lt175_c7 ;
  wire \u2_Display/lt175_c9 ;
  wire \u2_Display/lt176_c1 ;
  wire \u2_Display/lt176_c11 ;
  wire \u2_Display/lt176_c13 ;
  wire \u2_Display/lt176_c15 ;
  wire \u2_Display/lt176_c17 ;
  wire \u2_Display/lt176_c19 ;
  wire \u2_Display/lt176_c21 ;
  wire \u2_Display/lt176_c23 ;
  wire \u2_Display/lt176_c25 ;
  wire \u2_Display/lt176_c27 ;
  wire \u2_Display/lt176_c29 ;
  wire \u2_Display/lt176_c3 ;
  wire \u2_Display/lt176_c31 ;
  wire \u2_Display/lt176_c5 ;
  wire \u2_Display/lt176_c7 ;
  wire \u2_Display/lt176_c9 ;
  wire \u2_Display/lt1_c1 ;
  wire \u2_Display/lt1_c11 ;
  wire \u2_Display/lt1_c3 ;
  wire \u2_Display/lt1_c5 ;
  wire \u2_Display/lt1_c7 ;
  wire \u2_Display/lt1_c9 ;
  wire \u2_Display/lt22_c1 ;
  wire \u2_Display/lt22_c11 ;
  wire \u2_Display/lt22_c13 ;
  wire \u2_Display/lt22_c15 ;
  wire \u2_Display/lt22_c17 ;
  wire \u2_Display/lt22_c19 ;
  wire \u2_Display/lt22_c21 ;
  wire \u2_Display/lt22_c23 ;
  wire \u2_Display/lt22_c25 ;
  wire \u2_Display/lt22_c27 ;
  wire \u2_Display/lt22_c29 ;
  wire \u2_Display/lt22_c3 ;
  wire \u2_Display/lt22_c31 ;
  wire \u2_Display/lt22_c5 ;
  wire \u2_Display/lt22_c7 ;
  wire \u2_Display/lt22_c9 ;
  wire \u2_Display/lt23_c1 ;
  wire \u2_Display/lt23_c11 ;
  wire \u2_Display/lt23_c13 ;
  wire \u2_Display/lt23_c15 ;
  wire \u2_Display/lt23_c17 ;
  wire \u2_Display/lt23_c19 ;
  wire \u2_Display/lt23_c21 ;
  wire \u2_Display/lt23_c23 ;
  wire \u2_Display/lt23_c25 ;
  wire \u2_Display/lt23_c27 ;
  wire \u2_Display/lt23_c29 ;
  wire \u2_Display/lt23_c3 ;
  wire \u2_Display/lt23_c31 ;
  wire \u2_Display/lt23_c5 ;
  wire \u2_Display/lt23_c7 ;
  wire \u2_Display/lt23_c9 ;
  wire \u2_Display/lt24_c1 ;
  wire \u2_Display/lt24_c11 ;
  wire \u2_Display/lt24_c13 ;
  wire \u2_Display/lt24_c15 ;
  wire \u2_Display/lt24_c17 ;
  wire \u2_Display/lt24_c19 ;
  wire \u2_Display/lt24_c21 ;
  wire \u2_Display/lt24_c23 ;
  wire \u2_Display/lt24_c25 ;
  wire \u2_Display/lt24_c27 ;
  wire \u2_Display/lt24_c29 ;
  wire \u2_Display/lt24_c3 ;
  wire \u2_Display/lt24_c31 ;
  wire \u2_Display/lt24_c5 ;
  wire \u2_Display/lt24_c7 ;
  wire \u2_Display/lt24_c9 ;
  wire \u2_Display/lt25_c1 ;
  wire \u2_Display/lt25_c11 ;
  wire \u2_Display/lt25_c13 ;
  wire \u2_Display/lt25_c15 ;
  wire \u2_Display/lt25_c17 ;
  wire \u2_Display/lt25_c19 ;
  wire \u2_Display/lt25_c21 ;
  wire \u2_Display/lt25_c23 ;
  wire \u2_Display/lt25_c25 ;
  wire \u2_Display/lt25_c27 ;
  wire \u2_Display/lt25_c29 ;
  wire \u2_Display/lt25_c3 ;
  wire \u2_Display/lt25_c31 ;
  wire \u2_Display/lt25_c5 ;
  wire \u2_Display/lt25_c7 ;
  wire \u2_Display/lt25_c9 ;
  wire \u2_Display/lt26_c1 ;
  wire \u2_Display/lt26_c11 ;
  wire \u2_Display/lt26_c13 ;
  wire \u2_Display/lt26_c15 ;
  wire \u2_Display/lt26_c17 ;
  wire \u2_Display/lt26_c19 ;
  wire \u2_Display/lt26_c21 ;
  wire \u2_Display/lt26_c23 ;
  wire \u2_Display/lt26_c25 ;
  wire \u2_Display/lt26_c27 ;
  wire \u2_Display/lt26_c29 ;
  wire \u2_Display/lt26_c3 ;
  wire \u2_Display/lt26_c31 ;
  wire \u2_Display/lt26_c5 ;
  wire \u2_Display/lt26_c7 ;
  wire \u2_Display/lt26_c9 ;
  wire \u2_Display/lt27_c1 ;
  wire \u2_Display/lt27_c11 ;
  wire \u2_Display/lt27_c13 ;
  wire \u2_Display/lt27_c15 ;
  wire \u2_Display/lt27_c17 ;
  wire \u2_Display/lt27_c19 ;
  wire \u2_Display/lt27_c21 ;
  wire \u2_Display/lt27_c23 ;
  wire \u2_Display/lt27_c25 ;
  wire \u2_Display/lt27_c27 ;
  wire \u2_Display/lt27_c29 ;
  wire \u2_Display/lt27_c3 ;
  wire \u2_Display/lt27_c31 ;
  wire \u2_Display/lt27_c5 ;
  wire \u2_Display/lt27_c7 ;
  wire \u2_Display/lt27_c9 ;
  wire \u2_Display/lt28_c1 ;
  wire \u2_Display/lt28_c11 ;
  wire \u2_Display/lt28_c13 ;
  wire \u2_Display/lt28_c15 ;
  wire \u2_Display/lt28_c17 ;
  wire \u2_Display/lt28_c19 ;
  wire \u2_Display/lt28_c21 ;
  wire \u2_Display/lt28_c23 ;
  wire \u2_Display/lt28_c25 ;
  wire \u2_Display/lt28_c27 ;
  wire \u2_Display/lt28_c29 ;
  wire \u2_Display/lt28_c3 ;
  wire \u2_Display/lt28_c31 ;
  wire \u2_Display/lt28_c5 ;
  wire \u2_Display/lt28_c7 ;
  wire \u2_Display/lt28_c9 ;
  wire \u2_Display/lt29_c1 ;
  wire \u2_Display/lt29_c11 ;
  wire \u2_Display/lt29_c13 ;
  wire \u2_Display/lt29_c15 ;
  wire \u2_Display/lt29_c17 ;
  wire \u2_Display/lt29_c19 ;
  wire \u2_Display/lt29_c21 ;
  wire \u2_Display/lt29_c23 ;
  wire \u2_Display/lt29_c25 ;
  wire \u2_Display/lt29_c27 ;
  wire \u2_Display/lt29_c29 ;
  wire \u2_Display/lt29_c3 ;
  wire \u2_Display/lt29_c31 ;
  wire \u2_Display/lt29_c5 ;
  wire \u2_Display/lt29_c7 ;
  wire \u2_Display/lt29_c9 ;
  wire \u2_Display/lt2_2_c1 ;
  wire \u2_Display/lt2_2_c11 ;
  wire \u2_Display/lt2_2_c3 ;
  wire \u2_Display/lt2_2_c5 ;
  wire \u2_Display/lt2_2_c7 ;
  wire \u2_Display/lt2_2_c9 ;
  wire \u2_Display/lt30_c1 ;
  wire \u2_Display/lt30_c11 ;
  wire \u2_Display/lt30_c13 ;
  wire \u2_Display/lt30_c15 ;
  wire \u2_Display/lt30_c17 ;
  wire \u2_Display/lt30_c19 ;
  wire \u2_Display/lt30_c21 ;
  wire \u2_Display/lt30_c23 ;
  wire \u2_Display/lt30_c25 ;
  wire \u2_Display/lt30_c27 ;
  wire \u2_Display/lt30_c29 ;
  wire \u2_Display/lt30_c3 ;
  wire \u2_Display/lt30_c31 ;
  wire \u2_Display/lt30_c5 ;
  wire \u2_Display/lt30_c7 ;
  wire \u2_Display/lt30_c9 ;
  wire \u2_Display/lt31_c1 ;
  wire \u2_Display/lt31_c11 ;
  wire \u2_Display/lt31_c13 ;
  wire \u2_Display/lt31_c15 ;
  wire \u2_Display/lt31_c17 ;
  wire \u2_Display/lt31_c19 ;
  wire \u2_Display/lt31_c21 ;
  wire \u2_Display/lt31_c23 ;
  wire \u2_Display/lt31_c25 ;
  wire \u2_Display/lt31_c27 ;
  wire \u2_Display/lt31_c29 ;
  wire \u2_Display/lt31_c3 ;
  wire \u2_Display/lt31_c31 ;
  wire \u2_Display/lt31_c5 ;
  wire \u2_Display/lt31_c7 ;
  wire \u2_Display/lt31_c9 ;
  wire \u2_Display/lt32_c1 ;
  wire \u2_Display/lt32_c11 ;
  wire \u2_Display/lt32_c13 ;
  wire \u2_Display/lt32_c15 ;
  wire \u2_Display/lt32_c17 ;
  wire \u2_Display/lt32_c19 ;
  wire \u2_Display/lt32_c21 ;
  wire \u2_Display/lt32_c23 ;
  wire \u2_Display/lt32_c25 ;
  wire \u2_Display/lt32_c27 ;
  wire \u2_Display/lt32_c29 ;
  wire \u2_Display/lt32_c3 ;
  wire \u2_Display/lt32_c31 ;
  wire \u2_Display/lt32_c5 ;
  wire \u2_Display/lt32_c7 ;
  wire \u2_Display/lt32_c9 ;
  wire \u2_Display/lt33_c1 ;
  wire \u2_Display/lt33_c11 ;
  wire \u2_Display/lt33_c13 ;
  wire \u2_Display/lt33_c15 ;
  wire \u2_Display/lt33_c17 ;
  wire \u2_Display/lt33_c19 ;
  wire \u2_Display/lt33_c21 ;
  wire \u2_Display/lt33_c23 ;
  wire \u2_Display/lt33_c25 ;
  wire \u2_Display/lt33_c27 ;
  wire \u2_Display/lt33_c29 ;
  wire \u2_Display/lt33_c3 ;
  wire \u2_Display/lt33_c31 ;
  wire \u2_Display/lt33_c5 ;
  wire \u2_Display/lt33_c7 ;
  wire \u2_Display/lt33_c9 ;
  wire \u2_Display/lt34_c1 ;
  wire \u2_Display/lt34_c11 ;
  wire \u2_Display/lt34_c13 ;
  wire \u2_Display/lt34_c15 ;
  wire \u2_Display/lt34_c17 ;
  wire \u2_Display/lt34_c19 ;
  wire \u2_Display/lt34_c21 ;
  wire \u2_Display/lt34_c23 ;
  wire \u2_Display/lt34_c25 ;
  wire \u2_Display/lt34_c27 ;
  wire \u2_Display/lt34_c29 ;
  wire \u2_Display/lt34_c3 ;
  wire \u2_Display/lt34_c31 ;
  wire \u2_Display/lt34_c5 ;
  wire \u2_Display/lt34_c7 ;
  wire \u2_Display/lt34_c9 ;
  wire \u2_Display/lt35_c1 ;
  wire \u2_Display/lt35_c11 ;
  wire \u2_Display/lt35_c13 ;
  wire \u2_Display/lt35_c15 ;
  wire \u2_Display/lt35_c17 ;
  wire \u2_Display/lt35_c19 ;
  wire \u2_Display/lt35_c21 ;
  wire \u2_Display/lt35_c23 ;
  wire \u2_Display/lt35_c25 ;
  wire \u2_Display/lt35_c27 ;
  wire \u2_Display/lt35_c29 ;
  wire \u2_Display/lt35_c3 ;
  wire \u2_Display/lt35_c31 ;
  wire \u2_Display/lt35_c5 ;
  wire \u2_Display/lt35_c7 ;
  wire \u2_Display/lt35_c9 ;
  wire \u2_Display/lt36_c1 ;
  wire \u2_Display/lt36_c11 ;
  wire \u2_Display/lt36_c13 ;
  wire \u2_Display/lt36_c15 ;
  wire \u2_Display/lt36_c17 ;
  wire \u2_Display/lt36_c19 ;
  wire \u2_Display/lt36_c21 ;
  wire \u2_Display/lt36_c23 ;
  wire \u2_Display/lt36_c25 ;
  wire \u2_Display/lt36_c27 ;
  wire \u2_Display/lt36_c29 ;
  wire \u2_Display/lt36_c3 ;
  wire \u2_Display/lt36_c31 ;
  wire \u2_Display/lt36_c5 ;
  wire \u2_Display/lt36_c7 ;
  wire \u2_Display/lt36_c9 ;
  wire \u2_Display/lt37_c1 ;
  wire \u2_Display/lt37_c11 ;
  wire \u2_Display/lt37_c13 ;
  wire \u2_Display/lt37_c15 ;
  wire \u2_Display/lt37_c17 ;
  wire \u2_Display/lt37_c19 ;
  wire \u2_Display/lt37_c21 ;
  wire \u2_Display/lt37_c23 ;
  wire \u2_Display/lt37_c25 ;
  wire \u2_Display/lt37_c27 ;
  wire \u2_Display/lt37_c29 ;
  wire \u2_Display/lt37_c3 ;
  wire \u2_Display/lt37_c31 ;
  wire \u2_Display/lt37_c5 ;
  wire \u2_Display/lt37_c7 ;
  wire \u2_Display/lt37_c9 ;
  wire \u2_Display/lt38_c1 ;
  wire \u2_Display/lt38_c11 ;
  wire \u2_Display/lt38_c13 ;
  wire \u2_Display/lt38_c15 ;
  wire \u2_Display/lt38_c17 ;
  wire \u2_Display/lt38_c19 ;
  wire \u2_Display/lt38_c21 ;
  wire \u2_Display/lt38_c23 ;
  wire \u2_Display/lt38_c25 ;
  wire \u2_Display/lt38_c27 ;
  wire \u2_Display/lt38_c29 ;
  wire \u2_Display/lt38_c3 ;
  wire \u2_Display/lt38_c31 ;
  wire \u2_Display/lt38_c5 ;
  wire \u2_Display/lt38_c7 ;
  wire \u2_Display/lt38_c9 ;
  wire \u2_Display/lt39_c1 ;
  wire \u2_Display/lt39_c11 ;
  wire \u2_Display/lt39_c13 ;
  wire \u2_Display/lt39_c15 ;
  wire \u2_Display/lt39_c17 ;
  wire \u2_Display/lt39_c19 ;
  wire \u2_Display/lt39_c21 ;
  wire \u2_Display/lt39_c23 ;
  wire \u2_Display/lt39_c25 ;
  wire \u2_Display/lt39_c27 ;
  wire \u2_Display/lt39_c29 ;
  wire \u2_Display/lt39_c3 ;
  wire \u2_Display/lt39_c31 ;
  wire \u2_Display/lt39_c5 ;
  wire \u2_Display/lt39_c7 ;
  wire \u2_Display/lt39_c9 ;
  wire \u2_Display/lt3_c1 ;
  wire \u2_Display/lt3_c11 ;
  wire \u2_Display/lt3_c3 ;
  wire \u2_Display/lt3_c5 ;
  wire \u2_Display/lt3_c7 ;
  wire \u2_Display/lt3_c9 ;
  wire \u2_Display/lt40_c1 ;
  wire \u2_Display/lt40_c11 ;
  wire \u2_Display/lt40_c13 ;
  wire \u2_Display/lt40_c15 ;
  wire \u2_Display/lt40_c17 ;
  wire \u2_Display/lt40_c19 ;
  wire \u2_Display/lt40_c21 ;
  wire \u2_Display/lt40_c23 ;
  wire \u2_Display/lt40_c25 ;
  wire \u2_Display/lt40_c27 ;
  wire \u2_Display/lt40_c29 ;
  wire \u2_Display/lt40_c3 ;
  wire \u2_Display/lt40_c31 ;
  wire \u2_Display/lt40_c5 ;
  wire \u2_Display/lt40_c7 ;
  wire \u2_Display/lt40_c9 ;
  wire \u2_Display/lt41_c1 ;
  wire \u2_Display/lt41_c11 ;
  wire \u2_Display/lt41_c13 ;
  wire \u2_Display/lt41_c15 ;
  wire \u2_Display/lt41_c17 ;
  wire \u2_Display/lt41_c19 ;
  wire \u2_Display/lt41_c21 ;
  wire \u2_Display/lt41_c23 ;
  wire \u2_Display/lt41_c25 ;
  wire \u2_Display/lt41_c27 ;
  wire \u2_Display/lt41_c29 ;
  wire \u2_Display/lt41_c3 ;
  wire \u2_Display/lt41_c31 ;
  wire \u2_Display/lt41_c5 ;
  wire \u2_Display/lt41_c7 ;
  wire \u2_Display/lt41_c9 ;
  wire \u2_Display/lt42_c1 ;
  wire \u2_Display/lt42_c11 ;
  wire \u2_Display/lt42_c13 ;
  wire \u2_Display/lt42_c15 ;
  wire \u2_Display/lt42_c17 ;
  wire \u2_Display/lt42_c19 ;
  wire \u2_Display/lt42_c21 ;
  wire \u2_Display/lt42_c23 ;
  wire \u2_Display/lt42_c25 ;
  wire \u2_Display/lt42_c27 ;
  wire \u2_Display/lt42_c29 ;
  wire \u2_Display/lt42_c3 ;
  wire \u2_Display/lt42_c31 ;
  wire \u2_Display/lt42_c5 ;
  wire \u2_Display/lt42_c7 ;
  wire \u2_Display/lt42_c9 ;
  wire \u2_Display/lt43_c1 ;
  wire \u2_Display/lt43_c11 ;
  wire \u2_Display/lt43_c13 ;
  wire \u2_Display/lt43_c15 ;
  wire \u2_Display/lt43_c17 ;
  wire \u2_Display/lt43_c19 ;
  wire \u2_Display/lt43_c21 ;
  wire \u2_Display/lt43_c23 ;
  wire \u2_Display/lt43_c25 ;
  wire \u2_Display/lt43_c27 ;
  wire \u2_Display/lt43_c29 ;
  wire \u2_Display/lt43_c3 ;
  wire \u2_Display/lt43_c31 ;
  wire \u2_Display/lt43_c5 ;
  wire \u2_Display/lt43_c7 ;
  wire \u2_Display/lt43_c9 ;
  wire \u2_Display/lt44_c1 ;
  wire \u2_Display/lt44_c11 ;
  wire \u2_Display/lt44_c13 ;
  wire \u2_Display/lt44_c15 ;
  wire \u2_Display/lt44_c17 ;
  wire \u2_Display/lt44_c19 ;
  wire \u2_Display/lt44_c21 ;
  wire \u2_Display/lt44_c23 ;
  wire \u2_Display/lt44_c25 ;
  wire \u2_Display/lt44_c27 ;
  wire \u2_Display/lt44_c29 ;
  wire \u2_Display/lt44_c3 ;
  wire \u2_Display/lt44_c31 ;
  wire \u2_Display/lt44_c5 ;
  wire \u2_Display/lt44_c7 ;
  wire \u2_Display/lt44_c9 ;
  wire \u2_Display/lt4_2_c1 ;
  wire \u2_Display/lt4_2_c11 ;
  wire \u2_Display/lt4_2_c3 ;
  wire \u2_Display/lt4_2_c5 ;
  wire \u2_Display/lt4_2_c7 ;
  wire \u2_Display/lt4_2_c9 ;
  wire \u2_Display/lt55_c1 ;
  wire \u2_Display/lt55_c11 ;
  wire \u2_Display/lt55_c13 ;
  wire \u2_Display/lt55_c15 ;
  wire \u2_Display/lt55_c17 ;
  wire \u2_Display/lt55_c19 ;
  wire \u2_Display/lt55_c21 ;
  wire \u2_Display/lt55_c23 ;
  wire \u2_Display/lt55_c25 ;
  wire \u2_Display/lt55_c27 ;
  wire \u2_Display/lt55_c29 ;
  wire \u2_Display/lt55_c3 ;
  wire \u2_Display/lt55_c31 ;
  wire \u2_Display/lt55_c5 ;
  wire \u2_Display/lt55_c7 ;
  wire \u2_Display/lt55_c9 ;
  wire \u2_Display/lt56_c1 ;
  wire \u2_Display/lt56_c11 ;
  wire \u2_Display/lt56_c13 ;
  wire \u2_Display/lt56_c15 ;
  wire \u2_Display/lt56_c17 ;
  wire \u2_Display/lt56_c19 ;
  wire \u2_Display/lt56_c21 ;
  wire \u2_Display/lt56_c23 ;
  wire \u2_Display/lt56_c25 ;
  wire \u2_Display/lt56_c27 ;
  wire \u2_Display/lt56_c29 ;
  wire \u2_Display/lt56_c3 ;
  wire \u2_Display/lt56_c31 ;
  wire \u2_Display/lt56_c5 ;
  wire \u2_Display/lt56_c7 ;
  wire \u2_Display/lt56_c9 ;
  wire \u2_Display/lt57_c1 ;
  wire \u2_Display/lt57_c11 ;
  wire \u2_Display/lt57_c13 ;
  wire \u2_Display/lt57_c15 ;
  wire \u2_Display/lt57_c17 ;
  wire \u2_Display/lt57_c19 ;
  wire \u2_Display/lt57_c21 ;
  wire \u2_Display/lt57_c23 ;
  wire \u2_Display/lt57_c25 ;
  wire \u2_Display/lt57_c27 ;
  wire \u2_Display/lt57_c29 ;
  wire \u2_Display/lt57_c3 ;
  wire \u2_Display/lt57_c31 ;
  wire \u2_Display/lt57_c5 ;
  wire \u2_Display/lt57_c7 ;
  wire \u2_Display/lt57_c9 ;
  wire \u2_Display/lt58_c1 ;
  wire \u2_Display/lt58_c11 ;
  wire \u2_Display/lt58_c13 ;
  wire \u2_Display/lt58_c15 ;
  wire \u2_Display/lt58_c17 ;
  wire \u2_Display/lt58_c19 ;
  wire \u2_Display/lt58_c21 ;
  wire \u2_Display/lt58_c23 ;
  wire \u2_Display/lt58_c25 ;
  wire \u2_Display/lt58_c27 ;
  wire \u2_Display/lt58_c29 ;
  wire \u2_Display/lt58_c3 ;
  wire \u2_Display/lt58_c31 ;
  wire \u2_Display/lt58_c5 ;
  wire \u2_Display/lt58_c7 ;
  wire \u2_Display/lt58_c9 ;
  wire \u2_Display/lt59_c1 ;
  wire \u2_Display/lt59_c11 ;
  wire \u2_Display/lt59_c13 ;
  wire \u2_Display/lt59_c15 ;
  wire \u2_Display/lt59_c17 ;
  wire \u2_Display/lt59_c19 ;
  wire \u2_Display/lt59_c21 ;
  wire \u2_Display/lt59_c23 ;
  wire \u2_Display/lt59_c25 ;
  wire \u2_Display/lt59_c27 ;
  wire \u2_Display/lt59_c29 ;
  wire \u2_Display/lt59_c3 ;
  wire \u2_Display/lt59_c31 ;
  wire \u2_Display/lt59_c5 ;
  wire \u2_Display/lt59_c7 ;
  wire \u2_Display/lt59_c9 ;
  wire \u2_Display/lt5_2_c1 ;
  wire \u2_Display/lt5_2_c11 ;
  wire \u2_Display/lt5_2_c13 ;
  wire \u2_Display/lt5_2_c3 ;
  wire \u2_Display/lt5_2_c5 ;
  wire \u2_Display/lt5_2_c7 ;
  wire \u2_Display/lt5_2_c9 ;
  wire \u2_Display/lt60_c1 ;
  wire \u2_Display/lt60_c11 ;
  wire \u2_Display/lt60_c13 ;
  wire \u2_Display/lt60_c15 ;
  wire \u2_Display/lt60_c17 ;
  wire \u2_Display/lt60_c19 ;
  wire \u2_Display/lt60_c21 ;
  wire \u2_Display/lt60_c23 ;
  wire \u2_Display/lt60_c25 ;
  wire \u2_Display/lt60_c27 ;
  wire \u2_Display/lt60_c29 ;
  wire \u2_Display/lt60_c3 ;
  wire \u2_Display/lt60_c31 ;
  wire \u2_Display/lt60_c5 ;
  wire \u2_Display/lt60_c7 ;
  wire \u2_Display/lt60_c9 ;
  wire \u2_Display/lt61_c1 ;
  wire \u2_Display/lt61_c11 ;
  wire \u2_Display/lt61_c13 ;
  wire \u2_Display/lt61_c15 ;
  wire \u2_Display/lt61_c17 ;
  wire \u2_Display/lt61_c19 ;
  wire \u2_Display/lt61_c21 ;
  wire \u2_Display/lt61_c23 ;
  wire \u2_Display/lt61_c25 ;
  wire \u2_Display/lt61_c27 ;
  wire \u2_Display/lt61_c29 ;
  wire \u2_Display/lt61_c3 ;
  wire \u2_Display/lt61_c31 ;
  wire \u2_Display/lt61_c5 ;
  wire \u2_Display/lt61_c7 ;
  wire \u2_Display/lt61_c9 ;
  wire \u2_Display/lt62_c1 ;
  wire \u2_Display/lt62_c11 ;
  wire \u2_Display/lt62_c13 ;
  wire \u2_Display/lt62_c15 ;
  wire \u2_Display/lt62_c17 ;
  wire \u2_Display/lt62_c19 ;
  wire \u2_Display/lt62_c21 ;
  wire \u2_Display/lt62_c23 ;
  wire \u2_Display/lt62_c25 ;
  wire \u2_Display/lt62_c27 ;
  wire \u2_Display/lt62_c29 ;
  wire \u2_Display/lt62_c3 ;
  wire \u2_Display/lt62_c31 ;
  wire \u2_Display/lt62_c5 ;
  wire \u2_Display/lt62_c7 ;
  wire \u2_Display/lt62_c9 ;
  wire \u2_Display/lt63_c1 ;
  wire \u2_Display/lt63_c11 ;
  wire \u2_Display/lt63_c13 ;
  wire \u2_Display/lt63_c15 ;
  wire \u2_Display/lt63_c17 ;
  wire \u2_Display/lt63_c19 ;
  wire \u2_Display/lt63_c21 ;
  wire \u2_Display/lt63_c23 ;
  wire \u2_Display/lt63_c25 ;
  wire \u2_Display/lt63_c27 ;
  wire \u2_Display/lt63_c29 ;
  wire \u2_Display/lt63_c3 ;
  wire \u2_Display/lt63_c31 ;
  wire \u2_Display/lt63_c5 ;
  wire \u2_Display/lt63_c7 ;
  wire \u2_Display/lt63_c9 ;
  wire \u2_Display/lt64_c1 ;
  wire \u2_Display/lt64_c11 ;
  wire \u2_Display/lt64_c13 ;
  wire \u2_Display/lt64_c15 ;
  wire \u2_Display/lt64_c17 ;
  wire \u2_Display/lt64_c19 ;
  wire \u2_Display/lt64_c21 ;
  wire \u2_Display/lt64_c23 ;
  wire \u2_Display/lt64_c25 ;
  wire \u2_Display/lt64_c27 ;
  wire \u2_Display/lt64_c29 ;
  wire \u2_Display/lt64_c3 ;
  wire \u2_Display/lt64_c31 ;
  wire \u2_Display/lt64_c5 ;
  wire \u2_Display/lt64_c7 ;
  wire \u2_Display/lt64_c9 ;
  wire \u2_Display/lt65_c1 ;
  wire \u2_Display/lt65_c11 ;
  wire \u2_Display/lt65_c13 ;
  wire \u2_Display/lt65_c15 ;
  wire \u2_Display/lt65_c17 ;
  wire \u2_Display/lt65_c19 ;
  wire \u2_Display/lt65_c21 ;
  wire \u2_Display/lt65_c23 ;
  wire \u2_Display/lt65_c25 ;
  wire \u2_Display/lt65_c27 ;
  wire \u2_Display/lt65_c29 ;
  wire \u2_Display/lt65_c3 ;
  wire \u2_Display/lt65_c31 ;
  wire \u2_Display/lt65_c5 ;
  wire \u2_Display/lt65_c7 ;
  wire \u2_Display/lt65_c9 ;
  wire \u2_Display/lt66_c1 ;
  wire \u2_Display/lt66_c11 ;
  wire \u2_Display/lt66_c13 ;
  wire \u2_Display/lt66_c15 ;
  wire \u2_Display/lt66_c17 ;
  wire \u2_Display/lt66_c19 ;
  wire \u2_Display/lt66_c21 ;
  wire \u2_Display/lt66_c23 ;
  wire \u2_Display/lt66_c25 ;
  wire \u2_Display/lt66_c27 ;
  wire \u2_Display/lt66_c29 ;
  wire \u2_Display/lt66_c3 ;
  wire \u2_Display/lt66_c31 ;
  wire \u2_Display/lt66_c5 ;
  wire \u2_Display/lt66_c7 ;
  wire \u2_Display/lt66_c9 ;
  wire \u2_Display/lt67_c1 ;
  wire \u2_Display/lt67_c11 ;
  wire \u2_Display/lt67_c13 ;
  wire \u2_Display/lt67_c15 ;
  wire \u2_Display/lt67_c17 ;
  wire \u2_Display/lt67_c19 ;
  wire \u2_Display/lt67_c21 ;
  wire \u2_Display/lt67_c23 ;
  wire \u2_Display/lt67_c25 ;
  wire \u2_Display/lt67_c27 ;
  wire \u2_Display/lt67_c29 ;
  wire \u2_Display/lt67_c3 ;
  wire \u2_Display/lt67_c31 ;
  wire \u2_Display/lt67_c5 ;
  wire \u2_Display/lt67_c7 ;
  wire \u2_Display/lt67_c9 ;
  wire \u2_Display/lt68_c1 ;
  wire \u2_Display/lt68_c11 ;
  wire \u2_Display/lt68_c13 ;
  wire \u2_Display/lt68_c15 ;
  wire \u2_Display/lt68_c17 ;
  wire \u2_Display/lt68_c19 ;
  wire \u2_Display/lt68_c21 ;
  wire \u2_Display/lt68_c23 ;
  wire \u2_Display/lt68_c25 ;
  wire \u2_Display/lt68_c27 ;
  wire \u2_Display/lt68_c29 ;
  wire \u2_Display/lt68_c3 ;
  wire \u2_Display/lt68_c31 ;
  wire \u2_Display/lt68_c5 ;
  wire \u2_Display/lt68_c7 ;
  wire \u2_Display/lt68_c9 ;
  wire \u2_Display/lt69_c1 ;
  wire \u2_Display/lt69_c11 ;
  wire \u2_Display/lt69_c13 ;
  wire \u2_Display/lt69_c15 ;
  wire \u2_Display/lt69_c17 ;
  wire \u2_Display/lt69_c19 ;
  wire \u2_Display/lt69_c21 ;
  wire \u2_Display/lt69_c23 ;
  wire \u2_Display/lt69_c25 ;
  wire \u2_Display/lt69_c27 ;
  wire \u2_Display/lt69_c29 ;
  wire \u2_Display/lt69_c3 ;
  wire \u2_Display/lt69_c31 ;
  wire \u2_Display/lt69_c5 ;
  wire \u2_Display/lt69_c7 ;
  wire \u2_Display/lt69_c9 ;
  wire \u2_Display/lt6_2_c1 ;
  wire \u2_Display/lt6_2_c11 ;
  wire \u2_Display/lt6_2_c3 ;
  wire \u2_Display/lt6_2_c5 ;
  wire \u2_Display/lt6_2_c7 ;
  wire \u2_Display/lt6_2_c9 ;
  wire \u2_Display/lt70_c1 ;
  wire \u2_Display/lt70_c11 ;
  wire \u2_Display/lt70_c13 ;
  wire \u2_Display/lt70_c15 ;
  wire \u2_Display/lt70_c17 ;
  wire \u2_Display/lt70_c19 ;
  wire \u2_Display/lt70_c21 ;
  wire \u2_Display/lt70_c23 ;
  wire \u2_Display/lt70_c25 ;
  wire \u2_Display/lt70_c27 ;
  wire \u2_Display/lt70_c29 ;
  wire \u2_Display/lt70_c3 ;
  wire \u2_Display/lt70_c31 ;
  wire \u2_Display/lt70_c5 ;
  wire \u2_Display/lt70_c7 ;
  wire \u2_Display/lt70_c9 ;
  wire \u2_Display/lt71_c1 ;
  wire \u2_Display/lt71_c11 ;
  wire \u2_Display/lt71_c13 ;
  wire \u2_Display/lt71_c15 ;
  wire \u2_Display/lt71_c17 ;
  wire \u2_Display/lt71_c19 ;
  wire \u2_Display/lt71_c21 ;
  wire \u2_Display/lt71_c23 ;
  wire \u2_Display/lt71_c25 ;
  wire \u2_Display/lt71_c27 ;
  wire \u2_Display/lt71_c29 ;
  wire \u2_Display/lt71_c3 ;
  wire \u2_Display/lt71_c31 ;
  wire \u2_Display/lt71_c5 ;
  wire \u2_Display/lt71_c7 ;
  wire \u2_Display/lt71_c9 ;
  wire \u2_Display/lt72_c1 ;
  wire \u2_Display/lt72_c11 ;
  wire \u2_Display/lt72_c13 ;
  wire \u2_Display/lt72_c15 ;
  wire \u2_Display/lt72_c17 ;
  wire \u2_Display/lt72_c19 ;
  wire \u2_Display/lt72_c21 ;
  wire \u2_Display/lt72_c23 ;
  wire \u2_Display/lt72_c25 ;
  wire \u2_Display/lt72_c27 ;
  wire \u2_Display/lt72_c29 ;
  wire \u2_Display/lt72_c3 ;
  wire \u2_Display/lt72_c31 ;
  wire \u2_Display/lt72_c5 ;
  wire \u2_Display/lt72_c7 ;
  wire \u2_Display/lt72_c9 ;
  wire \u2_Display/lt73_c1 ;
  wire \u2_Display/lt73_c11 ;
  wire \u2_Display/lt73_c13 ;
  wire \u2_Display/lt73_c15 ;
  wire \u2_Display/lt73_c17 ;
  wire \u2_Display/lt73_c19 ;
  wire \u2_Display/lt73_c21 ;
  wire \u2_Display/lt73_c23 ;
  wire \u2_Display/lt73_c25 ;
  wire \u2_Display/lt73_c27 ;
  wire \u2_Display/lt73_c29 ;
  wire \u2_Display/lt73_c3 ;
  wire \u2_Display/lt73_c31 ;
  wire \u2_Display/lt73_c5 ;
  wire \u2_Display/lt73_c7 ;
  wire \u2_Display/lt73_c9 ;
  wire \u2_Display/lt74_c1 ;
  wire \u2_Display/lt74_c11 ;
  wire \u2_Display/lt74_c13 ;
  wire \u2_Display/lt74_c15 ;
  wire \u2_Display/lt74_c17 ;
  wire \u2_Display/lt74_c19 ;
  wire \u2_Display/lt74_c21 ;
  wire \u2_Display/lt74_c23 ;
  wire \u2_Display/lt74_c25 ;
  wire \u2_Display/lt74_c27 ;
  wire \u2_Display/lt74_c29 ;
  wire \u2_Display/lt74_c3 ;
  wire \u2_Display/lt74_c31 ;
  wire \u2_Display/lt74_c5 ;
  wire \u2_Display/lt74_c7 ;
  wire \u2_Display/lt74_c9 ;
  wire \u2_Display/lt75_c1 ;
  wire \u2_Display/lt75_c11 ;
  wire \u2_Display/lt75_c13 ;
  wire \u2_Display/lt75_c15 ;
  wire \u2_Display/lt75_c17 ;
  wire \u2_Display/lt75_c19 ;
  wire \u2_Display/lt75_c21 ;
  wire \u2_Display/lt75_c23 ;
  wire \u2_Display/lt75_c25 ;
  wire \u2_Display/lt75_c27 ;
  wire \u2_Display/lt75_c29 ;
  wire \u2_Display/lt75_c3 ;
  wire \u2_Display/lt75_c31 ;
  wire \u2_Display/lt75_c5 ;
  wire \u2_Display/lt75_c7 ;
  wire \u2_Display/lt75_c9 ;
  wire \u2_Display/lt76_c1 ;
  wire \u2_Display/lt76_c11 ;
  wire \u2_Display/lt76_c13 ;
  wire \u2_Display/lt76_c15 ;
  wire \u2_Display/lt76_c17 ;
  wire \u2_Display/lt76_c19 ;
  wire \u2_Display/lt76_c21 ;
  wire \u2_Display/lt76_c23 ;
  wire \u2_Display/lt76_c25 ;
  wire \u2_Display/lt76_c27 ;
  wire \u2_Display/lt76_c29 ;
  wire \u2_Display/lt76_c3 ;
  wire \u2_Display/lt76_c31 ;
  wire \u2_Display/lt76_c5 ;
  wire \u2_Display/lt76_c7 ;
  wire \u2_Display/lt76_c9 ;
  wire \u2_Display/lt77_c1 ;
  wire \u2_Display/lt77_c11 ;
  wire \u2_Display/lt77_c13 ;
  wire \u2_Display/lt77_c15 ;
  wire \u2_Display/lt77_c17 ;
  wire \u2_Display/lt77_c19 ;
  wire \u2_Display/lt77_c21 ;
  wire \u2_Display/lt77_c23 ;
  wire \u2_Display/lt77_c25 ;
  wire \u2_Display/lt77_c27 ;
  wire \u2_Display/lt77_c29 ;
  wire \u2_Display/lt77_c3 ;
  wire \u2_Display/lt77_c31 ;
  wire \u2_Display/lt77_c5 ;
  wire \u2_Display/lt77_c7 ;
  wire \u2_Display/lt77_c9 ;
  wire \u2_Display/lt7_2_c1 ;
  wire \u2_Display/lt7_2_c11 ;
  wire \u2_Display/lt7_2_c13 ;
  wire \u2_Display/lt7_2_c3 ;
  wire \u2_Display/lt7_2_c5 ;
  wire \u2_Display/lt7_2_c7 ;
  wire \u2_Display/lt7_2_c9 ;
  wire \u2_Display/lt88_c1 ;
  wire \u2_Display/lt88_c11 ;
  wire \u2_Display/lt88_c13 ;
  wire \u2_Display/lt88_c15 ;
  wire \u2_Display/lt88_c17 ;
  wire \u2_Display/lt88_c19 ;
  wire \u2_Display/lt88_c21 ;
  wire \u2_Display/lt88_c23 ;
  wire \u2_Display/lt88_c25 ;
  wire \u2_Display/lt88_c27 ;
  wire \u2_Display/lt88_c29 ;
  wire \u2_Display/lt88_c3 ;
  wire \u2_Display/lt88_c31 ;
  wire \u2_Display/lt88_c5 ;
  wire \u2_Display/lt88_c7 ;
  wire \u2_Display/lt88_c9 ;
  wire \u2_Display/lt89_c1 ;
  wire \u2_Display/lt89_c11 ;
  wire \u2_Display/lt89_c13 ;
  wire \u2_Display/lt89_c15 ;
  wire \u2_Display/lt89_c17 ;
  wire \u2_Display/lt89_c19 ;
  wire \u2_Display/lt89_c21 ;
  wire \u2_Display/lt89_c23 ;
  wire \u2_Display/lt89_c25 ;
  wire \u2_Display/lt89_c27 ;
  wire \u2_Display/lt89_c29 ;
  wire \u2_Display/lt89_c3 ;
  wire \u2_Display/lt89_c31 ;
  wire \u2_Display/lt89_c5 ;
  wire \u2_Display/lt89_c7 ;
  wire \u2_Display/lt89_c9 ;
  wire \u2_Display/lt8_2_c1 ;
  wire \u2_Display/lt8_2_c11 ;
  wire \u2_Display/lt8_2_c3 ;
  wire \u2_Display/lt8_2_c5 ;
  wire \u2_Display/lt8_2_c7 ;
  wire \u2_Display/lt8_2_c9 ;
  wire \u2_Display/lt90_c1 ;
  wire \u2_Display/lt90_c11 ;
  wire \u2_Display/lt90_c13 ;
  wire \u2_Display/lt90_c15 ;
  wire \u2_Display/lt90_c17 ;
  wire \u2_Display/lt90_c19 ;
  wire \u2_Display/lt90_c21 ;
  wire \u2_Display/lt90_c23 ;
  wire \u2_Display/lt90_c25 ;
  wire \u2_Display/lt90_c27 ;
  wire \u2_Display/lt90_c29 ;
  wire \u2_Display/lt90_c3 ;
  wire \u2_Display/lt90_c31 ;
  wire \u2_Display/lt90_c5 ;
  wire \u2_Display/lt90_c7 ;
  wire \u2_Display/lt90_c9 ;
  wire \u2_Display/lt91_c1 ;
  wire \u2_Display/lt91_c11 ;
  wire \u2_Display/lt91_c13 ;
  wire \u2_Display/lt91_c15 ;
  wire \u2_Display/lt91_c17 ;
  wire \u2_Display/lt91_c19 ;
  wire \u2_Display/lt91_c21 ;
  wire \u2_Display/lt91_c23 ;
  wire \u2_Display/lt91_c25 ;
  wire \u2_Display/lt91_c27 ;
  wire \u2_Display/lt91_c29 ;
  wire \u2_Display/lt91_c3 ;
  wire \u2_Display/lt91_c31 ;
  wire \u2_Display/lt91_c5 ;
  wire \u2_Display/lt91_c7 ;
  wire \u2_Display/lt91_c9 ;
  wire \u2_Display/lt92_c1 ;
  wire \u2_Display/lt92_c11 ;
  wire \u2_Display/lt92_c13 ;
  wire \u2_Display/lt92_c15 ;
  wire \u2_Display/lt92_c17 ;
  wire \u2_Display/lt92_c19 ;
  wire \u2_Display/lt92_c21 ;
  wire \u2_Display/lt92_c23 ;
  wire \u2_Display/lt92_c25 ;
  wire \u2_Display/lt92_c27 ;
  wire \u2_Display/lt92_c29 ;
  wire \u2_Display/lt92_c3 ;
  wire \u2_Display/lt92_c31 ;
  wire \u2_Display/lt92_c5 ;
  wire \u2_Display/lt92_c7 ;
  wire \u2_Display/lt92_c9 ;
  wire \u2_Display/lt93_c1 ;
  wire \u2_Display/lt93_c11 ;
  wire \u2_Display/lt93_c13 ;
  wire \u2_Display/lt93_c15 ;
  wire \u2_Display/lt93_c17 ;
  wire \u2_Display/lt93_c19 ;
  wire \u2_Display/lt93_c21 ;
  wire \u2_Display/lt93_c23 ;
  wire \u2_Display/lt93_c25 ;
  wire \u2_Display/lt93_c27 ;
  wire \u2_Display/lt93_c29 ;
  wire \u2_Display/lt93_c3 ;
  wire \u2_Display/lt93_c31 ;
  wire \u2_Display/lt93_c5 ;
  wire \u2_Display/lt93_c7 ;
  wire \u2_Display/lt93_c9 ;
  wire \u2_Display/lt94_c1 ;
  wire \u2_Display/lt94_c11 ;
  wire \u2_Display/lt94_c13 ;
  wire \u2_Display/lt94_c15 ;
  wire \u2_Display/lt94_c17 ;
  wire \u2_Display/lt94_c19 ;
  wire \u2_Display/lt94_c21 ;
  wire \u2_Display/lt94_c23 ;
  wire \u2_Display/lt94_c25 ;
  wire \u2_Display/lt94_c27 ;
  wire \u2_Display/lt94_c29 ;
  wire \u2_Display/lt94_c3 ;
  wire \u2_Display/lt94_c31 ;
  wire \u2_Display/lt94_c5 ;
  wire \u2_Display/lt94_c7 ;
  wire \u2_Display/lt94_c9 ;
  wire \u2_Display/lt95_c1 ;
  wire \u2_Display/lt95_c11 ;
  wire \u2_Display/lt95_c13 ;
  wire \u2_Display/lt95_c15 ;
  wire \u2_Display/lt95_c17 ;
  wire \u2_Display/lt95_c19 ;
  wire \u2_Display/lt95_c21 ;
  wire \u2_Display/lt95_c23 ;
  wire \u2_Display/lt95_c25 ;
  wire \u2_Display/lt95_c27 ;
  wire \u2_Display/lt95_c29 ;
  wire \u2_Display/lt95_c3 ;
  wire \u2_Display/lt95_c31 ;
  wire \u2_Display/lt95_c5 ;
  wire \u2_Display/lt95_c7 ;
  wire \u2_Display/lt95_c9 ;
  wire \u2_Display/lt96_c1 ;
  wire \u2_Display/lt96_c11 ;
  wire \u2_Display/lt96_c13 ;
  wire \u2_Display/lt96_c15 ;
  wire \u2_Display/lt96_c17 ;
  wire \u2_Display/lt96_c19 ;
  wire \u2_Display/lt96_c21 ;
  wire \u2_Display/lt96_c23 ;
  wire \u2_Display/lt96_c25 ;
  wire \u2_Display/lt96_c27 ;
  wire \u2_Display/lt96_c29 ;
  wire \u2_Display/lt96_c3 ;
  wire \u2_Display/lt96_c31 ;
  wire \u2_Display/lt96_c5 ;
  wire \u2_Display/lt96_c7 ;
  wire \u2_Display/lt96_c9 ;
  wire \u2_Display/lt97_c1 ;
  wire \u2_Display/lt97_c11 ;
  wire \u2_Display/lt97_c13 ;
  wire \u2_Display/lt97_c15 ;
  wire \u2_Display/lt97_c17 ;
  wire \u2_Display/lt97_c19 ;
  wire \u2_Display/lt97_c21 ;
  wire \u2_Display/lt97_c23 ;
  wire \u2_Display/lt97_c25 ;
  wire \u2_Display/lt97_c27 ;
  wire \u2_Display/lt97_c29 ;
  wire \u2_Display/lt97_c3 ;
  wire \u2_Display/lt97_c31 ;
  wire \u2_Display/lt97_c5 ;
  wire \u2_Display/lt97_c7 ;
  wire \u2_Display/lt97_c9 ;
  wire \u2_Display/lt98_c1 ;
  wire \u2_Display/lt98_c11 ;
  wire \u2_Display/lt98_c13 ;
  wire \u2_Display/lt98_c15 ;
  wire \u2_Display/lt98_c17 ;
  wire \u2_Display/lt98_c19 ;
  wire \u2_Display/lt98_c21 ;
  wire \u2_Display/lt98_c23 ;
  wire \u2_Display/lt98_c25 ;
  wire \u2_Display/lt98_c27 ;
  wire \u2_Display/lt98_c29 ;
  wire \u2_Display/lt98_c3 ;
  wire \u2_Display/lt98_c31 ;
  wire \u2_Display/lt98_c5 ;
  wire \u2_Display/lt98_c7 ;
  wire \u2_Display/lt98_c9 ;
  wire \u2_Display/lt99_c1 ;
  wire \u2_Display/lt99_c11 ;
  wire \u2_Display/lt99_c13 ;
  wire \u2_Display/lt99_c15 ;
  wire \u2_Display/lt99_c17 ;
  wire \u2_Display/lt99_c19 ;
  wire \u2_Display/lt99_c21 ;
  wire \u2_Display/lt99_c23 ;
  wire \u2_Display/lt99_c25 ;
  wire \u2_Display/lt99_c27 ;
  wire \u2_Display/lt99_c29 ;
  wire \u2_Display/lt99_c3 ;
  wire \u2_Display/lt99_c31 ;
  wire \u2_Display/lt99_c5 ;
  wire \u2_Display/lt99_c7 ;
  wire \u2_Display/lt99_c9 ;
  wire \u2_Display/lt9_2_c1 ;
  wire \u2_Display/lt9_2_c11 ;
  wire \u2_Display/lt9_2_c13 ;
  wire \u2_Display/lt9_2_c3 ;
  wire \u2_Display/lt9_2_c5 ;
  wire \u2_Display/lt9_2_c7 ;
  wire \u2_Display/lt9_2_c9 ;
  wire \u2_Display/mux11_b0_sel_is_0_o ;
  wire \u2_Display/mux19_b0_sel_is_0_o ;
  wire \u2_Display/mux21_b0_sel_is_0_o ;
  wire \u2_Display/mux5_b0_sel_is_0_o ;
  wire \u2_Display/n100 ;
  wire \u2_Display/n1000 ;
  wire \u2_Display/n1001 ;
  wire \u2_Display/n1002 ;
  wire \u2_Display/n1003 ;
  wire \u2_Display/n1004 ;
  wire \u2_Display/n1005 ;
  wire \u2_Display/n1006 ;
  wire \u2_Display/n1007 ;
  wire \u2_Display/n1008 ;
  wire \u2_Display/n1009 ;
  wire \u2_Display/n1010 ;
  wire \u2_Display/n1011 ;
  wire \u2_Display/n1012 ;
  wire \u2_Display/n1015 ;
  wire \u2_Display/n1016 ;
  wire \u2_Display/n1017 ;
  wire \u2_Display/n1018 ;
  wire \u2_Display/n1019 ;
  wire \u2_Display/n1020 ;
  wire \u2_Display/n1021 ;
  wire \u2_Display/n1022 ;
  wire \u2_Display/n1023 ;
  wire \u2_Display/n1024 ;
  wire \u2_Display/n1025 ;
  wire \u2_Display/n1026 ;
  wire \u2_Display/n1027 ;
  wire \u2_Display/n1028 ;
  wire \u2_Display/n1029 ;
  wire \u2_Display/n103 ;
  wire \u2_Display/n1030 ;
  wire \u2_Display/n1031 ;
  wire \u2_Display/n1032 ;
  wire \u2_Display/n1033 ;
  wire \u2_Display/n1034 ;
  wire \u2_Display/n1035 ;
  wire \u2_Display/n1036 ;
  wire \u2_Display/n1037 ;
  wire \u2_Display/n1038 ;
  wire \u2_Display/n1039 ;
  wire \u2_Display/n104 ;
  wire \u2_Display/n1040 ;
  wire \u2_Display/n1041 ;
  wire \u2_Display/n1042 ;
  wire \u2_Display/n1043 ;
  wire \u2_Display/n1044 ;
  wire \u2_Display/n1045 ;
  wire \u2_Display/n1046 ;
  wire \u2_Display/n1047 ;
  wire \u2_Display/n1050 ;
  wire \u2_Display/n1051 ;
  wire \u2_Display/n1052 ;
  wire \u2_Display/n1053 ;
  wire \u2_Display/n1054 ;
  wire \u2_Display/n1055 ;
  wire \u2_Display/n1056 ;
  wire \u2_Display/n1057 ;
  wire \u2_Display/n1058 ;
  wire \u2_Display/n1059 ;
  wire \u2_Display/n1060 ;
  wire \u2_Display/n1061 ;
  wire \u2_Display/n1062 ;
  wire \u2_Display/n1063 ;
  wire \u2_Display/n1064 ;
  wire \u2_Display/n1065 ;
  wire \u2_Display/n1066 ;
  wire \u2_Display/n1067 ;
  wire \u2_Display/n1068 ;
  wire \u2_Display/n1069 ;
  wire \u2_Display/n1070 ;
  wire \u2_Display/n1071 ;
  wire \u2_Display/n1072 ;
  wire \u2_Display/n1073 ;
  wire \u2_Display/n1074 ;
  wire \u2_Display/n1075 ;
  wire \u2_Display/n1076 ;
  wire \u2_Display/n1077 ;
  wire \u2_Display/n1078 ;
  wire \u2_Display/n1079 ;
  wire \u2_Display/n1080 ;
  wire \u2_Display/n1081 ;
  wire \u2_Display/n1082 ;
  wire \u2_Display/n1085 ;
  wire \u2_Display/n1086 ;
  wire \u2_Display/n1087 ;
  wire \u2_Display/n1088 ;
  wire \u2_Display/n1089 ;
  wire \u2_Display/n1090 ;
  wire \u2_Display/n1091 ;
  wire \u2_Display/n1092 ;
  wire \u2_Display/n1093 ;
  wire \u2_Display/n1094 ;
  wire \u2_Display/n1095 ;
  wire \u2_Display/n1096 ;
  wire \u2_Display/n1097 ;
  wire \u2_Display/n1098 ;
  wire \u2_Display/n1099 ;
  wire \u2_Display/n1100 ;
  wire \u2_Display/n1101 ;
  wire \u2_Display/n1102 ;
  wire \u2_Display/n1103 ;
  wire \u2_Display/n1104 ;
  wire \u2_Display/n1105 ;
  wire \u2_Display/n1106 ;
  wire \u2_Display/n1107 ;
  wire \u2_Display/n1108 ;
  wire \u2_Display/n1109 ;
  wire \u2_Display/n1110 ;
  wire \u2_Display/n1111 ;
  wire \u2_Display/n1112 ;
  wire \u2_Display/n1113 ;
  wire \u2_Display/n1114 ;
  wire \u2_Display/n1115 ;
  wire \u2_Display/n1116 ;
  wire \u2_Display/n1117 ;
  wire \u2_Display/n1120 ;
  wire \u2_Display/n1121 ;
  wire \u2_Display/n1122 ;
  wire \u2_Display/n1123 ;
  wire \u2_Display/n1124 ;
  wire \u2_Display/n1125 ;
  wire \u2_Display/n1126 ;
  wire \u2_Display/n1127 ;
  wire \u2_Display/n1128 ;
  wire \u2_Display/n1129 ;
  wire \u2_Display/n1130 ;
  wire \u2_Display/n1131 ;
  wire \u2_Display/n1132 ;
  wire \u2_Display/n1133 ;
  wire \u2_Display/n1134 ;
  wire \u2_Display/n1135 ;
  wire \u2_Display/n1136 ;
  wire \u2_Display/n1137 ;
  wire \u2_Display/n1138 ;
  wire \u2_Display/n1139 ;
  wire \u2_Display/n1140 ;
  wire \u2_Display/n1141 ;
  wire \u2_Display/n1142 ;
  wire \u2_Display/n1143 ;
  wire \u2_Display/n1144 ;
  wire \u2_Display/n1145 ;
  wire \u2_Display/n1146 ;
  wire \u2_Display/n1147 ;
  wire \u2_Display/n1148 ;
  wire \u2_Display/n1149 ;
  wire \u2_Display/n1150 ;
  wire \u2_Display/n1151 ;
  wire \u2_Display/n1152 ;
  wire \u2_Display/n1155 ;
  wire \u2_Display/n1156 ;
  wire \u2_Display/n1157 ;
  wire \u2_Display/n1158 ;
  wire \u2_Display/n1159 ;
  wire \u2_Display/n1160 ;
  wire \u2_Display/n1161 ;
  wire \u2_Display/n1162 ;
  wire \u2_Display/n1163 ;
  wire \u2_Display/n1164 ;
  wire \u2_Display/n1165 ;
  wire \u2_Display/n1166 ;
  wire \u2_Display/n1167 ;
  wire \u2_Display/n1168 ;
  wire \u2_Display/n1169 ;
  wire \u2_Display/n1170 ;
  wire \u2_Display/n1171 ;
  wire \u2_Display/n1172 ;
  wire \u2_Display/n1173 ;
  wire \u2_Display/n1174 ;
  wire \u2_Display/n1175 ;
  wire \u2_Display/n1176 ;
  wire \u2_Display/n1177 ;
  wire \u2_Display/n1178 ;
  wire \u2_Display/n1179 ;
  wire \u2_Display/n1180 ;
  wire \u2_Display/n1181 ;
  wire \u2_Display/n1182 ;
  wire \u2_Display/n1183 ;
  wire \u2_Display/n1184 ;
  wire \u2_Display/n1185 ;
  wire \u2_Display/n1186 ;
  wire \u2_Display/n1187 ;
  wire \u2_Display/n136 ;
  wire \u2_Display/n138 ;
  wire \u2_Display/n141 ;
  wire \u2_Display/n144 ;
  wire \u2_Display/n145 ;
  wire \u2_Display/n1540 ;
  wire \u2_Display/n1543 ;
  wire \u2_Display/n1544 ;
  wire \u2_Display/n1545 ;
  wire \u2_Display/n1546 ;
  wire \u2_Display/n1547 ;
  wire \u2_Display/n1548 ;
  wire \u2_Display/n1549 ;
  wire \u2_Display/n1550 ;
  wire \u2_Display/n1551 ;
  wire \u2_Display/n1552 ;
  wire \u2_Display/n1553 ;
  wire \u2_Display/n1554 ;
  wire \u2_Display/n1555 ;
  wire \u2_Display/n1556 ;
  wire \u2_Display/n1557 ;
  wire \u2_Display/n1558 ;
  wire \u2_Display/n1559 ;
  wire \u2_Display/n1560 ;
  wire \u2_Display/n1561 ;
  wire \u2_Display/n1562 ;
  wire \u2_Display/n1563 ;
  wire \u2_Display/n1564 ;
  wire \u2_Display/n1565 ;
  wire \u2_Display/n1566 ;
  wire \u2_Display/n1567 ;
  wire \u2_Display/n1568 ;
  wire \u2_Display/n1569 ;
  wire \u2_Display/n1570 ;
  wire \u2_Display/n1571 ;
  wire \u2_Display/n1572 ;
  wire \u2_Display/n1573 ;
  wire \u2_Display/n1574 ;
  wire \u2_Display/n1575 ;
  wire \u2_Display/n1578 ;
  wire \u2_Display/n1579 ;
  wire \u2_Display/n1580 ;
  wire \u2_Display/n1581 ;
  wire \u2_Display/n1582 ;
  wire \u2_Display/n1583 ;
  wire \u2_Display/n1584 ;
  wire \u2_Display/n1585 ;
  wire \u2_Display/n1586 ;
  wire \u2_Display/n1587 ;
  wire \u2_Display/n1588 ;
  wire \u2_Display/n1589 ;
  wire \u2_Display/n1590 ;
  wire \u2_Display/n1591 ;
  wire \u2_Display/n1592 ;
  wire \u2_Display/n1593 ;
  wire \u2_Display/n1594 ;
  wire \u2_Display/n1595 ;
  wire \u2_Display/n1596 ;
  wire \u2_Display/n1597 ;
  wire \u2_Display/n1598 ;
  wire \u2_Display/n1599 ;
  wire \u2_Display/n1600 ;
  wire \u2_Display/n1601 ;
  wire \u2_Display/n1602 ;
  wire \u2_Display/n1603 ;
  wire \u2_Display/n1604 ;
  wire \u2_Display/n1605 ;
  wire \u2_Display/n1606 ;
  wire \u2_Display/n1607 ;
  wire \u2_Display/n1608 ;
  wire \u2_Display/n1609 ;
  wire \u2_Display/n1610 ;
  wire \u2_Display/n1613 ;
  wire \u2_Display/n1614 ;
  wire \u2_Display/n1615 ;
  wire \u2_Display/n1616 ;
  wire \u2_Display/n1617 ;
  wire \u2_Display/n1618 ;
  wire \u2_Display/n1619 ;
  wire \u2_Display/n1620 ;
  wire \u2_Display/n1621 ;
  wire \u2_Display/n1622 ;
  wire \u2_Display/n1623 ;
  wire \u2_Display/n1624 ;
  wire \u2_Display/n1625 ;
  wire \u2_Display/n1626 ;
  wire \u2_Display/n1627 ;
  wire \u2_Display/n1628 ;
  wire \u2_Display/n1629 ;
  wire \u2_Display/n1630 ;
  wire \u2_Display/n1631 ;
  wire \u2_Display/n1632 ;
  wire \u2_Display/n1633 ;
  wire \u2_Display/n1634 ;
  wire \u2_Display/n1635 ;
  wire \u2_Display/n1636 ;
  wire \u2_Display/n1637 ;
  wire \u2_Display/n1638 ;
  wire \u2_Display/n1639 ;
  wire \u2_Display/n1640 ;
  wire \u2_Display/n1641 ;
  wire \u2_Display/n1642 ;
  wire \u2_Display/n1643 ;
  wire \u2_Display/n1644 ;
  wire \u2_Display/n1645 ;
  wire \u2_Display/n1648 ;
  wire \u2_Display/n1649 ;
  wire \u2_Display/n1650 ;
  wire \u2_Display/n1651 ;
  wire \u2_Display/n1652 ;
  wire \u2_Display/n1653 ;
  wire \u2_Display/n1654 ;
  wire \u2_Display/n1655 ;
  wire \u2_Display/n1656 ;
  wire \u2_Display/n1657 ;
  wire \u2_Display/n1658 ;
  wire \u2_Display/n1659 ;
  wire \u2_Display/n1660 ;
  wire \u2_Display/n1661 ;
  wire \u2_Display/n1662 ;
  wire \u2_Display/n1663 ;
  wire \u2_Display/n1664 ;
  wire \u2_Display/n1665 ;
  wire \u2_Display/n1666 ;
  wire \u2_Display/n1667 ;
  wire \u2_Display/n1668 ;
  wire \u2_Display/n1669 ;
  wire \u2_Display/n1670 ;
  wire \u2_Display/n1671 ;
  wire \u2_Display/n1672 ;
  wire \u2_Display/n1673 ;
  wire \u2_Display/n1674 ;
  wire \u2_Display/n1675 ;
  wire \u2_Display/n1676 ;
  wire \u2_Display/n1677 ;
  wire \u2_Display/n1678 ;
  wire \u2_Display/n1679 ;
  wire \u2_Display/n1680 ;
  wire \u2_Display/n1683 ;
  wire \u2_Display/n1684 ;
  wire \u2_Display/n1685 ;
  wire \u2_Display/n1686 ;
  wire \u2_Display/n1687 ;
  wire \u2_Display/n1688 ;
  wire \u2_Display/n1689 ;
  wire \u2_Display/n1690 ;
  wire \u2_Display/n1691 ;
  wire \u2_Display/n1692 ;
  wire \u2_Display/n1693 ;
  wire \u2_Display/n1694 ;
  wire \u2_Display/n1695 ;
  wire \u2_Display/n1696 ;
  wire \u2_Display/n1697 ;
  wire \u2_Display/n1698 ;
  wire \u2_Display/n1699 ;
  wire \u2_Display/n1700 ;
  wire \u2_Display/n1701 ;
  wire \u2_Display/n1702 ;
  wire \u2_Display/n1703 ;
  wire \u2_Display/n1704 ;
  wire \u2_Display/n1705 ;
  wire \u2_Display/n1706 ;
  wire \u2_Display/n1707 ;
  wire \u2_Display/n1708 ;
  wire \u2_Display/n1709 ;
  wire \u2_Display/n1710 ;
  wire \u2_Display/n1711 ;
  wire \u2_Display/n1712 ;
  wire \u2_Display/n1713 ;
  wire \u2_Display/n1714 ;
  wire \u2_Display/n1715 ;
  wire \u2_Display/n1718 ;
  wire \u2_Display/n1719 ;
  wire \u2_Display/n1720 ;
  wire \u2_Display/n1721 ;
  wire \u2_Display/n1722 ;
  wire \u2_Display/n1723 ;
  wire \u2_Display/n1724 ;
  wire \u2_Display/n1725 ;
  wire \u2_Display/n1726 ;
  wire \u2_Display/n1727 ;
  wire \u2_Display/n1728 ;
  wire \u2_Display/n1729 ;
  wire \u2_Display/n1730 ;
  wire \u2_Display/n1731 ;
  wire \u2_Display/n1732 ;
  wire \u2_Display/n1733 ;
  wire \u2_Display/n1734 ;
  wire \u2_Display/n1735 ;
  wire \u2_Display/n1736 ;
  wire \u2_Display/n1737 ;
  wire \u2_Display/n1738 ;
  wire \u2_Display/n1739 ;
  wire \u2_Display/n1740 ;
  wire \u2_Display/n1741 ;
  wire \u2_Display/n1742 ;
  wire \u2_Display/n1743 ;
  wire \u2_Display/n1744 ;
  wire \u2_Display/n1745 ;
  wire \u2_Display/n1746 ;
  wire \u2_Display/n1747 ;
  wire \u2_Display/n1748 ;
  wire \u2_Display/n1749 ;
  wire \u2_Display/n1750 ;
  wire \u2_Display/n1753 ;
  wire \u2_Display/n1754 ;
  wire \u2_Display/n1755 ;
  wire \u2_Display/n1756 ;
  wire \u2_Display/n1757 ;
  wire \u2_Display/n1758 ;
  wire \u2_Display/n1759 ;
  wire \u2_Display/n1760 ;
  wire \u2_Display/n1761 ;
  wire \u2_Display/n1762 ;
  wire \u2_Display/n1763 ;
  wire \u2_Display/n1764 ;
  wire \u2_Display/n1765 ;
  wire \u2_Display/n1766 ;
  wire \u2_Display/n1767 ;
  wire \u2_Display/n1768 ;
  wire \u2_Display/n1769 ;
  wire \u2_Display/n1770 ;
  wire \u2_Display/n1771 ;
  wire \u2_Display/n1772 ;
  wire \u2_Display/n1773 ;
  wire \u2_Display/n1774 ;
  wire \u2_Display/n1775 ;
  wire \u2_Display/n1776 ;
  wire \u2_Display/n1777 ;
  wire \u2_Display/n1778 ;
  wire \u2_Display/n1779 ;
  wire \u2_Display/n1780 ;
  wire \u2_Display/n1781 ;
  wire \u2_Display/n1782 ;
  wire \u2_Display/n1783 ;
  wire \u2_Display/n1784 ;
  wire \u2_Display/n1785 ;
  wire \u2_Display/n1788 ;
  wire \u2_Display/n1789 ;
  wire \u2_Display/n1790 ;
  wire \u2_Display/n1791 ;
  wire \u2_Display/n1792 ;
  wire \u2_Display/n1793 ;
  wire \u2_Display/n1794 ;
  wire \u2_Display/n1795 ;
  wire \u2_Display/n1796 ;
  wire \u2_Display/n1797 ;
  wire \u2_Display/n1798 ;
  wire \u2_Display/n1799 ;
  wire \u2_Display/n1800 ;
  wire \u2_Display/n1801 ;
  wire \u2_Display/n1802 ;
  wire \u2_Display/n1803 ;
  wire \u2_Display/n1804 ;
  wire \u2_Display/n1805 ;
  wire \u2_Display/n1806 ;
  wire \u2_Display/n1807 ;
  wire \u2_Display/n1808 ;
  wire \u2_Display/n1809 ;
  wire \u2_Display/n1810 ;
  wire \u2_Display/n1811 ;
  wire \u2_Display/n1812 ;
  wire \u2_Display/n1813 ;
  wire \u2_Display/n1814 ;
  wire \u2_Display/n1815 ;
  wire \u2_Display/n1816 ;
  wire \u2_Display/n1817 ;
  wire \u2_Display/n1818 ;
  wire \u2_Display/n1819 ;
  wire \u2_Display/n1820 ;
  wire \u2_Display/n1823 ;
  wire \u2_Display/n1824 ;
  wire \u2_Display/n1825 ;
  wire \u2_Display/n1826 ;
  wire \u2_Display/n1827 ;
  wire \u2_Display/n1828 ;
  wire \u2_Display/n1829 ;
  wire \u2_Display/n1830 ;
  wire \u2_Display/n1831 ;
  wire \u2_Display/n1832 ;
  wire \u2_Display/n1833 ;
  wire \u2_Display/n1834 ;
  wire \u2_Display/n1835 ;
  wire \u2_Display/n1836 ;
  wire \u2_Display/n1837 ;
  wire \u2_Display/n1838 ;
  wire \u2_Display/n1839 ;
  wire \u2_Display/n1840 ;
  wire \u2_Display/n1841 ;
  wire \u2_Display/n1842 ;
  wire \u2_Display/n1843 ;
  wire \u2_Display/n1844 ;
  wire \u2_Display/n1845 ;
  wire \u2_Display/n1846 ;
  wire \u2_Display/n1847 ;
  wire \u2_Display/n1848 ;
  wire \u2_Display/n1849 ;
  wire \u2_Display/n1850 ;
  wire \u2_Display/n1851 ;
  wire \u2_Display/n1852 ;
  wire \u2_Display/n1853 ;
  wire \u2_Display/n1854 ;
  wire \u2_Display/n1855 ;
  wire \u2_Display/n1858 ;
  wire \u2_Display/n1859 ;
  wire \u2_Display/n1860 ;
  wire \u2_Display/n1861 ;
  wire \u2_Display/n1862 ;
  wire \u2_Display/n1863 ;
  wire \u2_Display/n1864 ;
  wire \u2_Display/n1865 ;
  wire \u2_Display/n1866 ;
  wire \u2_Display/n1867 ;
  wire \u2_Display/n1868 ;
  wire \u2_Display/n1869 ;
  wire \u2_Display/n1870 ;
  wire \u2_Display/n1871 ;
  wire \u2_Display/n1872 ;
  wire \u2_Display/n1873 ;
  wire \u2_Display/n1874 ;
  wire \u2_Display/n1875 ;
  wire \u2_Display/n1876 ;
  wire \u2_Display/n1877 ;
  wire \u2_Display/n1878 ;
  wire \u2_Display/n1879 ;
  wire \u2_Display/n1880 ;
  wire \u2_Display/n1881 ;
  wire \u2_Display/n1882 ;
  wire \u2_Display/n1883 ;
  wire \u2_Display/n1884 ;
  wire \u2_Display/n1885 ;
  wire \u2_Display/n1886 ;
  wire \u2_Display/n1887 ;
  wire \u2_Display/n1888 ;
  wire \u2_Display/n1889 ;
  wire \u2_Display/n1890 ;
  wire \u2_Display/n1893 ;
  wire \u2_Display/n1894 ;
  wire \u2_Display/n1895 ;
  wire \u2_Display/n1896 ;
  wire \u2_Display/n1897 ;
  wire \u2_Display/n1898 ;
  wire \u2_Display/n1899 ;
  wire \u2_Display/n1900 ;
  wire \u2_Display/n1901 ;
  wire \u2_Display/n1902 ;
  wire \u2_Display/n1903 ;
  wire \u2_Display/n1904 ;
  wire \u2_Display/n1905 ;
  wire \u2_Display/n1906 ;
  wire \u2_Display/n1907 ;
  wire \u2_Display/n1908 ;
  wire \u2_Display/n1909 ;
  wire \u2_Display/n1910 ;
  wire \u2_Display/n1911 ;
  wire \u2_Display/n1912 ;
  wire \u2_Display/n1913 ;
  wire \u2_Display/n1914 ;
  wire \u2_Display/n1915 ;
  wire \u2_Display/n1916 ;
  wire \u2_Display/n1917 ;
  wire \u2_Display/n1918 ;
  wire \u2_Display/n1919 ;
  wire \u2_Display/n1920 ;
  wire \u2_Display/n1921 ;
  wire \u2_Display/n1922 ;
  wire \u2_Display/n1923 ;
  wire \u2_Display/n1924 ;
  wire \u2_Display/n1925 ;
  wire \u2_Display/n1928 ;
  wire \u2_Display/n1929 ;
  wire \u2_Display/n1930 ;
  wire \u2_Display/n1931 ;
  wire \u2_Display/n1932 ;
  wire \u2_Display/n1933 ;
  wire \u2_Display/n1934 ;
  wire \u2_Display/n1935 ;
  wire \u2_Display/n1936 ;
  wire \u2_Display/n1937 ;
  wire \u2_Display/n1938 ;
  wire \u2_Display/n1939 ;
  wire \u2_Display/n1940 ;
  wire \u2_Display/n1941 ;
  wire \u2_Display/n1942 ;
  wire \u2_Display/n1943 ;
  wire \u2_Display/n1944 ;
  wire \u2_Display/n1945 ;
  wire \u2_Display/n1946 ;
  wire \u2_Display/n1947 ;
  wire \u2_Display/n1948 ;
  wire \u2_Display/n1949 ;
  wire \u2_Display/n1950 ;
  wire \u2_Display/n1951 ;
  wire \u2_Display/n1952 ;
  wire \u2_Display/n1953 ;
  wire \u2_Display/n1954 ;
  wire \u2_Display/n1955 ;
  wire \u2_Display/n1956 ;
  wire \u2_Display/n1957 ;
  wire \u2_Display/n1958 ;
  wire \u2_Display/n1959 ;
  wire \u2_Display/n1960 ;
  wire \u2_Display/n1963 ;
  wire \u2_Display/n1964 ;
  wire \u2_Display/n1965 ;
  wire \u2_Display/n1966 ;
  wire \u2_Display/n1967 ;
  wire \u2_Display/n1968 ;
  wire \u2_Display/n1969 ;
  wire \u2_Display/n1970 ;
  wire \u2_Display/n1971 ;
  wire \u2_Display/n1972 ;
  wire \u2_Display/n1973 ;
  wire \u2_Display/n1974 ;
  wire \u2_Display/n1975 ;
  wire \u2_Display/n1976 ;
  wire \u2_Display/n1977 ;
  wire \u2_Display/n1978 ;
  wire \u2_Display/n1979 ;
  wire \u2_Display/n1980 ;
  wire \u2_Display/n1981 ;
  wire \u2_Display/n1982 ;
  wire \u2_Display/n1983 ;
  wire \u2_Display/n1984 ;
  wire \u2_Display/n1985 ;
  wire \u2_Display/n1986 ;
  wire \u2_Display/n1987 ;
  wire \u2_Display/n1988 ;
  wire \u2_Display/n1989 ;
  wire \u2_Display/n1990 ;
  wire \u2_Display/n1991 ;
  wire \u2_Display/n1992 ;
  wire \u2_Display/n1993 ;
  wire \u2_Display/n1994 ;
  wire \u2_Display/n1995 ;
  wire \u2_Display/n1998 ;
  wire \u2_Display/n1999 ;
  wire \u2_Display/n2000 ;
  wire \u2_Display/n2001 ;
  wire \u2_Display/n2002 ;
  wire \u2_Display/n2003 ;
  wire \u2_Display/n2004 ;
  wire \u2_Display/n2005 ;
  wire \u2_Display/n2006 ;
  wire \u2_Display/n2007 ;
  wire \u2_Display/n2008 ;
  wire \u2_Display/n2009 ;
  wire \u2_Display/n2010 ;
  wire \u2_Display/n2011 ;
  wire \u2_Display/n2012 ;
  wire \u2_Display/n2013 ;
  wire \u2_Display/n2014 ;
  wire \u2_Display/n2015 ;
  wire \u2_Display/n2016 ;
  wire \u2_Display/n2017 ;
  wire \u2_Display/n2018 ;
  wire \u2_Display/n2019 ;
  wire \u2_Display/n2020 ;
  wire \u2_Display/n2021 ;
  wire \u2_Display/n2022 ;
  wire \u2_Display/n2023 ;
  wire \u2_Display/n2024 ;
  wire \u2_Display/n2025 ;
  wire \u2_Display/n2026 ;
  wire \u2_Display/n2027 ;
  wire \u2_Display/n2028 ;
  wire \u2_Display/n2029 ;
  wire \u2_Display/n2030 ;
  wire \u2_Display/n2033 ;
  wire \u2_Display/n2034 ;
  wire \u2_Display/n2035 ;
  wire \u2_Display/n2036 ;
  wire \u2_Display/n2037 ;
  wire \u2_Display/n2038 ;
  wire \u2_Display/n2039 ;
  wire \u2_Display/n2040 ;
  wire \u2_Display/n2041 ;
  wire \u2_Display/n2042 ;
  wire \u2_Display/n2043 ;
  wire \u2_Display/n2044 ;
  wire \u2_Display/n2045 ;
  wire \u2_Display/n2046 ;
  wire \u2_Display/n2047 ;
  wire \u2_Display/n2048 ;
  wire \u2_Display/n2049 ;
  wire \u2_Display/n2050 ;
  wire \u2_Display/n2051 ;
  wire \u2_Display/n2052 ;
  wire \u2_Display/n2053 ;
  wire \u2_Display/n2054 ;
  wire \u2_Display/n2055 ;
  wire \u2_Display/n2056 ;
  wire \u2_Display/n2057 ;
  wire \u2_Display/n2058 ;
  wire \u2_Display/n2059 ;
  wire \u2_Display/n2060 ;
  wire \u2_Display/n2061 ;
  wire \u2_Display/n2062 ;
  wire \u2_Display/n2063 ;
  wire \u2_Display/n2064 ;
  wire \u2_Display/n2065 ;
  wire \u2_Display/n2068 ;
  wire \u2_Display/n2069 ;
  wire \u2_Display/n2070 ;
  wire \u2_Display/n2071 ;
  wire \u2_Display/n2072 ;
  wire \u2_Display/n2073 ;
  wire \u2_Display/n2074 ;
  wire \u2_Display/n2075 ;
  wire \u2_Display/n2076 ;
  wire \u2_Display/n2077 ;
  wire \u2_Display/n2078 ;
  wire \u2_Display/n2079 ;
  wire \u2_Display/n2080 ;
  wire \u2_Display/n2081 ;
  wire \u2_Display/n2082 ;
  wire \u2_Display/n2083 ;
  wire \u2_Display/n2084 ;
  wire \u2_Display/n2085 ;
  wire \u2_Display/n2086 ;
  wire \u2_Display/n2087 ;
  wire \u2_Display/n2088 ;
  wire \u2_Display/n2089 ;
  wire \u2_Display/n2090 ;
  wire \u2_Display/n2091 ;
  wire \u2_Display/n2092 ;
  wire \u2_Display/n2093 ;
  wire \u2_Display/n2094 ;
  wire \u2_Display/n2095 ;
  wire \u2_Display/n2096 ;
  wire \u2_Display/n2097 ;
  wire \u2_Display/n2098 ;
  wire \u2_Display/n2099 ;
  wire \u2_Display/n2100 ;
  wire \u2_Display/n2103 ;
  wire \u2_Display/n2104 ;
  wire \u2_Display/n2105 ;
  wire \u2_Display/n2106 ;
  wire \u2_Display/n2107 ;
  wire \u2_Display/n2108 ;
  wire \u2_Display/n2109 ;
  wire \u2_Display/n2110 ;
  wire \u2_Display/n2111 ;
  wire \u2_Display/n2112 ;
  wire \u2_Display/n2113 ;
  wire \u2_Display/n2114 ;
  wire \u2_Display/n2115 ;
  wire \u2_Display/n2116 ;
  wire \u2_Display/n2117 ;
  wire \u2_Display/n2118 ;
  wire \u2_Display/n2119 ;
  wire \u2_Display/n2120 ;
  wire \u2_Display/n2121 ;
  wire \u2_Display/n2122 ;
  wire \u2_Display/n2123 ;
  wire \u2_Display/n2124 ;
  wire \u2_Display/n2125 ;
  wire \u2_Display/n2126 ;
  wire \u2_Display/n2127 ;
  wire \u2_Display/n2128 ;
  wire \u2_Display/n2129 ;
  wire \u2_Display/n2130 ;
  wire \u2_Display/n2131 ;
  wire \u2_Display/n2132 ;
  wire \u2_Display/n2133 ;
  wire \u2_Display/n2134 ;
  wire \u2_Display/n2135 ;
  wire \u2_Display/n2138 ;
  wire \u2_Display/n2139 ;
  wire \u2_Display/n2140 ;
  wire \u2_Display/n2141 ;
  wire \u2_Display/n2142 ;
  wire \u2_Display/n2143 ;
  wire \u2_Display/n2144 ;
  wire \u2_Display/n2145 ;
  wire \u2_Display/n2146 ;
  wire \u2_Display/n2147 ;
  wire \u2_Display/n2148 ;
  wire \u2_Display/n2149 ;
  wire \u2_Display/n2150 ;
  wire \u2_Display/n2151 ;
  wire \u2_Display/n2152 ;
  wire \u2_Display/n2153 ;
  wire \u2_Display/n2154 ;
  wire \u2_Display/n2155 ;
  wire \u2_Display/n2156 ;
  wire \u2_Display/n2157 ;
  wire \u2_Display/n2158 ;
  wire \u2_Display/n2159 ;
  wire \u2_Display/n2160 ;
  wire \u2_Display/n2161 ;
  wire \u2_Display/n2162 ;
  wire \u2_Display/n2163 ;
  wire \u2_Display/n2164 ;
  wire \u2_Display/n2165 ;
  wire \u2_Display/n2166 ;
  wire \u2_Display/n2167 ;
  wire \u2_Display/n2168 ;
  wire \u2_Display/n2169 ;
  wire \u2_Display/n2170 ;
  wire \u2_Display/n2173 ;
  wire \u2_Display/n2174 ;
  wire \u2_Display/n2175 ;
  wire \u2_Display/n2176 ;
  wire \u2_Display/n2177 ;
  wire \u2_Display/n2178 ;
  wire \u2_Display/n2179 ;
  wire \u2_Display/n2180 ;
  wire \u2_Display/n2181 ;
  wire \u2_Display/n2182 ;
  wire \u2_Display/n2183 ;
  wire \u2_Display/n2184 ;
  wire \u2_Display/n2185 ;
  wire \u2_Display/n2186 ;
  wire \u2_Display/n2187 ;
  wire \u2_Display/n2188 ;
  wire \u2_Display/n2189 ;
  wire \u2_Display/n2190 ;
  wire \u2_Display/n2191 ;
  wire \u2_Display/n2192 ;
  wire \u2_Display/n2193 ;
  wire \u2_Display/n2194 ;
  wire \u2_Display/n2195 ;
  wire \u2_Display/n2196 ;
  wire \u2_Display/n2197 ;
  wire \u2_Display/n2198 ;
  wire \u2_Display/n2199 ;
  wire \u2_Display/n2200 ;
  wire \u2_Display/n2201 ;
  wire \u2_Display/n2202 ;
  wire \u2_Display/n2203 ;
  wire \u2_Display/n2204 ;
  wire \u2_Display/n2205 ;
  wire \u2_Display/n2208 ;
  wire \u2_Display/n2209 ;
  wire \u2_Display/n2210 ;
  wire \u2_Display/n2211 ;
  wire \u2_Display/n2212 ;
  wire \u2_Display/n2213 ;
  wire \u2_Display/n2214 ;
  wire \u2_Display/n2215 ;
  wire \u2_Display/n2216 ;
  wire \u2_Display/n2217 ;
  wire \u2_Display/n2218 ;
  wire \u2_Display/n2219 ;
  wire \u2_Display/n2220 ;
  wire \u2_Display/n2221 ;
  wire \u2_Display/n2222 ;
  wire \u2_Display/n2223 ;
  wire \u2_Display/n2224 ;
  wire \u2_Display/n2225 ;
  wire \u2_Display/n2226 ;
  wire \u2_Display/n2227 ;
  wire \u2_Display/n2228 ;
  wire \u2_Display/n2229 ;
  wire \u2_Display/n2230 ;
  wire \u2_Display/n2231 ;
  wire \u2_Display/n2232 ;
  wire \u2_Display/n2233 ;
  wire \u2_Display/n2234 ;
  wire \u2_Display/n2235 ;
  wire \u2_Display/n2236 ;
  wire \u2_Display/n2237 ;
  wire \u2_Display/n2238 ;
  wire \u2_Display/n2239 ;
  wire \u2_Display/n2240 ;
  wire \u2_Display/n2243 ;
  wire \u2_Display/n2244 ;
  wire \u2_Display/n2245 ;
  wire \u2_Display/n2246 ;
  wire \u2_Display/n2247 ;
  wire \u2_Display/n2248 ;
  wire \u2_Display/n2249 ;
  wire \u2_Display/n2250 ;
  wire \u2_Display/n2251 ;
  wire \u2_Display/n2252 ;
  wire \u2_Display/n2253 ;
  wire \u2_Display/n2254 ;
  wire \u2_Display/n2255 ;
  wire \u2_Display/n2256 ;
  wire \u2_Display/n2257 ;
  wire \u2_Display/n2258 ;
  wire \u2_Display/n2259 ;
  wire \u2_Display/n2260 ;
  wire \u2_Display/n2261 ;
  wire \u2_Display/n2262 ;
  wire \u2_Display/n2263 ;
  wire \u2_Display/n2264 ;
  wire \u2_Display/n2265 ;
  wire \u2_Display/n2266 ;
  wire \u2_Display/n2267 ;
  wire \u2_Display/n2268 ;
  wire \u2_Display/n2269 ;
  wire \u2_Display/n2270 ;
  wire \u2_Display/n2271 ;
  wire \u2_Display/n2272 ;
  wire \u2_Display/n2273 ;
  wire \u2_Display/n2274 ;
  wire \u2_Display/n2275 ;
  wire \u2_Display/n2278 ;
  wire \u2_Display/n2279 ;
  wire \u2_Display/n2280 ;
  wire \u2_Display/n2281 ;
  wire \u2_Display/n2282 ;
  wire \u2_Display/n2283 ;
  wire \u2_Display/n2284 ;
  wire \u2_Display/n2285 ;
  wire \u2_Display/n2286 ;
  wire \u2_Display/n2287 ;
  wire \u2_Display/n2288 ;
  wire \u2_Display/n2289 ;
  wire \u2_Display/n2290 ;
  wire \u2_Display/n2291 ;
  wire \u2_Display/n2292 ;
  wire \u2_Display/n2293 ;
  wire \u2_Display/n2294 ;
  wire \u2_Display/n2295 ;
  wire \u2_Display/n2296 ;
  wire \u2_Display/n2297 ;
  wire \u2_Display/n2298 ;
  wire \u2_Display/n2299 ;
  wire \u2_Display/n2300 ;
  wire \u2_Display/n2301 ;
  wire \u2_Display/n2302 ;
  wire \u2_Display/n2303 ;
  wire \u2_Display/n2304 ;
  wire \u2_Display/n2305 ;
  wire \u2_Display/n2306 ;
  wire \u2_Display/n2307 ;
  wire \u2_Display/n2308 ;
  wire \u2_Display/n2309 ;
  wire \u2_Display/n2310 ;
  wire \u2_Display/n2663 ;
  wire \u2_Display/n2666 ;
  wire \u2_Display/n2667 ;
  wire \u2_Display/n2668 ;
  wire \u2_Display/n2669 ;
  wire \u2_Display/n2670 ;
  wire \u2_Display/n2671 ;
  wire \u2_Display/n2672 ;
  wire \u2_Display/n2673 ;
  wire \u2_Display/n2674 ;
  wire \u2_Display/n2675 ;
  wire \u2_Display/n2676 ;
  wire \u2_Display/n2677 ;
  wire \u2_Display/n2678 ;
  wire \u2_Display/n2679 ;
  wire \u2_Display/n2680 ;
  wire \u2_Display/n2681 ;
  wire \u2_Display/n2682 ;
  wire \u2_Display/n2683 ;
  wire \u2_Display/n2684 ;
  wire \u2_Display/n2685 ;
  wire \u2_Display/n2686 ;
  wire \u2_Display/n2687 ;
  wire \u2_Display/n2688 ;
  wire \u2_Display/n2689 ;
  wire \u2_Display/n2690 ;
  wire \u2_Display/n2691 ;
  wire \u2_Display/n2692 ;
  wire \u2_Display/n2693 ;
  wire \u2_Display/n2694 ;
  wire \u2_Display/n2695 ;
  wire \u2_Display/n2696 ;
  wire \u2_Display/n2697 ;
  wire \u2_Display/n2698 ;
  wire \u2_Display/n2701 ;
  wire \u2_Display/n2702 ;
  wire \u2_Display/n2703 ;
  wire \u2_Display/n2704 ;
  wire \u2_Display/n2705 ;
  wire \u2_Display/n2706 ;
  wire \u2_Display/n2707 ;
  wire \u2_Display/n2708 ;
  wire \u2_Display/n2709 ;
  wire \u2_Display/n2710 ;
  wire \u2_Display/n2711 ;
  wire \u2_Display/n2712 ;
  wire \u2_Display/n2713 ;
  wire \u2_Display/n2714 ;
  wire \u2_Display/n2715 ;
  wire \u2_Display/n2716 ;
  wire \u2_Display/n2717 ;
  wire \u2_Display/n2718 ;
  wire \u2_Display/n2719 ;
  wire \u2_Display/n2720 ;
  wire \u2_Display/n2721 ;
  wire \u2_Display/n2722 ;
  wire \u2_Display/n2723 ;
  wire \u2_Display/n2724 ;
  wire \u2_Display/n2725 ;
  wire \u2_Display/n2726 ;
  wire \u2_Display/n2727 ;
  wire \u2_Display/n2728 ;
  wire \u2_Display/n2729 ;
  wire \u2_Display/n2730 ;
  wire \u2_Display/n2731 ;
  wire \u2_Display/n2732 ;
  wire \u2_Display/n2733 ;
  wire \u2_Display/n2736 ;
  wire \u2_Display/n2737 ;
  wire \u2_Display/n2738 ;
  wire \u2_Display/n2739 ;
  wire \u2_Display/n2740 ;
  wire \u2_Display/n2741 ;
  wire \u2_Display/n2742 ;
  wire \u2_Display/n2743 ;
  wire \u2_Display/n2744 ;
  wire \u2_Display/n2745 ;
  wire \u2_Display/n2746 ;
  wire \u2_Display/n2747 ;
  wire \u2_Display/n2748 ;
  wire \u2_Display/n2749 ;
  wire \u2_Display/n2750 ;
  wire \u2_Display/n2751 ;
  wire \u2_Display/n2752 ;
  wire \u2_Display/n2753 ;
  wire \u2_Display/n2754 ;
  wire \u2_Display/n2755 ;
  wire \u2_Display/n2756 ;
  wire \u2_Display/n2757 ;
  wire \u2_Display/n2758 ;
  wire \u2_Display/n2759 ;
  wire \u2_Display/n2760 ;
  wire \u2_Display/n2761 ;
  wire \u2_Display/n2762 ;
  wire \u2_Display/n2763 ;
  wire \u2_Display/n2764 ;
  wire \u2_Display/n2765 ;
  wire \u2_Display/n2766 ;
  wire \u2_Display/n2767 ;
  wire \u2_Display/n2768 ;
  wire \u2_Display/n2771 ;
  wire \u2_Display/n2772 ;
  wire \u2_Display/n2773 ;
  wire \u2_Display/n2774 ;
  wire \u2_Display/n2775 ;
  wire \u2_Display/n2776 ;
  wire \u2_Display/n2777 ;
  wire \u2_Display/n2778 ;
  wire \u2_Display/n2779 ;
  wire \u2_Display/n2780 ;
  wire \u2_Display/n2781 ;
  wire \u2_Display/n2782 ;
  wire \u2_Display/n2783 ;
  wire \u2_Display/n2784 ;
  wire \u2_Display/n2785 ;
  wire \u2_Display/n2786 ;
  wire \u2_Display/n2787 ;
  wire \u2_Display/n2788 ;
  wire \u2_Display/n2789 ;
  wire \u2_Display/n2790 ;
  wire \u2_Display/n2791 ;
  wire \u2_Display/n2792 ;
  wire \u2_Display/n2793 ;
  wire \u2_Display/n2794 ;
  wire \u2_Display/n2795 ;
  wire \u2_Display/n2796 ;
  wire \u2_Display/n2797 ;
  wire \u2_Display/n2798 ;
  wire \u2_Display/n2799 ;
  wire \u2_Display/n2800 ;
  wire \u2_Display/n2801 ;
  wire \u2_Display/n2802 ;
  wire \u2_Display/n2803 ;
  wire \u2_Display/n2806 ;
  wire \u2_Display/n2807 ;
  wire \u2_Display/n2808 ;
  wire \u2_Display/n2809 ;
  wire \u2_Display/n2810 ;
  wire \u2_Display/n2811 ;
  wire \u2_Display/n2812 ;
  wire \u2_Display/n2813 ;
  wire \u2_Display/n2814 ;
  wire \u2_Display/n2815 ;
  wire \u2_Display/n2816 ;
  wire \u2_Display/n2817 ;
  wire \u2_Display/n2818 ;
  wire \u2_Display/n2819 ;
  wire \u2_Display/n2820 ;
  wire \u2_Display/n2821 ;
  wire \u2_Display/n2822 ;
  wire \u2_Display/n2823 ;
  wire \u2_Display/n2824 ;
  wire \u2_Display/n2825 ;
  wire \u2_Display/n2826 ;
  wire \u2_Display/n2827 ;
  wire \u2_Display/n2828 ;
  wire \u2_Display/n2829 ;
  wire \u2_Display/n2830 ;
  wire \u2_Display/n2831 ;
  wire \u2_Display/n2832 ;
  wire \u2_Display/n2833 ;
  wire \u2_Display/n2834 ;
  wire \u2_Display/n2835 ;
  wire \u2_Display/n2836 ;
  wire \u2_Display/n2837 ;
  wire \u2_Display/n2838 ;
  wire \u2_Display/n2841 ;
  wire \u2_Display/n2842 ;
  wire \u2_Display/n2843 ;
  wire \u2_Display/n2844 ;
  wire \u2_Display/n2845 ;
  wire \u2_Display/n2846 ;
  wire \u2_Display/n2847 ;
  wire \u2_Display/n2848 ;
  wire \u2_Display/n2849 ;
  wire \u2_Display/n2850 ;
  wire \u2_Display/n2851 ;
  wire \u2_Display/n2852 ;
  wire \u2_Display/n2853 ;
  wire \u2_Display/n2854 ;
  wire \u2_Display/n2855 ;
  wire \u2_Display/n2856 ;
  wire \u2_Display/n2857 ;
  wire \u2_Display/n2858 ;
  wire \u2_Display/n2859 ;
  wire \u2_Display/n2860 ;
  wire \u2_Display/n2861 ;
  wire \u2_Display/n2862 ;
  wire \u2_Display/n2863 ;
  wire \u2_Display/n2864 ;
  wire \u2_Display/n2865 ;
  wire \u2_Display/n2866 ;
  wire \u2_Display/n2867 ;
  wire \u2_Display/n2868 ;
  wire \u2_Display/n2869 ;
  wire \u2_Display/n2870 ;
  wire \u2_Display/n2871 ;
  wire \u2_Display/n2872 ;
  wire \u2_Display/n2873 ;
  wire \u2_Display/n2876 ;
  wire \u2_Display/n2877 ;
  wire \u2_Display/n2878 ;
  wire \u2_Display/n2879 ;
  wire \u2_Display/n2880 ;
  wire \u2_Display/n2881 ;
  wire \u2_Display/n2882 ;
  wire \u2_Display/n2883 ;
  wire \u2_Display/n2884 ;
  wire \u2_Display/n2885 ;
  wire \u2_Display/n2886 ;
  wire \u2_Display/n2887 ;
  wire \u2_Display/n2888 ;
  wire \u2_Display/n2889 ;
  wire \u2_Display/n2890 ;
  wire \u2_Display/n2891 ;
  wire \u2_Display/n2892 ;
  wire \u2_Display/n2893 ;
  wire \u2_Display/n2894 ;
  wire \u2_Display/n2895 ;
  wire \u2_Display/n2896 ;
  wire \u2_Display/n2897 ;
  wire \u2_Display/n2898 ;
  wire \u2_Display/n2899 ;
  wire \u2_Display/n2900 ;
  wire \u2_Display/n2901 ;
  wire \u2_Display/n2902 ;
  wire \u2_Display/n2903 ;
  wire \u2_Display/n2904 ;
  wire \u2_Display/n2905 ;
  wire \u2_Display/n2906 ;
  wire \u2_Display/n2907 ;
  wire \u2_Display/n2908 ;
  wire \u2_Display/n2911 ;
  wire \u2_Display/n2912 ;
  wire \u2_Display/n2913 ;
  wire \u2_Display/n2914 ;
  wire \u2_Display/n2915 ;
  wire \u2_Display/n2916 ;
  wire \u2_Display/n2917 ;
  wire \u2_Display/n2918 ;
  wire \u2_Display/n2919 ;
  wire \u2_Display/n2920 ;
  wire \u2_Display/n2921 ;
  wire \u2_Display/n2922 ;
  wire \u2_Display/n2923 ;
  wire \u2_Display/n2924 ;
  wire \u2_Display/n2925 ;
  wire \u2_Display/n2926 ;
  wire \u2_Display/n2927 ;
  wire \u2_Display/n2928 ;
  wire \u2_Display/n2929 ;
  wire \u2_Display/n2930 ;
  wire \u2_Display/n2931 ;
  wire \u2_Display/n2932 ;
  wire \u2_Display/n2933 ;
  wire \u2_Display/n2934 ;
  wire \u2_Display/n2935 ;
  wire \u2_Display/n2936 ;
  wire \u2_Display/n2937 ;
  wire \u2_Display/n2938 ;
  wire \u2_Display/n2939 ;
  wire \u2_Display/n2940 ;
  wire \u2_Display/n2941 ;
  wire \u2_Display/n2942 ;
  wire \u2_Display/n2943 ;
  wire \u2_Display/n2946 ;
  wire \u2_Display/n2947 ;
  wire \u2_Display/n2948 ;
  wire \u2_Display/n2949 ;
  wire \u2_Display/n2950 ;
  wire \u2_Display/n2951 ;
  wire \u2_Display/n2952 ;
  wire \u2_Display/n2953 ;
  wire \u2_Display/n2954 ;
  wire \u2_Display/n2955 ;
  wire \u2_Display/n2956 ;
  wire \u2_Display/n2957 ;
  wire \u2_Display/n2958 ;
  wire \u2_Display/n2959 ;
  wire \u2_Display/n2960 ;
  wire \u2_Display/n2961 ;
  wire \u2_Display/n2962 ;
  wire \u2_Display/n2963 ;
  wire \u2_Display/n2964 ;
  wire \u2_Display/n2965 ;
  wire \u2_Display/n2966 ;
  wire \u2_Display/n2967 ;
  wire \u2_Display/n2968 ;
  wire \u2_Display/n2969 ;
  wire \u2_Display/n2970 ;
  wire \u2_Display/n2971 ;
  wire \u2_Display/n2972 ;
  wire \u2_Display/n2973 ;
  wire \u2_Display/n2974 ;
  wire \u2_Display/n2975 ;
  wire \u2_Display/n2976 ;
  wire \u2_Display/n2977 ;
  wire \u2_Display/n2978 ;
  wire \u2_Display/n2981 ;
  wire \u2_Display/n2982 ;
  wire \u2_Display/n2983 ;
  wire \u2_Display/n2984 ;
  wire \u2_Display/n2985 ;
  wire \u2_Display/n2986 ;
  wire \u2_Display/n2987 ;
  wire \u2_Display/n2988 ;
  wire \u2_Display/n2989 ;
  wire \u2_Display/n2990 ;
  wire \u2_Display/n2991 ;
  wire \u2_Display/n2992 ;
  wire \u2_Display/n2993 ;
  wire \u2_Display/n2994 ;
  wire \u2_Display/n2995 ;
  wire \u2_Display/n2996 ;
  wire \u2_Display/n2997 ;
  wire \u2_Display/n2998 ;
  wire \u2_Display/n2999 ;
  wire \u2_Display/n3000 ;
  wire \u2_Display/n3001 ;
  wire \u2_Display/n3002 ;
  wire \u2_Display/n3003 ;
  wire \u2_Display/n3004 ;
  wire \u2_Display/n3005 ;
  wire \u2_Display/n3006 ;
  wire \u2_Display/n3007 ;
  wire \u2_Display/n3008 ;
  wire \u2_Display/n3009 ;
  wire \u2_Display/n3010 ;
  wire \u2_Display/n3011 ;
  wire \u2_Display/n3012 ;
  wire \u2_Display/n3013 ;
  wire \u2_Display/n3016 ;
  wire \u2_Display/n3017 ;
  wire \u2_Display/n3018 ;
  wire \u2_Display/n3019 ;
  wire \u2_Display/n3020 ;
  wire \u2_Display/n3021 ;
  wire \u2_Display/n3022 ;
  wire \u2_Display/n3023 ;
  wire \u2_Display/n3024 ;
  wire \u2_Display/n3025 ;
  wire \u2_Display/n3026 ;
  wire \u2_Display/n3027 ;
  wire \u2_Display/n3028 ;
  wire \u2_Display/n3029 ;
  wire \u2_Display/n3030 ;
  wire \u2_Display/n3031 ;
  wire \u2_Display/n3032 ;
  wire \u2_Display/n3033 ;
  wire \u2_Display/n3034 ;
  wire \u2_Display/n3035 ;
  wire \u2_Display/n3036 ;
  wire \u2_Display/n3037 ;
  wire \u2_Display/n3038 ;
  wire \u2_Display/n3039 ;
  wire \u2_Display/n3040 ;
  wire \u2_Display/n3041 ;
  wire \u2_Display/n3042 ;
  wire \u2_Display/n3043 ;
  wire \u2_Display/n3044 ;
  wire \u2_Display/n3045 ;
  wire \u2_Display/n3046 ;
  wire \u2_Display/n3047 ;
  wire \u2_Display/n3048 ;
  wire \u2_Display/n3051 ;
  wire \u2_Display/n3052 ;
  wire \u2_Display/n3053 ;
  wire \u2_Display/n3054 ;
  wire \u2_Display/n3055 ;
  wire \u2_Display/n3056 ;
  wire \u2_Display/n3057 ;
  wire \u2_Display/n3058 ;
  wire \u2_Display/n3059 ;
  wire \u2_Display/n3060 ;
  wire \u2_Display/n3061 ;
  wire \u2_Display/n3062 ;
  wire \u2_Display/n3063 ;
  wire \u2_Display/n3064 ;
  wire \u2_Display/n3065 ;
  wire \u2_Display/n3066 ;
  wire \u2_Display/n3067 ;
  wire \u2_Display/n3068 ;
  wire \u2_Display/n3069 ;
  wire \u2_Display/n3070 ;
  wire \u2_Display/n3071 ;
  wire \u2_Display/n3072 ;
  wire \u2_Display/n3073 ;
  wire \u2_Display/n3074 ;
  wire \u2_Display/n3075 ;
  wire \u2_Display/n3076 ;
  wire \u2_Display/n3077 ;
  wire \u2_Display/n3078 ;
  wire \u2_Display/n3079 ;
  wire \u2_Display/n3080 ;
  wire \u2_Display/n3081 ;
  wire \u2_Display/n3082 ;
  wire \u2_Display/n3083 ;
  wire \u2_Display/n3086 ;
  wire \u2_Display/n3087 ;
  wire \u2_Display/n3088 ;
  wire \u2_Display/n3089 ;
  wire \u2_Display/n3090 ;
  wire \u2_Display/n3091 ;
  wire \u2_Display/n3092 ;
  wire \u2_Display/n3093 ;
  wire \u2_Display/n3094 ;
  wire \u2_Display/n3095 ;
  wire \u2_Display/n3096 ;
  wire \u2_Display/n3097 ;
  wire \u2_Display/n3098 ;
  wire \u2_Display/n3099 ;
  wire \u2_Display/n3100 ;
  wire \u2_Display/n3101 ;
  wire \u2_Display/n3102 ;
  wire \u2_Display/n3103 ;
  wire \u2_Display/n3104 ;
  wire \u2_Display/n3105 ;
  wire \u2_Display/n3106 ;
  wire \u2_Display/n3107 ;
  wire \u2_Display/n3108 ;
  wire \u2_Display/n3109 ;
  wire \u2_Display/n3110 ;
  wire \u2_Display/n3111 ;
  wire \u2_Display/n3112 ;
  wire \u2_Display/n3113 ;
  wire \u2_Display/n3114 ;
  wire \u2_Display/n3115 ;
  wire \u2_Display/n3116 ;
  wire \u2_Display/n3117 ;
  wire \u2_Display/n3118 ;
  wire \u2_Display/n3121 ;
  wire \u2_Display/n3122 ;
  wire \u2_Display/n3123 ;
  wire \u2_Display/n3124 ;
  wire \u2_Display/n3125 ;
  wire \u2_Display/n3126 ;
  wire \u2_Display/n3127 ;
  wire \u2_Display/n3128 ;
  wire \u2_Display/n3129 ;
  wire \u2_Display/n3130 ;
  wire \u2_Display/n3131 ;
  wire \u2_Display/n3132 ;
  wire \u2_Display/n3133 ;
  wire \u2_Display/n3134 ;
  wire \u2_Display/n3135 ;
  wire \u2_Display/n3136 ;
  wire \u2_Display/n3137 ;
  wire \u2_Display/n3138 ;
  wire \u2_Display/n3139 ;
  wire \u2_Display/n3140 ;
  wire \u2_Display/n3141 ;
  wire \u2_Display/n3142 ;
  wire \u2_Display/n3143 ;
  wire \u2_Display/n3144 ;
  wire \u2_Display/n3145 ;
  wire \u2_Display/n3146 ;
  wire \u2_Display/n3147 ;
  wire \u2_Display/n3148 ;
  wire \u2_Display/n3149 ;
  wire \u2_Display/n3150 ;
  wire \u2_Display/n3151 ;
  wire \u2_Display/n3152 ;
  wire \u2_Display/n3153 ;
  wire \u2_Display/n3156 ;
  wire \u2_Display/n3157 ;
  wire \u2_Display/n3158 ;
  wire \u2_Display/n3159 ;
  wire \u2_Display/n3160 ;
  wire \u2_Display/n3161 ;
  wire \u2_Display/n3162 ;
  wire \u2_Display/n3163 ;
  wire \u2_Display/n3164 ;
  wire \u2_Display/n3165 ;
  wire \u2_Display/n3166 ;
  wire \u2_Display/n3167 ;
  wire \u2_Display/n3168 ;
  wire \u2_Display/n3169 ;
  wire \u2_Display/n3170 ;
  wire \u2_Display/n3171 ;
  wire \u2_Display/n3172 ;
  wire \u2_Display/n3173 ;
  wire \u2_Display/n3174 ;
  wire \u2_Display/n3175 ;
  wire \u2_Display/n3176 ;
  wire \u2_Display/n3177 ;
  wire \u2_Display/n3178 ;
  wire \u2_Display/n3179 ;
  wire \u2_Display/n3180 ;
  wire \u2_Display/n3181 ;
  wire \u2_Display/n3182 ;
  wire \u2_Display/n3183 ;
  wire \u2_Display/n3184 ;
  wire \u2_Display/n3185 ;
  wire \u2_Display/n3186 ;
  wire \u2_Display/n3187 ;
  wire \u2_Display/n3188 ;
  wire \u2_Display/n3191 ;
  wire \u2_Display/n3192 ;
  wire \u2_Display/n3193 ;
  wire \u2_Display/n3194 ;
  wire \u2_Display/n3195 ;
  wire \u2_Display/n3196 ;
  wire \u2_Display/n3197 ;
  wire \u2_Display/n3198 ;
  wire \u2_Display/n3199 ;
  wire \u2_Display/n3200 ;
  wire \u2_Display/n3201 ;
  wire \u2_Display/n3202 ;
  wire \u2_Display/n3203 ;
  wire \u2_Display/n3204 ;
  wire \u2_Display/n3205 ;
  wire \u2_Display/n3206 ;
  wire \u2_Display/n3207 ;
  wire \u2_Display/n3208 ;
  wire \u2_Display/n3209 ;
  wire \u2_Display/n3210 ;
  wire \u2_Display/n3211 ;
  wire \u2_Display/n3212 ;
  wire \u2_Display/n3213 ;
  wire \u2_Display/n3214 ;
  wire \u2_Display/n3215 ;
  wire \u2_Display/n3216 ;
  wire \u2_Display/n3217 ;
  wire \u2_Display/n3218 ;
  wire \u2_Display/n3219 ;
  wire \u2_Display/n3220 ;
  wire \u2_Display/n3221 ;
  wire \u2_Display/n3222 ;
  wire \u2_Display/n3223 ;
  wire \u2_Display/n3226 ;
  wire \u2_Display/n3227 ;
  wire \u2_Display/n3228 ;
  wire \u2_Display/n3229 ;
  wire \u2_Display/n3230 ;
  wire \u2_Display/n3231 ;
  wire \u2_Display/n3232 ;
  wire \u2_Display/n3233 ;
  wire \u2_Display/n3234 ;
  wire \u2_Display/n3235 ;
  wire \u2_Display/n3236 ;
  wire \u2_Display/n3237 ;
  wire \u2_Display/n3238 ;
  wire \u2_Display/n3239 ;
  wire \u2_Display/n3240 ;
  wire \u2_Display/n3241 ;
  wire \u2_Display/n3242 ;
  wire \u2_Display/n3243 ;
  wire \u2_Display/n3244 ;
  wire \u2_Display/n3245 ;
  wire \u2_Display/n3246 ;
  wire \u2_Display/n3247 ;
  wire \u2_Display/n3248 ;
  wire \u2_Display/n3249 ;
  wire \u2_Display/n3250 ;
  wire \u2_Display/n3251 ;
  wire \u2_Display/n3252 ;
  wire \u2_Display/n3253 ;
  wire \u2_Display/n3254 ;
  wire \u2_Display/n3255 ;
  wire \u2_Display/n3256 ;
  wire \u2_Display/n3257 ;
  wire \u2_Display/n3258 ;
  wire \u2_Display/n3261 ;
  wire \u2_Display/n3262 ;
  wire \u2_Display/n3263 ;
  wire \u2_Display/n3264 ;
  wire \u2_Display/n3265 ;
  wire \u2_Display/n3266 ;
  wire \u2_Display/n3267 ;
  wire \u2_Display/n3268 ;
  wire \u2_Display/n3269 ;
  wire \u2_Display/n3270 ;
  wire \u2_Display/n3271 ;
  wire \u2_Display/n3272 ;
  wire \u2_Display/n3273 ;
  wire \u2_Display/n3274 ;
  wire \u2_Display/n3275 ;
  wire \u2_Display/n3276 ;
  wire \u2_Display/n3277 ;
  wire \u2_Display/n3278 ;
  wire \u2_Display/n3279 ;
  wire \u2_Display/n3280 ;
  wire \u2_Display/n3281 ;
  wire \u2_Display/n3282 ;
  wire \u2_Display/n3283 ;
  wire \u2_Display/n3284 ;
  wire \u2_Display/n3285 ;
  wire \u2_Display/n3286 ;
  wire \u2_Display/n3287 ;
  wire \u2_Display/n3288 ;
  wire \u2_Display/n3289 ;
  wire \u2_Display/n3290 ;
  wire \u2_Display/n3291 ;
  wire \u2_Display/n3292 ;
  wire \u2_Display/n3293 ;
  wire \u2_Display/n3296 ;
  wire \u2_Display/n3297 ;
  wire \u2_Display/n3298 ;
  wire \u2_Display/n3299 ;
  wire \u2_Display/n3300 ;
  wire \u2_Display/n3301 ;
  wire \u2_Display/n3302 ;
  wire \u2_Display/n3303 ;
  wire \u2_Display/n3304 ;
  wire \u2_Display/n3305 ;
  wire \u2_Display/n3306 ;
  wire \u2_Display/n3307 ;
  wire \u2_Display/n3308 ;
  wire \u2_Display/n3309 ;
  wire \u2_Display/n3310 ;
  wire \u2_Display/n3311 ;
  wire \u2_Display/n3312 ;
  wire \u2_Display/n3313 ;
  wire \u2_Display/n3314 ;
  wire \u2_Display/n3315 ;
  wire \u2_Display/n3316 ;
  wire \u2_Display/n3317 ;
  wire \u2_Display/n3318 ;
  wire \u2_Display/n3319 ;
  wire \u2_Display/n3320 ;
  wire \u2_Display/n3321 ;
  wire \u2_Display/n3322 ;
  wire \u2_Display/n3323 ;
  wire \u2_Display/n3324 ;
  wire \u2_Display/n3325 ;
  wire \u2_Display/n3326 ;
  wire \u2_Display/n3327 ;
  wire \u2_Display/n3328 ;
  wire \u2_Display/n3331 ;
  wire \u2_Display/n3332 ;
  wire \u2_Display/n3333 ;
  wire \u2_Display/n3334 ;
  wire \u2_Display/n3335 ;
  wire \u2_Display/n3336 ;
  wire \u2_Display/n3337 ;
  wire \u2_Display/n3338 ;
  wire \u2_Display/n3339 ;
  wire \u2_Display/n3340 ;
  wire \u2_Display/n3341 ;
  wire \u2_Display/n3342 ;
  wire \u2_Display/n3343 ;
  wire \u2_Display/n3344 ;
  wire \u2_Display/n3345 ;
  wire \u2_Display/n3346 ;
  wire \u2_Display/n3347 ;
  wire \u2_Display/n3348 ;
  wire \u2_Display/n3349 ;
  wire \u2_Display/n3350 ;
  wire \u2_Display/n3351 ;
  wire \u2_Display/n3352 ;
  wire \u2_Display/n3353 ;
  wire \u2_Display/n3354 ;
  wire \u2_Display/n3355 ;
  wire \u2_Display/n3356 ;
  wire \u2_Display/n3357 ;
  wire \u2_Display/n3358 ;
  wire \u2_Display/n3359 ;
  wire \u2_Display/n3360 ;
  wire \u2_Display/n3361 ;
  wire \u2_Display/n3362 ;
  wire \u2_Display/n3363 ;
  wire \u2_Display/n3366 ;
  wire \u2_Display/n3367 ;
  wire \u2_Display/n3368 ;
  wire \u2_Display/n3369 ;
  wire \u2_Display/n3370 ;
  wire \u2_Display/n3371 ;
  wire \u2_Display/n3372 ;
  wire \u2_Display/n3373 ;
  wire \u2_Display/n3374 ;
  wire \u2_Display/n3375 ;
  wire \u2_Display/n3376 ;
  wire \u2_Display/n3377 ;
  wire \u2_Display/n3378 ;
  wire \u2_Display/n3379 ;
  wire \u2_Display/n3380 ;
  wire \u2_Display/n3381 ;
  wire \u2_Display/n3382 ;
  wire \u2_Display/n3383 ;
  wire \u2_Display/n3384 ;
  wire \u2_Display/n3385 ;
  wire \u2_Display/n3386 ;
  wire \u2_Display/n3387 ;
  wire \u2_Display/n3388 ;
  wire \u2_Display/n3389 ;
  wire \u2_Display/n3390 ;
  wire \u2_Display/n3391 ;
  wire \u2_Display/n3392 ;
  wire \u2_Display/n3393 ;
  wire \u2_Display/n3394 ;
  wire \u2_Display/n3395 ;
  wire \u2_Display/n3396 ;
  wire \u2_Display/n3397 ;
  wire \u2_Display/n3398 ;
  wire \u2_Display/n3401 ;
  wire \u2_Display/n3402 ;
  wire \u2_Display/n3403 ;
  wire \u2_Display/n3404 ;
  wire \u2_Display/n3405 ;
  wire \u2_Display/n3406 ;
  wire \u2_Display/n3407 ;
  wire \u2_Display/n3408 ;
  wire \u2_Display/n3409 ;
  wire \u2_Display/n3410 ;
  wire \u2_Display/n3411 ;
  wire \u2_Display/n3412 ;
  wire \u2_Display/n3413 ;
  wire \u2_Display/n3414 ;
  wire \u2_Display/n3415 ;
  wire \u2_Display/n3416 ;
  wire \u2_Display/n3417 ;
  wire \u2_Display/n3418 ;
  wire \u2_Display/n3419 ;
  wire \u2_Display/n3420 ;
  wire \u2_Display/n3421 ;
  wire \u2_Display/n3422 ;
  wire \u2_Display/n3423 ;
  wire \u2_Display/n3424 ;
  wire \u2_Display/n3425 ;
  wire \u2_Display/n3426 ;
  wire \u2_Display/n3427 ;
  wire \u2_Display/n3428 ;
  wire \u2_Display/n3429 ;
  wire \u2_Display/n3430 ;
  wire \u2_Display/n3431 ;
  wire \u2_Display/n3432 ;
  wire \u2_Display/n3433 ;
  wire \u2_Display/n35 ;
  wire \u2_Display/n3786 ;
  wire \u2_Display/n3789 ;
  wire \u2_Display/n3790 ;
  wire \u2_Display/n3791 ;
  wire \u2_Display/n3792 ;
  wire \u2_Display/n3793 ;
  wire \u2_Display/n3794 ;
  wire \u2_Display/n3795 ;
  wire \u2_Display/n3796 ;
  wire \u2_Display/n3797 ;
  wire \u2_Display/n3798 ;
  wire \u2_Display/n3799 ;
  wire \u2_Display/n3800 ;
  wire \u2_Display/n3801 ;
  wire \u2_Display/n3802 ;
  wire \u2_Display/n3803 ;
  wire \u2_Display/n3804 ;
  wire \u2_Display/n3805 ;
  wire \u2_Display/n3806 ;
  wire \u2_Display/n3807 ;
  wire \u2_Display/n3808 ;
  wire \u2_Display/n3809 ;
  wire \u2_Display/n3810 ;
  wire \u2_Display/n3811 ;
  wire \u2_Display/n3812 ;
  wire \u2_Display/n3813 ;
  wire \u2_Display/n3814 ;
  wire \u2_Display/n3815 ;
  wire \u2_Display/n3816 ;
  wire \u2_Display/n3817 ;
  wire \u2_Display/n3818 ;
  wire \u2_Display/n3819 ;
  wire \u2_Display/n3820 ;
  wire \u2_Display/n3821 ;
  wire \u2_Display/n3824 ;
  wire \u2_Display/n3825 ;
  wire \u2_Display/n3826 ;
  wire \u2_Display/n3827 ;
  wire \u2_Display/n3828 ;
  wire \u2_Display/n3829 ;
  wire \u2_Display/n3830 ;
  wire \u2_Display/n3831 ;
  wire \u2_Display/n3832 ;
  wire \u2_Display/n3833 ;
  wire \u2_Display/n3834 ;
  wire \u2_Display/n3835 ;
  wire \u2_Display/n3836 ;
  wire \u2_Display/n3837 ;
  wire \u2_Display/n3838 ;
  wire \u2_Display/n3839 ;
  wire \u2_Display/n3840 ;
  wire \u2_Display/n3841 ;
  wire \u2_Display/n3842 ;
  wire \u2_Display/n3843 ;
  wire \u2_Display/n3844 ;
  wire \u2_Display/n3845 ;
  wire \u2_Display/n3846 ;
  wire \u2_Display/n3847 ;
  wire \u2_Display/n3848 ;
  wire \u2_Display/n3849 ;
  wire \u2_Display/n3850 ;
  wire \u2_Display/n3851 ;
  wire \u2_Display/n3852 ;
  wire \u2_Display/n3853 ;
  wire \u2_Display/n3854 ;
  wire \u2_Display/n3855 ;
  wire \u2_Display/n3856 ;
  wire \u2_Display/n3859 ;
  wire \u2_Display/n3860 ;
  wire \u2_Display/n3861 ;
  wire \u2_Display/n3862 ;
  wire \u2_Display/n3863 ;
  wire \u2_Display/n3864 ;
  wire \u2_Display/n3865 ;
  wire \u2_Display/n3866 ;
  wire \u2_Display/n3867 ;
  wire \u2_Display/n3868 ;
  wire \u2_Display/n3869 ;
  wire \u2_Display/n3870 ;
  wire \u2_Display/n3871 ;
  wire \u2_Display/n3872 ;
  wire \u2_Display/n3873 ;
  wire \u2_Display/n3874 ;
  wire \u2_Display/n3875 ;
  wire \u2_Display/n3876 ;
  wire \u2_Display/n3877 ;
  wire \u2_Display/n3878 ;
  wire \u2_Display/n3879 ;
  wire \u2_Display/n3880 ;
  wire \u2_Display/n3881 ;
  wire \u2_Display/n3882 ;
  wire \u2_Display/n3883 ;
  wire \u2_Display/n3884 ;
  wire \u2_Display/n3885 ;
  wire \u2_Display/n3886 ;
  wire \u2_Display/n3887 ;
  wire \u2_Display/n3888 ;
  wire \u2_Display/n3889 ;
  wire \u2_Display/n3890 ;
  wire \u2_Display/n3891 ;
  wire \u2_Display/n3894 ;
  wire \u2_Display/n3895 ;
  wire \u2_Display/n3896 ;
  wire \u2_Display/n3897 ;
  wire \u2_Display/n3898 ;
  wire \u2_Display/n3899 ;
  wire \u2_Display/n3900 ;
  wire \u2_Display/n3901 ;
  wire \u2_Display/n3902 ;
  wire \u2_Display/n3903 ;
  wire \u2_Display/n3904 ;
  wire \u2_Display/n3905 ;
  wire \u2_Display/n3906 ;
  wire \u2_Display/n3907 ;
  wire \u2_Display/n3908 ;
  wire \u2_Display/n3909 ;
  wire \u2_Display/n3910 ;
  wire \u2_Display/n3911 ;
  wire \u2_Display/n3912 ;
  wire \u2_Display/n3913 ;
  wire \u2_Display/n3914 ;
  wire \u2_Display/n3915 ;
  wire \u2_Display/n3916 ;
  wire \u2_Display/n3917 ;
  wire \u2_Display/n3918 ;
  wire \u2_Display/n3919 ;
  wire \u2_Display/n3920 ;
  wire \u2_Display/n3921 ;
  wire \u2_Display/n3922 ;
  wire \u2_Display/n3923 ;
  wire \u2_Display/n3924 ;
  wire \u2_Display/n3925 ;
  wire \u2_Display/n3926 ;
  wire \u2_Display/n3929 ;
  wire \u2_Display/n3930 ;
  wire \u2_Display/n3931 ;
  wire \u2_Display/n3932 ;
  wire \u2_Display/n3933 ;
  wire \u2_Display/n3934 ;
  wire \u2_Display/n3935 ;
  wire \u2_Display/n3936 ;
  wire \u2_Display/n3937 ;
  wire \u2_Display/n3938 ;
  wire \u2_Display/n3939 ;
  wire \u2_Display/n3940 ;
  wire \u2_Display/n3941 ;
  wire \u2_Display/n3942 ;
  wire \u2_Display/n3943 ;
  wire \u2_Display/n3944 ;
  wire \u2_Display/n3945 ;
  wire \u2_Display/n3946 ;
  wire \u2_Display/n3947 ;
  wire \u2_Display/n3948 ;
  wire \u2_Display/n3949 ;
  wire \u2_Display/n3950 ;
  wire \u2_Display/n3951 ;
  wire \u2_Display/n3952 ;
  wire \u2_Display/n3953 ;
  wire \u2_Display/n3954 ;
  wire \u2_Display/n3955 ;
  wire \u2_Display/n3956 ;
  wire \u2_Display/n3957 ;
  wire \u2_Display/n3958 ;
  wire \u2_Display/n3959 ;
  wire \u2_Display/n3960 ;
  wire \u2_Display/n3961 ;
  wire \u2_Display/n3964 ;
  wire \u2_Display/n3965 ;
  wire \u2_Display/n3966 ;
  wire \u2_Display/n3967 ;
  wire \u2_Display/n3968 ;
  wire \u2_Display/n3969 ;
  wire \u2_Display/n3970 ;
  wire \u2_Display/n3971 ;
  wire \u2_Display/n3972 ;
  wire \u2_Display/n3973 ;
  wire \u2_Display/n3974 ;
  wire \u2_Display/n3975 ;
  wire \u2_Display/n3976 ;
  wire \u2_Display/n3977 ;
  wire \u2_Display/n3978 ;
  wire \u2_Display/n3979 ;
  wire \u2_Display/n3980 ;
  wire \u2_Display/n3981 ;
  wire \u2_Display/n3982 ;
  wire \u2_Display/n3983 ;
  wire \u2_Display/n3984 ;
  wire \u2_Display/n3985 ;
  wire \u2_Display/n3986 ;
  wire \u2_Display/n3987 ;
  wire \u2_Display/n3988 ;
  wire \u2_Display/n3989 ;
  wire \u2_Display/n3990 ;
  wire \u2_Display/n3991 ;
  wire \u2_Display/n3992 ;
  wire \u2_Display/n3993 ;
  wire \u2_Display/n3994 ;
  wire \u2_Display/n3995 ;
  wire \u2_Display/n3996 ;
  wire \u2_Display/n3999 ;
  wire \u2_Display/n4000 ;
  wire \u2_Display/n4001 ;
  wire \u2_Display/n4002 ;
  wire \u2_Display/n4003 ;
  wire \u2_Display/n4004 ;
  wire \u2_Display/n4005 ;
  wire \u2_Display/n4006 ;
  wire \u2_Display/n4007 ;
  wire \u2_Display/n4008 ;
  wire \u2_Display/n4009 ;
  wire \u2_Display/n4010 ;
  wire \u2_Display/n4011 ;
  wire \u2_Display/n4012 ;
  wire \u2_Display/n4013 ;
  wire \u2_Display/n4014 ;
  wire \u2_Display/n4015 ;
  wire \u2_Display/n4016 ;
  wire \u2_Display/n4017 ;
  wire \u2_Display/n4018 ;
  wire \u2_Display/n4019 ;
  wire \u2_Display/n4020 ;
  wire \u2_Display/n4021 ;
  wire \u2_Display/n4022 ;
  wire \u2_Display/n4023 ;
  wire \u2_Display/n4024 ;
  wire \u2_Display/n4025 ;
  wire \u2_Display/n4026 ;
  wire \u2_Display/n4027 ;
  wire \u2_Display/n4028 ;
  wire \u2_Display/n4029 ;
  wire \u2_Display/n4030 ;
  wire \u2_Display/n4031 ;
  wire \u2_Display/n4034 ;
  wire \u2_Display/n4035 ;
  wire \u2_Display/n4036 ;
  wire \u2_Display/n4037 ;
  wire \u2_Display/n4038 ;
  wire \u2_Display/n4039 ;
  wire \u2_Display/n4040 ;
  wire \u2_Display/n4041 ;
  wire \u2_Display/n4042 ;
  wire \u2_Display/n4043 ;
  wire \u2_Display/n4044 ;
  wire \u2_Display/n4045 ;
  wire \u2_Display/n4046 ;
  wire \u2_Display/n4047 ;
  wire \u2_Display/n4048 ;
  wire \u2_Display/n4049 ;
  wire \u2_Display/n4050 ;
  wire \u2_Display/n4051 ;
  wire \u2_Display/n4052 ;
  wire \u2_Display/n4053 ;
  wire \u2_Display/n4054 ;
  wire \u2_Display/n4055 ;
  wire \u2_Display/n4056 ;
  wire \u2_Display/n4057 ;
  wire \u2_Display/n4058 ;
  wire \u2_Display/n4059 ;
  wire \u2_Display/n4060 ;
  wire \u2_Display/n4061 ;
  wire \u2_Display/n4062 ;
  wire \u2_Display/n4063 ;
  wire \u2_Display/n4064 ;
  wire \u2_Display/n4065 ;
  wire \u2_Display/n4066 ;
  wire \u2_Display/n4069 ;
  wire \u2_Display/n4070 ;
  wire \u2_Display/n4071 ;
  wire \u2_Display/n4072 ;
  wire \u2_Display/n4073 ;
  wire \u2_Display/n4074 ;
  wire \u2_Display/n4075 ;
  wire \u2_Display/n4076 ;
  wire \u2_Display/n4077 ;
  wire \u2_Display/n4078 ;
  wire \u2_Display/n4079 ;
  wire \u2_Display/n4080 ;
  wire \u2_Display/n4081 ;
  wire \u2_Display/n4082 ;
  wire \u2_Display/n4083 ;
  wire \u2_Display/n4084 ;
  wire \u2_Display/n4085 ;
  wire \u2_Display/n4086 ;
  wire \u2_Display/n4087 ;
  wire \u2_Display/n4088 ;
  wire \u2_Display/n4089 ;
  wire \u2_Display/n4090 ;
  wire \u2_Display/n4091 ;
  wire \u2_Display/n4092 ;
  wire \u2_Display/n4093 ;
  wire \u2_Display/n4094 ;
  wire \u2_Display/n4095 ;
  wire \u2_Display/n4096 ;
  wire \u2_Display/n4097 ;
  wire \u2_Display/n4098 ;
  wire \u2_Display/n4099 ;
  wire \u2_Display/n4100 ;
  wire \u2_Display/n4101 ;
  wire \u2_Display/n4104 ;
  wire \u2_Display/n4105 ;
  wire \u2_Display/n4106 ;
  wire \u2_Display/n4107 ;
  wire \u2_Display/n4108 ;
  wire \u2_Display/n4109 ;
  wire \u2_Display/n4110 ;
  wire \u2_Display/n4111 ;
  wire \u2_Display/n4112 ;
  wire \u2_Display/n4113 ;
  wire \u2_Display/n4114 ;
  wire \u2_Display/n4115 ;
  wire \u2_Display/n4116 ;
  wire \u2_Display/n4117 ;
  wire \u2_Display/n4118 ;
  wire \u2_Display/n4119 ;
  wire \u2_Display/n4120 ;
  wire \u2_Display/n4121 ;
  wire \u2_Display/n4122 ;
  wire \u2_Display/n4123 ;
  wire \u2_Display/n4124 ;
  wire \u2_Display/n4125 ;
  wire \u2_Display/n4126 ;
  wire \u2_Display/n4127 ;
  wire \u2_Display/n4128 ;
  wire \u2_Display/n4129 ;
  wire \u2_Display/n4130 ;
  wire \u2_Display/n4131 ;
  wire \u2_Display/n4132 ;
  wire \u2_Display/n4133 ;
  wire \u2_Display/n4134 ;
  wire \u2_Display/n4135 ;
  wire \u2_Display/n4136 ;
  wire \u2_Display/n4139 ;
  wire \u2_Display/n4140 ;
  wire \u2_Display/n4141 ;
  wire \u2_Display/n4142 ;
  wire \u2_Display/n4143 ;
  wire \u2_Display/n4144 ;
  wire \u2_Display/n4145 ;
  wire \u2_Display/n4146 ;
  wire \u2_Display/n4147 ;
  wire \u2_Display/n4148 ;
  wire \u2_Display/n4149 ;
  wire \u2_Display/n4150 ;
  wire \u2_Display/n4151 ;
  wire \u2_Display/n4152 ;
  wire \u2_Display/n4153 ;
  wire \u2_Display/n4154 ;
  wire \u2_Display/n4155 ;
  wire \u2_Display/n4156 ;
  wire \u2_Display/n4157 ;
  wire \u2_Display/n4158 ;
  wire \u2_Display/n4159 ;
  wire \u2_Display/n4160 ;
  wire \u2_Display/n4161 ;
  wire \u2_Display/n4162 ;
  wire \u2_Display/n4163 ;
  wire \u2_Display/n4164 ;
  wire \u2_Display/n4165 ;
  wire \u2_Display/n4166 ;
  wire \u2_Display/n4167 ;
  wire \u2_Display/n4168 ;
  wire \u2_Display/n4169 ;
  wire \u2_Display/n417 ;
  wire \u2_Display/n4170 ;
  wire \u2_Display/n4171 ;
  wire \u2_Display/n4174 ;
  wire \u2_Display/n4175 ;
  wire \u2_Display/n4176 ;
  wire \u2_Display/n4177 ;
  wire \u2_Display/n4178 ;
  wire \u2_Display/n4179 ;
  wire \u2_Display/n4180 ;
  wire \u2_Display/n4181 ;
  wire \u2_Display/n4182 ;
  wire \u2_Display/n4183 ;
  wire \u2_Display/n4184 ;
  wire \u2_Display/n4185 ;
  wire \u2_Display/n4186 ;
  wire \u2_Display/n4187 ;
  wire \u2_Display/n4188 ;
  wire \u2_Display/n4189 ;
  wire \u2_Display/n4190 ;
  wire \u2_Display/n4191 ;
  wire \u2_Display/n4192 ;
  wire \u2_Display/n4193 ;
  wire \u2_Display/n4194 ;
  wire \u2_Display/n4195 ;
  wire \u2_Display/n4196 ;
  wire \u2_Display/n4197 ;
  wire \u2_Display/n4198 ;
  wire \u2_Display/n4199 ;
  wire \u2_Display/n420 ;
  wire \u2_Display/n4200 ;
  wire \u2_Display/n4201 ;
  wire \u2_Display/n4202 ;
  wire \u2_Display/n4203 ;
  wire \u2_Display/n4204 ;
  wire \u2_Display/n4205 ;
  wire \u2_Display/n4206 ;
  wire \u2_Display/n4209 ;
  wire \u2_Display/n421 ;
  wire \u2_Display/n4210 ;
  wire \u2_Display/n4211 ;
  wire \u2_Display/n4212 ;
  wire \u2_Display/n4213 ;
  wire \u2_Display/n4214 ;
  wire \u2_Display/n4215 ;
  wire \u2_Display/n4216 ;
  wire \u2_Display/n4217 ;
  wire \u2_Display/n4218 ;
  wire \u2_Display/n4219 ;
  wire \u2_Display/n422 ;
  wire \u2_Display/n4220 ;
  wire \u2_Display/n4221 ;
  wire \u2_Display/n4222 ;
  wire \u2_Display/n4223 ;
  wire \u2_Display/n4224 ;
  wire \u2_Display/n4225 ;
  wire \u2_Display/n4226 ;
  wire \u2_Display/n4227 ;
  wire \u2_Display/n4228 ;
  wire \u2_Display/n4229 ;
  wire \u2_Display/n423 ;
  wire \u2_Display/n4230 ;
  wire \u2_Display/n4231 ;
  wire \u2_Display/n4232 ;
  wire \u2_Display/n4233 ;
  wire \u2_Display/n4234 ;
  wire \u2_Display/n4235 ;
  wire \u2_Display/n4236 ;
  wire \u2_Display/n4237 ;
  wire \u2_Display/n4238 ;
  wire \u2_Display/n4239 ;
  wire \u2_Display/n424 ;
  wire \u2_Display/n4240 ;
  wire \u2_Display/n4241 ;
  wire \u2_Display/n4244 ;
  wire \u2_Display/n4245 ;
  wire \u2_Display/n4246 ;
  wire \u2_Display/n4247 ;
  wire \u2_Display/n4248 ;
  wire \u2_Display/n4249 ;
  wire \u2_Display/n425 ;
  wire \u2_Display/n4250 ;
  wire \u2_Display/n4251 ;
  wire \u2_Display/n4252 ;
  wire \u2_Display/n4253 ;
  wire \u2_Display/n4254 ;
  wire \u2_Display/n4255 ;
  wire \u2_Display/n4256 ;
  wire \u2_Display/n4257 ;
  wire \u2_Display/n4258 ;
  wire \u2_Display/n4259 ;
  wire \u2_Display/n426 ;
  wire \u2_Display/n4260 ;
  wire \u2_Display/n4261 ;
  wire \u2_Display/n4262 ;
  wire \u2_Display/n4263 ;
  wire \u2_Display/n4264 ;
  wire \u2_Display/n4265 ;
  wire \u2_Display/n4266 ;
  wire \u2_Display/n4267 ;
  wire \u2_Display/n4268 ;
  wire \u2_Display/n4269 ;
  wire \u2_Display/n427 ;
  wire \u2_Display/n4270 ;
  wire \u2_Display/n4271 ;
  wire \u2_Display/n4272 ;
  wire \u2_Display/n4273 ;
  wire \u2_Display/n4274 ;
  wire \u2_Display/n4275 ;
  wire \u2_Display/n4276 ;
  wire \u2_Display/n4279 ;
  wire \u2_Display/n428 ;
  wire \u2_Display/n4280 ;
  wire \u2_Display/n4281 ;
  wire \u2_Display/n4282 ;
  wire \u2_Display/n4283 ;
  wire \u2_Display/n4284 ;
  wire \u2_Display/n4285 ;
  wire \u2_Display/n4286 ;
  wire \u2_Display/n4287 ;
  wire \u2_Display/n4288 ;
  wire \u2_Display/n4289 ;
  wire \u2_Display/n429 ;
  wire \u2_Display/n4290 ;
  wire \u2_Display/n4291 ;
  wire \u2_Display/n4292 ;
  wire \u2_Display/n4293 ;
  wire \u2_Display/n4294 ;
  wire \u2_Display/n4295 ;
  wire \u2_Display/n4296 ;
  wire \u2_Display/n4297 ;
  wire \u2_Display/n4298 ;
  wire \u2_Display/n4299 ;
  wire \u2_Display/n430 ;
  wire \u2_Display/n4300 ;
  wire \u2_Display/n4301 ;
  wire \u2_Display/n4302 ;
  wire \u2_Display/n4303 ;
  wire \u2_Display/n4304 ;
  wire \u2_Display/n4305 ;
  wire \u2_Display/n4306 ;
  wire \u2_Display/n4307 ;
  wire \u2_Display/n4308 ;
  wire \u2_Display/n4309 ;
  wire \u2_Display/n431 ;
  wire \u2_Display/n4310 ;
  wire \u2_Display/n4311 ;
  wire \u2_Display/n4314 ;
  wire \u2_Display/n4315 ;
  wire \u2_Display/n4316 ;
  wire \u2_Display/n4317 ;
  wire \u2_Display/n4318 ;
  wire \u2_Display/n4319 ;
  wire \u2_Display/n432 ;
  wire \u2_Display/n4320 ;
  wire \u2_Display/n4321 ;
  wire \u2_Display/n4322 ;
  wire \u2_Display/n4323 ;
  wire \u2_Display/n4324 ;
  wire \u2_Display/n4325 ;
  wire \u2_Display/n4326 ;
  wire \u2_Display/n4327 ;
  wire \u2_Display/n4328 ;
  wire \u2_Display/n4329 ;
  wire \u2_Display/n433 ;
  wire \u2_Display/n4330 ;
  wire \u2_Display/n4331 ;
  wire \u2_Display/n4332 ;
  wire \u2_Display/n4333 ;
  wire \u2_Display/n4334 ;
  wire \u2_Display/n4335 ;
  wire \u2_Display/n4336 ;
  wire \u2_Display/n4337 ;
  wire \u2_Display/n4338 ;
  wire \u2_Display/n4339 ;
  wire \u2_Display/n434 ;
  wire \u2_Display/n4340 ;
  wire \u2_Display/n4341 ;
  wire \u2_Display/n4342 ;
  wire \u2_Display/n4343 ;
  wire \u2_Display/n4344 ;
  wire \u2_Display/n4345 ;
  wire \u2_Display/n4346 ;
  wire \u2_Display/n4349 ;
  wire \u2_Display/n435 ;
  wire \u2_Display/n4350 ;
  wire \u2_Display/n4351 ;
  wire \u2_Display/n4352 ;
  wire \u2_Display/n4353 ;
  wire \u2_Display/n4354 ;
  wire \u2_Display/n4355 ;
  wire \u2_Display/n4356 ;
  wire \u2_Display/n4357 ;
  wire \u2_Display/n4358 ;
  wire \u2_Display/n4359 ;
  wire \u2_Display/n436 ;
  wire \u2_Display/n4360 ;
  wire \u2_Display/n4361 ;
  wire \u2_Display/n4362 ;
  wire \u2_Display/n4363 ;
  wire \u2_Display/n4364 ;
  wire \u2_Display/n4365 ;
  wire \u2_Display/n4366 ;
  wire \u2_Display/n4367 ;
  wire \u2_Display/n4368 ;
  wire \u2_Display/n4369 ;
  wire \u2_Display/n437 ;
  wire \u2_Display/n4370 ;
  wire \u2_Display/n4371 ;
  wire \u2_Display/n4372 ;
  wire \u2_Display/n4373 ;
  wire \u2_Display/n4374 ;
  wire \u2_Display/n4375 ;
  wire \u2_Display/n4376 ;
  wire \u2_Display/n4377 ;
  wire \u2_Display/n4378 ;
  wire \u2_Display/n4379 ;
  wire \u2_Display/n438 ;
  wire \u2_Display/n4380 ;
  wire \u2_Display/n4381 ;
  wire \u2_Display/n4384 ;
  wire \u2_Display/n4385 ;
  wire \u2_Display/n4386 ;
  wire \u2_Display/n4387 ;
  wire \u2_Display/n4388 ;
  wire \u2_Display/n4389 ;
  wire \u2_Display/n439 ;
  wire \u2_Display/n4390 ;
  wire \u2_Display/n4391 ;
  wire \u2_Display/n4392 ;
  wire \u2_Display/n4393 ;
  wire \u2_Display/n4394 ;
  wire \u2_Display/n4395 ;
  wire \u2_Display/n4396 ;
  wire \u2_Display/n4397 ;
  wire \u2_Display/n4398 ;
  wire \u2_Display/n4399 ;
  wire \u2_Display/n44 ;
  wire \u2_Display/n440 ;
  wire \u2_Display/n4400 ;
  wire \u2_Display/n4401 ;
  wire \u2_Display/n4402 ;
  wire \u2_Display/n4403 ;
  wire \u2_Display/n4404 ;
  wire \u2_Display/n4405 ;
  wire \u2_Display/n4406 ;
  wire \u2_Display/n4407 ;
  wire \u2_Display/n4408 ;
  wire \u2_Display/n4409 ;
  wire \u2_Display/n441 ;
  wire \u2_Display/n4410 ;
  wire \u2_Display/n4411 ;
  wire \u2_Display/n4412 ;
  wire \u2_Display/n4413 ;
  wire \u2_Display/n4414 ;
  wire \u2_Display/n4415 ;
  wire \u2_Display/n4416 ;
  wire \u2_Display/n4419 ;
  wire \u2_Display/n442 ;
  wire \u2_Display/n4420 ;
  wire \u2_Display/n4421 ;
  wire \u2_Display/n4422 ;
  wire \u2_Display/n4423 ;
  wire \u2_Display/n4424 ;
  wire \u2_Display/n4425 ;
  wire \u2_Display/n4426 ;
  wire \u2_Display/n4427 ;
  wire \u2_Display/n4428 ;
  wire \u2_Display/n4429 ;
  wire \u2_Display/n443 ;
  wire \u2_Display/n4430 ;
  wire \u2_Display/n4431 ;
  wire \u2_Display/n4432 ;
  wire \u2_Display/n4433 ;
  wire \u2_Display/n4434 ;
  wire \u2_Display/n4435 ;
  wire \u2_Display/n4436 ;
  wire \u2_Display/n4437 ;
  wire \u2_Display/n4438 ;
  wire \u2_Display/n4439 ;
  wire \u2_Display/n444 ;
  wire \u2_Display/n4440 ;
  wire \u2_Display/n4441 ;
  wire \u2_Display/n4442 ;
  wire \u2_Display/n4443 ;
  wire \u2_Display/n4444 ;
  wire \u2_Display/n4445 ;
  wire \u2_Display/n4446 ;
  wire \u2_Display/n4447 ;
  wire \u2_Display/n4448 ;
  wire \u2_Display/n4449 ;
  wire \u2_Display/n445 ;
  wire \u2_Display/n4450 ;
  wire \u2_Display/n4451 ;
  wire \u2_Display/n4454 ;
  wire \u2_Display/n4455 ;
  wire \u2_Display/n4456 ;
  wire \u2_Display/n4457 ;
  wire \u2_Display/n4458 ;
  wire \u2_Display/n4459 ;
  wire \u2_Display/n446 ;
  wire \u2_Display/n4460 ;
  wire \u2_Display/n4461 ;
  wire \u2_Display/n4462 ;
  wire \u2_Display/n4463 ;
  wire \u2_Display/n4464 ;
  wire \u2_Display/n4465 ;
  wire \u2_Display/n4466 ;
  wire \u2_Display/n4467 ;
  wire \u2_Display/n4468 ;
  wire \u2_Display/n4469 ;
  wire \u2_Display/n447 ;
  wire \u2_Display/n4470 ;
  wire \u2_Display/n4471 ;
  wire \u2_Display/n4472 ;
  wire \u2_Display/n4473 ;
  wire \u2_Display/n4474 ;
  wire \u2_Display/n4475 ;
  wire \u2_Display/n4476 ;
  wire \u2_Display/n4477 ;
  wire \u2_Display/n4478 ;
  wire \u2_Display/n4479 ;
  wire \u2_Display/n448 ;
  wire \u2_Display/n4480 ;
  wire \u2_Display/n4481 ;
  wire \u2_Display/n4482 ;
  wire \u2_Display/n4483 ;
  wire \u2_Display/n4484 ;
  wire \u2_Display/n4485 ;
  wire \u2_Display/n4486 ;
  wire \u2_Display/n4489 ;
  wire \u2_Display/n449 ;
  wire \u2_Display/n4490 ;
  wire \u2_Display/n4491 ;
  wire \u2_Display/n4492 ;
  wire \u2_Display/n4493 ;
  wire \u2_Display/n4494 ;
  wire \u2_Display/n4495 ;
  wire \u2_Display/n4496 ;
  wire \u2_Display/n4497 ;
  wire \u2_Display/n4498 ;
  wire \u2_Display/n4499 ;
  wire \u2_Display/n45 ;
  wire \u2_Display/n450 ;
  wire \u2_Display/n4500 ;
  wire \u2_Display/n4501 ;
  wire \u2_Display/n4502 ;
  wire \u2_Display/n4503 ;
  wire \u2_Display/n4504 ;
  wire \u2_Display/n4505 ;
  wire \u2_Display/n4506 ;
  wire \u2_Display/n4507 ;
  wire \u2_Display/n4508 ;
  wire \u2_Display/n4509 ;
  wire \u2_Display/n451 ;
  wire \u2_Display/n4510 ;
  wire \u2_Display/n4511 ;
  wire \u2_Display/n4512 ;
  wire \u2_Display/n4513 ;
  wire \u2_Display/n4514 ;
  wire \u2_Display/n4515 ;
  wire \u2_Display/n4516 ;
  wire \u2_Display/n4517 ;
  wire \u2_Display/n4518 ;
  wire \u2_Display/n4519 ;
  wire \u2_Display/n452 ;
  wire \u2_Display/n4520 ;
  wire \u2_Display/n4521 ;
  wire \u2_Display/n4524 ;
  wire \u2_Display/n4525 ;
  wire \u2_Display/n4526 ;
  wire \u2_Display/n4527 ;
  wire \u2_Display/n4528 ;
  wire \u2_Display/n4529 ;
  wire \u2_Display/n4530 ;
  wire \u2_Display/n4531 ;
  wire \u2_Display/n4532 ;
  wire \u2_Display/n4533 ;
  wire \u2_Display/n4534 ;
  wire \u2_Display/n4535 ;
  wire \u2_Display/n4536 ;
  wire \u2_Display/n4537 ;
  wire \u2_Display/n4538 ;
  wire \u2_Display/n4539 ;
  wire \u2_Display/n4540 ;
  wire \u2_Display/n4541 ;
  wire \u2_Display/n4542 ;
  wire \u2_Display/n4543 ;
  wire \u2_Display/n4544 ;
  wire \u2_Display/n4545 ;
  wire \u2_Display/n4546 ;
  wire \u2_Display/n4547 ;
  wire \u2_Display/n4548 ;
  wire \u2_Display/n4549 ;
  wire \u2_Display/n455 ;
  wire \u2_Display/n4550 ;
  wire \u2_Display/n4551 ;
  wire \u2_Display/n4552 ;
  wire \u2_Display/n4553 ;
  wire \u2_Display/n4554 ;
  wire \u2_Display/n4555 ;
  wire \u2_Display/n4556 ;
  wire \u2_Display/n456 ;
  wire \u2_Display/n457 ;
  wire \u2_Display/n458 ;
  wire \u2_Display/n459 ;
  wire \u2_Display/n460 ;
  wire \u2_Display/n461 ;
  wire \u2_Display/n462 ;
  wire \u2_Display/n463 ;
  wire \u2_Display/n464 ;
  wire \u2_Display/n465 ;
  wire \u2_Display/n466 ;
  wire \u2_Display/n467 ;
  wire \u2_Display/n468 ;
  wire \u2_Display/n469 ;
  wire \u2_Display/n470 ;
  wire \u2_Display/n471 ;
  wire \u2_Display/n472 ;
  wire \u2_Display/n473 ;
  wire \u2_Display/n474 ;
  wire \u2_Display/n475 ;
  wire \u2_Display/n476 ;
  wire \u2_Display/n477 ;
  wire \u2_Display/n478 ;
  wire \u2_Display/n479 ;
  wire \u2_Display/n48 ;
  wire \u2_Display/n480 ;
  wire \u2_Display/n481 ;
  wire \u2_Display/n482 ;
  wire \u2_Display/n483 ;
  wire \u2_Display/n484 ;
  wire \u2_Display/n485 ;
  wire \u2_Display/n486 ;
  wire \u2_Display/n487 ;
  wire \u2_Display/n490 ;
  wire \u2_Display/n4909 ;
  wire \u2_Display/n491 ;
  wire \u2_Display/n492 ;
  wire \u2_Display/n493 ;
  wire \u2_Display/n494 ;
  wire \u2_Display/n4944 ;
  wire \u2_Display/n495 ;
  wire \u2_Display/n496 ;
  wire \u2_Display/n497 ;
  wire \u2_Display/n4979 ;
  wire \u2_Display/n498 ;
  wire \u2_Display/n499 ;
  wire \u2_Display/n50 ;
  wire \u2_Display/n500 ;
  wire \u2_Display/n501 ;
  wire \u2_Display/n5014 ;
  wire \u2_Display/n502 ;
  wire \u2_Display/n503 ;
  wire \u2_Display/n504 ;
  wire \u2_Display/n5049 ;
  wire \u2_Display/n505 ;
  wire \u2_Display/n506 ;
  wire \u2_Display/n507 ;
  wire \u2_Display/n508 ;
  wire \u2_Display/n5084 ;
  wire \u2_Display/n509 ;
  wire \u2_Display/n51 ;
  wire \u2_Display/n510 ;
  wire \u2_Display/n511 ;
  wire \u2_Display/n5119 ;
  wire \u2_Display/n512 ;
  wire \u2_Display/n513 ;
  wire \u2_Display/n514 ;
  wire \u2_Display/n515 ;
  wire \u2_Display/n5154 ;
  wire \u2_Display/n516 ;
  wire \u2_Display/n517 ;
  wire \u2_Display/n518 ;
  wire \u2_Display/n5189 ;
  wire \u2_Display/n519 ;
  wire \u2_Display/n5196 ;
  wire \u2_Display/n5197 ;
  wire \u2_Display/n5198 ;
  wire \u2_Display/n5199 ;
  wire \u2_Display/n520 ;
  wire \u2_Display/n5200 ;
  wire \u2_Display/n5201 ;
  wire \u2_Display/n5202 ;
  wire \u2_Display/n5203 ;
  wire \u2_Display/n5204 ;
  wire \u2_Display/n5205 ;
  wire \u2_Display/n5206 ;
  wire \u2_Display/n5207 ;
  wire \u2_Display/n5208 ;
  wire \u2_Display/n5209 ;
  wire \u2_Display/n521 ;
  wire \u2_Display/n5210 ;
  wire \u2_Display/n5211 ;
  wire \u2_Display/n5212 ;
  wire \u2_Display/n5213 ;
  wire \u2_Display/n5214 ;
  wire \u2_Display/n5215 ;
  wire \u2_Display/n5216 ;
  wire \u2_Display/n5217 ;
  wire \u2_Display/n5218 ;
  wire \u2_Display/n5219 ;
  wire \u2_Display/n522 ;
  wire \u2_Display/n5220 ;
  wire \u2_Display/n5221 ;
  wire \u2_Display/n5222 ;
  wire \u2_Display/n5223 ;
  wire \u2_Display/n5224 ;
  wire \u2_Display/n5227 ;
  wire \u2_Display/n5228 ;
  wire \u2_Display/n5229 ;
  wire \u2_Display/n5230 ;
  wire \u2_Display/n5231 ;
  wire \u2_Display/n5232 ;
  wire \u2_Display/n5233 ;
  wire \u2_Display/n5234 ;
  wire \u2_Display/n5235 ;
  wire \u2_Display/n5236 ;
  wire \u2_Display/n5237 ;
  wire \u2_Display/n5238 ;
  wire \u2_Display/n5239 ;
  wire \u2_Display/n5240 ;
  wire \u2_Display/n5241 ;
  wire \u2_Display/n5242 ;
  wire \u2_Display/n5243 ;
  wire \u2_Display/n5244 ;
  wire \u2_Display/n5245 ;
  wire \u2_Display/n5246 ;
  wire \u2_Display/n5247 ;
  wire \u2_Display/n5248 ;
  wire \u2_Display/n5249 ;
  wire \u2_Display/n525 ;
  wire \u2_Display/n5250 ;
  wire \u2_Display/n5251 ;
  wire \u2_Display/n5252 ;
  wire \u2_Display/n5253 ;
  wire \u2_Display/n5254 ;
  wire \u2_Display/n5255 ;
  wire \u2_Display/n5256 ;
  wire \u2_Display/n5257 ;
  wire \u2_Display/n5258 ;
  wire \u2_Display/n5259 ;
  wire \u2_Display/n526 ;
  wire \u2_Display/n5262 ;
  wire \u2_Display/n5263 ;
  wire \u2_Display/n5264 ;
  wire \u2_Display/n5265 ;
  wire \u2_Display/n5266 ;
  wire \u2_Display/n5267 ;
  wire \u2_Display/n5268 ;
  wire \u2_Display/n5269 ;
  wire \u2_Display/n527 ;
  wire \u2_Display/n5270 ;
  wire \u2_Display/n5271 ;
  wire \u2_Display/n5272 ;
  wire \u2_Display/n5273 ;
  wire \u2_Display/n5274 ;
  wire \u2_Display/n5275 ;
  wire \u2_Display/n5276 ;
  wire \u2_Display/n5277 ;
  wire \u2_Display/n5278 ;
  wire \u2_Display/n5279 ;
  wire \u2_Display/n528 ;
  wire \u2_Display/n5280 ;
  wire \u2_Display/n5281 ;
  wire \u2_Display/n5282 ;
  wire \u2_Display/n5283 ;
  wire \u2_Display/n5284 ;
  wire \u2_Display/n5285 ;
  wire \u2_Display/n5286 ;
  wire \u2_Display/n5287 ;
  wire \u2_Display/n5288 ;
  wire \u2_Display/n5289 ;
  wire \u2_Display/n529 ;
  wire \u2_Display/n5290 ;
  wire \u2_Display/n5291 ;
  wire \u2_Display/n5292 ;
  wire \u2_Display/n5293 ;
  wire \u2_Display/n5294 ;
  wire \u2_Display/n5297 ;
  wire \u2_Display/n5298 ;
  wire \u2_Display/n5299 ;
  wire \u2_Display/n530 ;
  wire \u2_Display/n5300 ;
  wire \u2_Display/n5301 ;
  wire \u2_Display/n5302 ;
  wire \u2_Display/n5303 ;
  wire \u2_Display/n5304 ;
  wire \u2_Display/n5305 ;
  wire \u2_Display/n5306 ;
  wire \u2_Display/n5307 ;
  wire \u2_Display/n5308 ;
  wire \u2_Display/n5309 ;
  wire \u2_Display/n531 ;
  wire \u2_Display/n5310 ;
  wire \u2_Display/n5311 ;
  wire \u2_Display/n5312 ;
  wire \u2_Display/n5313 ;
  wire \u2_Display/n5314 ;
  wire \u2_Display/n5315 ;
  wire \u2_Display/n5316 ;
  wire \u2_Display/n5317 ;
  wire \u2_Display/n5318 ;
  wire \u2_Display/n5319 ;
  wire \u2_Display/n532 ;
  wire \u2_Display/n5320 ;
  wire \u2_Display/n5321 ;
  wire \u2_Display/n5322 ;
  wire \u2_Display/n5323 ;
  wire \u2_Display/n5324 ;
  wire \u2_Display/n5325 ;
  wire \u2_Display/n5326 ;
  wire \u2_Display/n5327 ;
  wire \u2_Display/n5328 ;
  wire \u2_Display/n5329 ;
  wire \u2_Display/n533 ;
  wire \u2_Display/n5332 ;
  wire \u2_Display/n5333 ;
  wire \u2_Display/n5334 ;
  wire \u2_Display/n5335 ;
  wire \u2_Display/n5336 ;
  wire \u2_Display/n5337 ;
  wire \u2_Display/n5338 ;
  wire \u2_Display/n5339 ;
  wire \u2_Display/n534 ;
  wire \u2_Display/n5340 ;
  wire \u2_Display/n5341 ;
  wire \u2_Display/n5342 ;
  wire \u2_Display/n5343 ;
  wire \u2_Display/n5344 ;
  wire \u2_Display/n5345 ;
  wire \u2_Display/n5346 ;
  wire \u2_Display/n5347 ;
  wire \u2_Display/n5348 ;
  wire \u2_Display/n5349 ;
  wire \u2_Display/n535 ;
  wire \u2_Display/n5350 ;
  wire \u2_Display/n5351 ;
  wire \u2_Display/n5352 ;
  wire \u2_Display/n5353 ;
  wire \u2_Display/n5354 ;
  wire \u2_Display/n5355 ;
  wire \u2_Display/n5356 ;
  wire \u2_Display/n5357 ;
  wire \u2_Display/n5358 ;
  wire \u2_Display/n5359 ;
  wire \u2_Display/n536 ;
  wire \u2_Display/n5360 ;
  wire \u2_Display/n5361 ;
  wire \u2_Display/n5362 ;
  wire \u2_Display/n5363 ;
  wire \u2_Display/n5364 ;
  wire \u2_Display/n5367 ;
  wire \u2_Display/n5368 ;
  wire \u2_Display/n5369 ;
  wire \u2_Display/n537 ;
  wire \u2_Display/n5370 ;
  wire \u2_Display/n5371 ;
  wire \u2_Display/n5372 ;
  wire \u2_Display/n5373 ;
  wire \u2_Display/n5374 ;
  wire \u2_Display/n5375 ;
  wire \u2_Display/n5376 ;
  wire \u2_Display/n5377 ;
  wire \u2_Display/n5378 ;
  wire \u2_Display/n5379 ;
  wire \u2_Display/n538 ;
  wire \u2_Display/n5380 ;
  wire \u2_Display/n5381 ;
  wire \u2_Display/n5382 ;
  wire \u2_Display/n5383 ;
  wire \u2_Display/n5384 ;
  wire \u2_Display/n5385 ;
  wire \u2_Display/n5386 ;
  wire \u2_Display/n5387 ;
  wire \u2_Display/n5388 ;
  wire \u2_Display/n5389 ;
  wire \u2_Display/n539 ;
  wire \u2_Display/n5390 ;
  wire \u2_Display/n5391 ;
  wire \u2_Display/n5392 ;
  wire \u2_Display/n5393 ;
  wire \u2_Display/n5394 ;
  wire \u2_Display/n5395 ;
  wire \u2_Display/n5396 ;
  wire \u2_Display/n5397 ;
  wire \u2_Display/n5398 ;
  wire \u2_Display/n5399 ;
  wire \u2_Display/n540 ;
  wire \u2_Display/n5402 ;
  wire \u2_Display/n5403 ;
  wire \u2_Display/n5404 ;
  wire \u2_Display/n5405 ;
  wire \u2_Display/n5406 ;
  wire \u2_Display/n5407 ;
  wire \u2_Display/n5408 ;
  wire \u2_Display/n5409 ;
  wire \u2_Display/n541 ;
  wire \u2_Display/n5410 ;
  wire \u2_Display/n5411 ;
  wire \u2_Display/n5412 ;
  wire \u2_Display/n5413 ;
  wire \u2_Display/n5414 ;
  wire \u2_Display/n5415 ;
  wire \u2_Display/n5416 ;
  wire \u2_Display/n5417 ;
  wire \u2_Display/n5418 ;
  wire \u2_Display/n5419 ;
  wire \u2_Display/n542 ;
  wire \u2_Display/n5420 ;
  wire \u2_Display/n5421 ;
  wire \u2_Display/n5422 ;
  wire \u2_Display/n5423 ;
  wire \u2_Display/n5424 ;
  wire \u2_Display/n5425 ;
  wire \u2_Display/n5426 ;
  wire \u2_Display/n5427 ;
  wire \u2_Display/n5428 ;
  wire \u2_Display/n5429 ;
  wire \u2_Display/n543 ;
  wire \u2_Display/n5430 ;
  wire \u2_Display/n5431 ;
  wire \u2_Display/n5432 ;
  wire \u2_Display/n5433 ;
  wire \u2_Display/n5434 ;
  wire \u2_Display/n5437 ;
  wire \u2_Display/n5438 ;
  wire \u2_Display/n5439 ;
  wire \u2_Display/n544 ;
  wire \u2_Display/n5440 ;
  wire \u2_Display/n5441 ;
  wire \u2_Display/n5442 ;
  wire \u2_Display/n5443 ;
  wire \u2_Display/n5444 ;
  wire \u2_Display/n5445 ;
  wire \u2_Display/n5446 ;
  wire \u2_Display/n5447 ;
  wire \u2_Display/n5448 ;
  wire \u2_Display/n5449 ;
  wire \u2_Display/n545 ;
  wire \u2_Display/n5450 ;
  wire \u2_Display/n5451 ;
  wire \u2_Display/n5452 ;
  wire \u2_Display/n5453 ;
  wire \u2_Display/n5454 ;
  wire \u2_Display/n5455 ;
  wire \u2_Display/n5456 ;
  wire \u2_Display/n5457 ;
  wire \u2_Display/n5458 ;
  wire \u2_Display/n5459 ;
  wire \u2_Display/n546 ;
  wire \u2_Display/n5460 ;
  wire \u2_Display/n5461 ;
  wire \u2_Display/n5462 ;
  wire \u2_Display/n5463 ;
  wire \u2_Display/n5464 ;
  wire \u2_Display/n5465 ;
  wire \u2_Display/n5466 ;
  wire \u2_Display/n5467 ;
  wire \u2_Display/n5468 ;
  wire \u2_Display/n5469 ;
  wire \u2_Display/n547 ;
  wire \u2_Display/n5472 ;
  wire \u2_Display/n5473 ;
  wire \u2_Display/n5474 ;
  wire \u2_Display/n5475 ;
  wire \u2_Display/n5476 ;
  wire \u2_Display/n5477 ;
  wire \u2_Display/n5478 ;
  wire \u2_Display/n5479 ;
  wire \u2_Display/n548 ;
  wire \u2_Display/n5480 ;
  wire \u2_Display/n5481 ;
  wire \u2_Display/n5482 ;
  wire \u2_Display/n5483 ;
  wire \u2_Display/n5484 ;
  wire \u2_Display/n5485 ;
  wire \u2_Display/n5486 ;
  wire \u2_Display/n5487 ;
  wire \u2_Display/n5488 ;
  wire \u2_Display/n5489 ;
  wire \u2_Display/n549 ;
  wire \u2_Display/n5490 ;
  wire \u2_Display/n5491 ;
  wire \u2_Display/n5492 ;
  wire \u2_Display/n5493 ;
  wire \u2_Display/n5494 ;
  wire \u2_Display/n5495 ;
  wire \u2_Display/n5496 ;
  wire \u2_Display/n5497 ;
  wire \u2_Display/n5498 ;
  wire \u2_Display/n5499 ;
  wire \u2_Display/n550 ;
  wire \u2_Display/n5500 ;
  wire \u2_Display/n5501 ;
  wire \u2_Display/n5502 ;
  wire \u2_Display/n5503 ;
  wire \u2_Display/n5504 ;
  wire \u2_Display/n5507 ;
  wire \u2_Display/n5508 ;
  wire \u2_Display/n5509 ;
  wire \u2_Display/n551 ;
  wire \u2_Display/n5510 ;
  wire \u2_Display/n5511 ;
  wire \u2_Display/n5512 ;
  wire \u2_Display/n5513 ;
  wire \u2_Display/n5514 ;
  wire \u2_Display/n5515 ;
  wire \u2_Display/n5516 ;
  wire \u2_Display/n5517 ;
  wire \u2_Display/n5518 ;
  wire \u2_Display/n5519 ;
  wire \u2_Display/n552 ;
  wire \u2_Display/n5520 ;
  wire \u2_Display/n5521 ;
  wire \u2_Display/n5522 ;
  wire \u2_Display/n5523 ;
  wire \u2_Display/n5524 ;
  wire \u2_Display/n5525 ;
  wire \u2_Display/n5526 ;
  wire \u2_Display/n5527 ;
  wire \u2_Display/n5528 ;
  wire \u2_Display/n5529 ;
  wire \u2_Display/n553 ;
  wire \u2_Display/n5530 ;
  wire \u2_Display/n5531 ;
  wire \u2_Display/n5532 ;
  wire \u2_Display/n5533 ;
  wire \u2_Display/n5534 ;
  wire \u2_Display/n5535 ;
  wire \u2_Display/n5536 ;
  wire \u2_Display/n5537 ;
  wire \u2_Display/n5538 ;
  wire \u2_Display/n5539 ;
  wire \u2_Display/n554 ;
  wire \u2_Display/n5542 ;
  wire \u2_Display/n5543 ;
  wire \u2_Display/n5544 ;
  wire \u2_Display/n5545 ;
  wire \u2_Display/n5546 ;
  wire \u2_Display/n5547 ;
  wire \u2_Display/n5548 ;
  wire \u2_Display/n5549 ;
  wire \u2_Display/n555 ;
  wire \u2_Display/n5550 ;
  wire \u2_Display/n5551 ;
  wire \u2_Display/n5552 ;
  wire \u2_Display/n5553 ;
  wire \u2_Display/n5554 ;
  wire \u2_Display/n5555 ;
  wire \u2_Display/n5556 ;
  wire \u2_Display/n5557 ;
  wire \u2_Display/n5558 ;
  wire \u2_Display/n5559 ;
  wire \u2_Display/n556 ;
  wire \u2_Display/n5560 ;
  wire \u2_Display/n5561 ;
  wire \u2_Display/n5562 ;
  wire \u2_Display/n5563 ;
  wire \u2_Display/n5564 ;
  wire \u2_Display/n5565 ;
  wire \u2_Display/n5566 ;
  wire \u2_Display/n5567 ;
  wire \u2_Display/n5568 ;
  wire \u2_Display/n5569 ;
  wire \u2_Display/n557 ;
  wire \u2_Display/n5570 ;
  wire \u2_Display/n5571 ;
  wire \u2_Display/n5572 ;
  wire \u2_Display/n5573 ;
  wire \u2_Display/n5574 ;
  wire \u2_Display/n5577 ;
  wire \u2_Display/n5578 ;
  wire \u2_Display/n5579 ;
  wire \u2_Display/n5580 ;
  wire \u2_Display/n5581 ;
  wire \u2_Display/n5582 ;
  wire \u2_Display/n5583 ;
  wire \u2_Display/n5584 ;
  wire \u2_Display/n5585 ;
  wire \u2_Display/n5586 ;
  wire \u2_Display/n5587 ;
  wire \u2_Display/n5588 ;
  wire \u2_Display/n5589 ;
  wire \u2_Display/n5590 ;
  wire \u2_Display/n5591 ;
  wire \u2_Display/n5592 ;
  wire \u2_Display/n5593 ;
  wire \u2_Display/n5594 ;
  wire \u2_Display/n5595 ;
  wire \u2_Display/n5596 ;
  wire \u2_Display/n5597 ;
  wire \u2_Display/n5598 ;
  wire \u2_Display/n5599 ;
  wire \u2_Display/n560 ;
  wire \u2_Display/n5600 ;
  wire \u2_Display/n5601 ;
  wire \u2_Display/n5602 ;
  wire \u2_Display/n5603 ;
  wire \u2_Display/n5604 ;
  wire \u2_Display/n5605 ;
  wire \u2_Display/n5606 ;
  wire \u2_Display/n5607 ;
  wire \u2_Display/n5608 ;
  wire \u2_Display/n5609 ;
  wire \u2_Display/n561 ;
  wire \u2_Display/n5612 ;
  wire \u2_Display/n5613 ;
  wire \u2_Display/n5614 ;
  wire \u2_Display/n5615 ;
  wire \u2_Display/n5616 ;
  wire \u2_Display/n5617 ;
  wire \u2_Display/n5618 ;
  wire \u2_Display/n5619 ;
  wire \u2_Display/n562 ;
  wire \u2_Display/n5620 ;
  wire \u2_Display/n5621 ;
  wire \u2_Display/n5622 ;
  wire \u2_Display/n5623 ;
  wire \u2_Display/n5624 ;
  wire \u2_Display/n5625 ;
  wire \u2_Display/n5626 ;
  wire \u2_Display/n5627 ;
  wire \u2_Display/n5628 ;
  wire \u2_Display/n5629 ;
  wire \u2_Display/n563 ;
  wire \u2_Display/n5630 ;
  wire \u2_Display/n5631 ;
  wire \u2_Display/n5632 ;
  wire \u2_Display/n5633 ;
  wire \u2_Display/n5634 ;
  wire \u2_Display/n5635 ;
  wire \u2_Display/n5636 ;
  wire \u2_Display/n5637 ;
  wire \u2_Display/n5638 ;
  wire \u2_Display/n5639 ;
  wire \u2_Display/n564 ;
  wire \u2_Display/n5640 ;
  wire \u2_Display/n5641 ;
  wire \u2_Display/n5642 ;
  wire \u2_Display/n5643 ;
  wire \u2_Display/n5644 ;
  wire \u2_Display/n5647 ;
  wire \u2_Display/n5648 ;
  wire \u2_Display/n5649 ;
  wire \u2_Display/n565 ;
  wire \u2_Display/n5650 ;
  wire \u2_Display/n5651 ;
  wire \u2_Display/n5652 ;
  wire \u2_Display/n5653 ;
  wire \u2_Display/n5654 ;
  wire \u2_Display/n5655 ;
  wire \u2_Display/n5656 ;
  wire \u2_Display/n5657 ;
  wire \u2_Display/n5658 ;
  wire \u2_Display/n5659 ;
  wire \u2_Display/n566 ;
  wire \u2_Display/n5660 ;
  wire \u2_Display/n5661 ;
  wire \u2_Display/n5662 ;
  wire \u2_Display/n5663 ;
  wire \u2_Display/n5664 ;
  wire \u2_Display/n5665 ;
  wire \u2_Display/n5666 ;
  wire \u2_Display/n5667 ;
  wire \u2_Display/n5668 ;
  wire \u2_Display/n5669 ;
  wire \u2_Display/n567 ;
  wire \u2_Display/n5670 ;
  wire \u2_Display/n5671 ;
  wire \u2_Display/n5672 ;
  wire \u2_Display/n5673 ;
  wire \u2_Display/n5674 ;
  wire \u2_Display/n5675 ;
  wire \u2_Display/n5676 ;
  wire \u2_Display/n5677 ;
  wire \u2_Display/n5678 ;
  wire \u2_Display/n5679 ;
  wire \u2_Display/n568 ;
  wire \u2_Display/n569 ;
  wire \u2_Display/n570 ;
  wire \u2_Display/n571 ;
  wire \u2_Display/n572 ;
  wire \u2_Display/n573 ;
  wire \u2_Display/n574 ;
  wire \u2_Display/n575 ;
  wire \u2_Display/n576 ;
  wire \u2_Display/n577 ;
  wire \u2_Display/n578 ;
  wire \u2_Display/n579 ;
  wire \u2_Display/n580 ;
  wire \u2_Display/n581 ;
  wire \u2_Display/n582 ;
  wire \u2_Display/n583 ;
  wire \u2_Display/n584 ;
  wire \u2_Display/n585 ;
  wire \u2_Display/n586 ;
  wire \u2_Display/n587 ;
  wire \u2_Display/n588 ;
  wire \u2_Display/n589 ;
  wire \u2_Display/n590 ;
  wire \u2_Display/n591 ;
  wire \u2_Display/n592 ;
  wire \u2_Display/n595 ;
  wire \u2_Display/n596 ;
  wire \u2_Display/n597 ;
  wire \u2_Display/n598 ;
  wire \u2_Display/n599 ;
  wire \u2_Display/n600 ;
  wire \u2_Display/n601 ;
  wire \u2_Display/n602 ;
  wire \u2_Display/n603 ;
  wire \u2_Display/n604 ;
  wire \u2_Display/n605 ;
  wire \u2_Display/n606 ;
  wire \u2_Display/n607 ;
  wire \u2_Display/n6070 ;
  wire \u2_Display/n6071 ;
  wire \u2_Display/n6072 ;
  wire \u2_Display/n6073 ;
  wire \u2_Display/n6074 ;
  wire \u2_Display/n6075 ;
  wire \u2_Display/n6076 ;
  wire \u2_Display/n6077 ;
  wire \u2_Display/n6078 ;
  wire \u2_Display/n6079 ;
  wire \u2_Display/n608 ;
  wire \u2_Display/n6080 ;
  wire \u2_Display/n6081 ;
  wire \u2_Display/n6082 ;
  wire \u2_Display/n6083 ;
  wire \u2_Display/n6084 ;
  wire \u2_Display/n6085 ;
  wire \u2_Display/n6086 ;
  wire \u2_Display/n6087 ;
  wire \u2_Display/n6088 ;
  wire \u2_Display/n6089 ;
  wire \u2_Display/n609 ;
  wire \u2_Display/n6090 ;
  wire \u2_Display/n6091 ;
  wire \u2_Display/n6092 ;
  wire \u2_Display/n6093 ;
  wire \u2_Display/n6094 ;
  wire \u2_Display/n6095 ;
  wire \u2_Display/n6096 ;
  wire \u2_Display/n6097 ;
  wire \u2_Display/n6098 ;
  wire \u2_Display/n6099 ;
  wire \u2_Display/n610 ;
  wire \u2_Display/n6100 ;
  wire \u2_Display/n6101 ;
  wire \u2_Display/n6105 ;
  wire \u2_Display/n6106 ;
  wire \u2_Display/n6107 ;
  wire \u2_Display/n6108 ;
  wire \u2_Display/n6109 ;
  wire \u2_Display/n611 ;
  wire \u2_Display/n6110 ;
  wire \u2_Display/n6111 ;
  wire \u2_Display/n6112 ;
  wire \u2_Display/n6113 ;
  wire \u2_Display/n6114 ;
  wire \u2_Display/n6115 ;
  wire \u2_Display/n6116 ;
  wire \u2_Display/n6117 ;
  wire \u2_Display/n6118 ;
  wire \u2_Display/n6119 ;
  wire \u2_Display/n612 ;
  wire \u2_Display/n6120 ;
  wire \u2_Display/n6121 ;
  wire \u2_Display/n6122 ;
  wire \u2_Display/n6123 ;
  wire \u2_Display/n6124 ;
  wire \u2_Display/n6125 ;
  wire \u2_Display/n6126 ;
  wire \u2_Display/n6127 ;
  wire \u2_Display/n6128 ;
  wire \u2_Display/n6129 ;
  wire \u2_Display/n613 ;
  wire \u2_Display/n6130 ;
  wire \u2_Display/n6131 ;
  wire \u2_Display/n6132 ;
  wire \u2_Display/n6133 ;
  wire \u2_Display/n6134 ;
  wire \u2_Display/n6135 ;
  wire \u2_Display/n6136 ;
  wire \u2_Display/n614 ;
  wire \u2_Display/n6140 ;
  wire \u2_Display/n6141 ;
  wire \u2_Display/n6142 ;
  wire \u2_Display/n6143 ;
  wire \u2_Display/n6144 ;
  wire \u2_Display/n6145 ;
  wire \u2_Display/n6146 ;
  wire \u2_Display/n6147 ;
  wire \u2_Display/n6148 ;
  wire \u2_Display/n6149 ;
  wire \u2_Display/n615 ;
  wire \u2_Display/n6150 ;
  wire \u2_Display/n6151 ;
  wire \u2_Display/n6152 ;
  wire \u2_Display/n6153 ;
  wire \u2_Display/n6154 ;
  wire \u2_Display/n6155 ;
  wire \u2_Display/n6156 ;
  wire \u2_Display/n6157 ;
  wire \u2_Display/n6158 ;
  wire \u2_Display/n6159 ;
  wire \u2_Display/n616 ;
  wire \u2_Display/n6160 ;
  wire \u2_Display/n6161 ;
  wire \u2_Display/n6162 ;
  wire \u2_Display/n6163 ;
  wire \u2_Display/n6164 ;
  wire \u2_Display/n6165 ;
  wire \u2_Display/n6166 ;
  wire \u2_Display/n6167 ;
  wire \u2_Display/n6168 ;
  wire \u2_Display/n6169 ;
  wire \u2_Display/n617 ;
  wire \u2_Display/n6170 ;
  wire \u2_Display/n6171 ;
  wire \u2_Display/n6175 ;
  wire \u2_Display/n6176 ;
  wire \u2_Display/n6177 ;
  wire \u2_Display/n6178 ;
  wire \u2_Display/n6179 ;
  wire \u2_Display/n618 ;
  wire \u2_Display/n6180 ;
  wire \u2_Display/n6181 ;
  wire \u2_Display/n6182 ;
  wire \u2_Display/n6183 ;
  wire \u2_Display/n6184 ;
  wire \u2_Display/n6185 ;
  wire \u2_Display/n6186 ;
  wire \u2_Display/n6187 ;
  wire \u2_Display/n6188 ;
  wire \u2_Display/n6189 ;
  wire \u2_Display/n619 ;
  wire \u2_Display/n6190 ;
  wire \u2_Display/n6191 ;
  wire \u2_Display/n6192 ;
  wire \u2_Display/n6193 ;
  wire \u2_Display/n6194 ;
  wire \u2_Display/n6195 ;
  wire \u2_Display/n6196 ;
  wire \u2_Display/n6197 ;
  wire \u2_Display/n6198 ;
  wire \u2_Display/n6199 ;
  wire \u2_Display/n620 ;
  wire \u2_Display/n6200 ;
  wire \u2_Display/n6201 ;
  wire \u2_Display/n6202 ;
  wire \u2_Display/n6203 ;
  wire \u2_Display/n6204 ;
  wire \u2_Display/n6205 ;
  wire \u2_Display/n6206 ;
  wire \u2_Display/n621 ;
  wire \u2_Display/n6210 ;
  wire \u2_Display/n6211 ;
  wire \u2_Display/n6212 ;
  wire \u2_Display/n6213 ;
  wire \u2_Display/n6214 ;
  wire \u2_Display/n6215 ;
  wire \u2_Display/n6216 ;
  wire \u2_Display/n6217 ;
  wire \u2_Display/n6218 ;
  wire \u2_Display/n6219 ;
  wire \u2_Display/n622 ;
  wire \u2_Display/n6220 ;
  wire \u2_Display/n6221 ;
  wire \u2_Display/n6222 ;
  wire \u2_Display/n6223 ;
  wire \u2_Display/n6224 ;
  wire \u2_Display/n6225 ;
  wire \u2_Display/n6226 ;
  wire \u2_Display/n6227 ;
  wire \u2_Display/n6228 ;
  wire \u2_Display/n6229 ;
  wire \u2_Display/n623 ;
  wire \u2_Display/n6230 ;
  wire \u2_Display/n6231 ;
  wire \u2_Display/n6232 ;
  wire \u2_Display/n6233 ;
  wire \u2_Display/n6234 ;
  wire \u2_Display/n6235 ;
  wire \u2_Display/n6236 ;
  wire \u2_Display/n6237 ;
  wire \u2_Display/n6238 ;
  wire \u2_Display/n6239 ;
  wire \u2_Display/n624 ;
  wire \u2_Display/n6240 ;
  wire \u2_Display/n6241 ;
  wire \u2_Display/n6245 ;
  wire \u2_Display/n6246 ;
  wire \u2_Display/n6247 ;
  wire \u2_Display/n6248 ;
  wire \u2_Display/n6249 ;
  wire \u2_Display/n625 ;
  wire \u2_Display/n6250 ;
  wire \u2_Display/n6251 ;
  wire \u2_Display/n6252 ;
  wire \u2_Display/n6253 ;
  wire \u2_Display/n6254 ;
  wire \u2_Display/n6255 ;
  wire \u2_Display/n6256 ;
  wire \u2_Display/n6257 ;
  wire \u2_Display/n6258 ;
  wire \u2_Display/n6259 ;
  wire \u2_Display/n626 ;
  wire \u2_Display/n6260 ;
  wire \u2_Display/n6261 ;
  wire \u2_Display/n6262 ;
  wire \u2_Display/n6263 ;
  wire \u2_Display/n6264 ;
  wire \u2_Display/n6265 ;
  wire \u2_Display/n6266 ;
  wire \u2_Display/n6267 ;
  wire \u2_Display/n6268 ;
  wire \u2_Display/n6269 ;
  wire \u2_Display/n627 ;
  wire \u2_Display/n6270 ;
  wire \u2_Display/n6271 ;
  wire \u2_Display/n6272 ;
  wire \u2_Display/n6273 ;
  wire \u2_Display/n6274 ;
  wire \u2_Display/n6275 ;
  wire \u2_Display/n6276 ;
  wire \u2_Display/n6280 ;
  wire \u2_Display/n6281 ;
  wire \u2_Display/n6282 ;
  wire \u2_Display/n6283 ;
  wire \u2_Display/n6284 ;
  wire \u2_Display/n6285 ;
  wire \u2_Display/n6286 ;
  wire \u2_Display/n6287 ;
  wire \u2_Display/n6288 ;
  wire \u2_Display/n6289 ;
  wire \u2_Display/n6290 ;
  wire \u2_Display/n6291 ;
  wire \u2_Display/n6292 ;
  wire \u2_Display/n6293 ;
  wire \u2_Display/n6294 ;
  wire \u2_Display/n6295 ;
  wire \u2_Display/n6296 ;
  wire \u2_Display/n6297 ;
  wire \u2_Display/n6298 ;
  wire \u2_Display/n6299 ;
  wire \u2_Display/n630 ;
  wire \u2_Display/n6300 ;
  wire \u2_Display/n6301 ;
  wire \u2_Display/n6302 ;
  wire \u2_Display/n6303 ;
  wire \u2_Display/n6304 ;
  wire \u2_Display/n6305 ;
  wire \u2_Display/n6306 ;
  wire \u2_Display/n6307 ;
  wire \u2_Display/n6308 ;
  wire \u2_Display/n6309 ;
  wire \u2_Display/n631 ;
  wire \u2_Display/n6310 ;
  wire \u2_Display/n6311 ;
  wire \u2_Display/n6315 ;
  wire \u2_Display/n6316 ;
  wire \u2_Display/n6317 ;
  wire \u2_Display/n6318 ;
  wire \u2_Display/n6319 ;
  wire \u2_Display/n632 ;
  wire \u2_Display/n6320 ;
  wire \u2_Display/n6321 ;
  wire \u2_Display/n6322 ;
  wire \u2_Display/n6323 ;
  wire \u2_Display/n6324 ;
  wire \u2_Display/n6325 ;
  wire \u2_Display/n6326 ;
  wire \u2_Display/n6327 ;
  wire \u2_Display/n6328 ;
  wire \u2_Display/n6329 ;
  wire \u2_Display/n633 ;
  wire \u2_Display/n6330 ;
  wire \u2_Display/n6331 ;
  wire \u2_Display/n6332 ;
  wire \u2_Display/n6333 ;
  wire \u2_Display/n6334 ;
  wire \u2_Display/n6335 ;
  wire \u2_Display/n6336 ;
  wire \u2_Display/n6337 ;
  wire \u2_Display/n6338 ;
  wire \u2_Display/n6339 ;
  wire \u2_Display/n634 ;
  wire \u2_Display/n6340 ;
  wire \u2_Display/n6341 ;
  wire \u2_Display/n6342 ;
  wire \u2_Display/n6343 ;
  wire \u2_Display/n6344 ;
  wire \u2_Display/n6345 ;
  wire \u2_Display/n6346 ;
  wire \u2_Display/n635 ;
  wire \u2_Display/n6350 ;
  wire \u2_Display/n6351 ;
  wire \u2_Display/n6352 ;
  wire \u2_Display/n6353 ;
  wire \u2_Display/n636 ;
  wire \u2_Display/n637 ;
  wire \u2_Display/n638 ;
  wire \u2_Display/n639 ;
  wire \u2_Display/n640 ;
  wire \u2_Display/n641 ;
  wire \u2_Display/n642 ;
  wire \u2_Display/n643 ;
  wire \u2_Display/n644 ;
  wire \u2_Display/n645 ;
  wire \u2_Display/n646 ;
  wire \u2_Display/n647 ;
  wire \u2_Display/n648 ;
  wire \u2_Display/n649 ;
  wire \u2_Display/n650 ;
  wire \u2_Display/n651 ;
  wire \u2_Display/n652 ;
  wire \u2_Display/n653 ;
  wire \u2_Display/n654 ;
  wire \u2_Display/n655 ;
  wire \u2_Display/n656 ;
  wire \u2_Display/n657 ;
  wire \u2_Display/n658 ;
  wire \u2_Display/n659 ;
  wire \u2_Display/n660 ;
  wire \u2_Display/n661 ;
  wire \u2_Display/n662 ;
  wire \u2_Display/n665 ;
  wire \u2_Display/n666 ;
  wire \u2_Display/n667 ;
  wire \u2_Display/n668 ;
  wire \u2_Display/n669 ;
  wire \u2_Display/n670 ;
  wire \u2_Display/n671 ;
  wire \u2_Display/n672 ;
  wire \u2_Display/n673 ;
  wire \u2_Display/n674 ;
  wire \u2_Display/n675 ;
  wire \u2_Display/n676 ;
  wire \u2_Display/n677 ;
  wire \u2_Display/n678 ;
  wire \u2_Display/n679 ;
  wire \u2_Display/n680 ;
  wire \u2_Display/n681 ;
  wire \u2_Display/n682 ;
  wire \u2_Display/n683 ;
  wire \u2_Display/n684 ;
  wire \u2_Display/n685 ;
  wire \u2_Display/n686 ;
  wire \u2_Display/n687 ;
  wire \u2_Display/n688 ;
  wire \u2_Display/n689 ;
  wire \u2_Display/n690 ;
  wire \u2_Display/n691 ;
  wire \u2_Display/n692 ;
  wire \u2_Display/n693 ;
  wire \u2_Display/n694 ;
  wire \u2_Display/n695 ;
  wire \u2_Display/n696 ;
  wire \u2_Display/n697 ;
  wire \u2_Display/n700 ;
  wire \u2_Display/n701 ;
  wire \u2_Display/n702 ;
  wire \u2_Display/n703 ;
  wire \u2_Display/n704 ;
  wire \u2_Display/n705 ;
  wire \u2_Display/n706 ;
  wire \u2_Display/n707 ;
  wire \u2_Display/n708 ;
  wire \u2_Display/n709 ;
  wire \u2_Display/n710 ;
  wire \u2_Display/n711 ;
  wire \u2_Display/n712 ;
  wire \u2_Display/n713 ;
  wire \u2_Display/n714 ;
  wire \u2_Display/n715 ;
  wire \u2_Display/n716 ;
  wire \u2_Display/n717 ;
  wire \u2_Display/n718 ;
  wire \u2_Display/n719 ;
  wire \u2_Display/n720 ;
  wire \u2_Display/n721 ;
  wire \u2_Display/n722 ;
  wire \u2_Display/n723 ;
  wire \u2_Display/n724 ;
  wire \u2_Display/n725 ;
  wire \u2_Display/n726 ;
  wire \u2_Display/n727 ;
  wire \u2_Display/n728 ;
  wire \u2_Display/n729 ;
  wire \u2_Display/n730 ;
  wire \u2_Display/n731 ;
  wire \u2_Display/n732 ;
  wire \u2_Display/n735 ;
  wire \u2_Display/n736 ;
  wire \u2_Display/n737 ;
  wire \u2_Display/n738 ;
  wire \u2_Display/n739 ;
  wire \u2_Display/n740 ;
  wire \u2_Display/n741 ;
  wire \u2_Display/n742 ;
  wire \u2_Display/n743 ;
  wire \u2_Display/n744 ;
  wire \u2_Display/n745 ;
  wire \u2_Display/n746 ;
  wire \u2_Display/n747 ;
  wire \u2_Display/n748 ;
  wire \u2_Display/n749 ;
  wire \u2_Display/n750 ;
  wire \u2_Display/n751 ;
  wire \u2_Display/n752 ;
  wire \u2_Display/n753 ;
  wire \u2_Display/n754 ;
  wire \u2_Display/n755 ;
  wire \u2_Display/n756 ;
  wire \u2_Display/n757 ;
  wire \u2_Display/n758 ;
  wire \u2_Display/n759 ;
  wire \u2_Display/n760 ;
  wire \u2_Display/n761 ;
  wire \u2_Display/n762 ;
  wire \u2_Display/n763 ;
  wire \u2_Display/n764 ;
  wire \u2_Display/n765 ;
  wire \u2_Display/n766 ;
  wire \u2_Display/n767 ;
  wire \u2_Display/n770 ;
  wire \u2_Display/n771 ;
  wire \u2_Display/n772 ;
  wire \u2_Display/n773 ;
  wire \u2_Display/n774 ;
  wire \u2_Display/n775 ;
  wire \u2_Display/n776 ;
  wire \u2_Display/n777 ;
  wire \u2_Display/n778 ;
  wire \u2_Display/n779 ;
  wire \u2_Display/n780 ;
  wire \u2_Display/n781 ;
  wire \u2_Display/n782 ;
  wire \u2_Display/n783 ;
  wire \u2_Display/n784 ;
  wire \u2_Display/n785 ;
  wire \u2_Display/n786 ;
  wire \u2_Display/n787 ;
  wire \u2_Display/n788 ;
  wire \u2_Display/n789 ;
  wire \u2_Display/n790 ;
  wire \u2_Display/n791 ;
  wire \u2_Display/n792 ;
  wire \u2_Display/n793 ;
  wire \u2_Display/n794 ;
  wire \u2_Display/n795 ;
  wire \u2_Display/n796 ;
  wire \u2_Display/n797 ;
  wire \u2_Display/n798 ;
  wire \u2_Display/n799 ;
  wire \u2_Display/n800 ;
  wire \u2_Display/n801 ;
  wire \u2_Display/n802 ;
  wire \u2_Display/n805 ;
  wire \u2_Display/n806 ;
  wire \u2_Display/n807 ;
  wire \u2_Display/n808 ;
  wire \u2_Display/n809 ;
  wire \u2_Display/n810 ;
  wire \u2_Display/n811 ;
  wire \u2_Display/n812 ;
  wire \u2_Display/n813 ;
  wire \u2_Display/n814 ;
  wire \u2_Display/n815 ;
  wire \u2_Display/n816 ;
  wire \u2_Display/n817 ;
  wire \u2_Display/n818 ;
  wire \u2_Display/n819 ;
  wire \u2_Display/n820 ;
  wire \u2_Display/n821 ;
  wire \u2_Display/n822 ;
  wire \u2_Display/n823 ;
  wire \u2_Display/n824 ;
  wire \u2_Display/n825 ;
  wire \u2_Display/n826 ;
  wire \u2_Display/n827 ;
  wire \u2_Display/n828 ;
  wire \u2_Display/n829 ;
  wire \u2_Display/n830 ;
  wire \u2_Display/n831 ;
  wire \u2_Display/n832 ;
  wire \u2_Display/n833 ;
  wire \u2_Display/n834 ;
  wire \u2_Display/n835 ;
  wire \u2_Display/n836 ;
  wire \u2_Display/n837 ;
  wire \u2_Display/n840 ;
  wire \u2_Display/n841 ;
  wire \u2_Display/n842 ;
  wire \u2_Display/n843 ;
  wire \u2_Display/n844 ;
  wire \u2_Display/n845 ;
  wire \u2_Display/n846 ;
  wire \u2_Display/n847 ;
  wire \u2_Display/n848 ;
  wire \u2_Display/n849 ;
  wire \u2_Display/n850 ;
  wire \u2_Display/n851 ;
  wire \u2_Display/n852 ;
  wire \u2_Display/n853 ;
  wire \u2_Display/n854 ;
  wire \u2_Display/n855 ;
  wire \u2_Display/n856 ;
  wire \u2_Display/n857 ;
  wire \u2_Display/n858 ;
  wire \u2_Display/n859 ;
  wire \u2_Display/n860 ;
  wire \u2_Display/n861 ;
  wire \u2_Display/n862 ;
  wire \u2_Display/n863 ;
  wire \u2_Display/n864 ;
  wire \u2_Display/n865 ;
  wire \u2_Display/n866 ;
  wire \u2_Display/n867 ;
  wire \u2_Display/n868 ;
  wire \u2_Display/n869 ;
  wire \u2_Display/n870 ;
  wire \u2_Display/n871 ;
  wire \u2_Display/n872 ;
  wire \u2_Display/n875 ;
  wire \u2_Display/n876 ;
  wire \u2_Display/n877 ;
  wire \u2_Display/n878 ;
  wire \u2_Display/n879 ;
  wire \u2_Display/n880 ;
  wire \u2_Display/n881 ;
  wire \u2_Display/n882 ;
  wire \u2_Display/n883 ;
  wire \u2_Display/n884 ;
  wire \u2_Display/n885 ;
  wire \u2_Display/n886 ;
  wire \u2_Display/n887 ;
  wire \u2_Display/n888 ;
  wire \u2_Display/n889 ;
  wire \u2_Display/n890 ;
  wire \u2_Display/n891 ;
  wire \u2_Display/n892 ;
  wire \u2_Display/n893 ;
  wire \u2_Display/n894 ;
  wire \u2_Display/n895 ;
  wire \u2_Display/n896 ;
  wire \u2_Display/n897 ;
  wire \u2_Display/n898 ;
  wire \u2_Display/n899 ;
  wire \u2_Display/n900 ;
  wire \u2_Display/n901 ;
  wire \u2_Display/n902 ;
  wire \u2_Display/n903 ;
  wire \u2_Display/n904 ;
  wire \u2_Display/n905 ;
  wire \u2_Display/n906 ;
  wire \u2_Display/n907 ;
  wire \u2_Display/n910 ;
  wire \u2_Display/n911 ;
  wire \u2_Display/n912 ;
  wire \u2_Display/n913 ;
  wire \u2_Display/n914 ;
  wire \u2_Display/n915 ;
  wire \u2_Display/n916 ;
  wire \u2_Display/n917 ;
  wire \u2_Display/n918 ;
  wire \u2_Display/n919 ;
  wire \u2_Display/n920 ;
  wire \u2_Display/n921 ;
  wire \u2_Display/n922 ;
  wire \u2_Display/n923 ;
  wire \u2_Display/n924 ;
  wire \u2_Display/n925 ;
  wire \u2_Display/n926 ;
  wire \u2_Display/n927 ;
  wire \u2_Display/n928 ;
  wire \u2_Display/n929 ;
  wire \u2_Display/n930 ;
  wire \u2_Display/n931 ;
  wire \u2_Display/n932 ;
  wire \u2_Display/n933 ;
  wire \u2_Display/n934 ;
  wire \u2_Display/n935 ;
  wire \u2_Display/n936 ;
  wire \u2_Display/n937 ;
  wire \u2_Display/n938 ;
  wire \u2_Display/n939 ;
  wire \u2_Display/n940 ;
  wire \u2_Display/n941 ;
  wire \u2_Display/n942 ;
  wire \u2_Display/n945 ;
  wire \u2_Display/n946 ;
  wire \u2_Display/n947 ;
  wire \u2_Display/n948 ;
  wire \u2_Display/n949 ;
  wire \u2_Display/n95 ;
  wire \u2_Display/n950 ;
  wire \u2_Display/n951 ;
  wire \u2_Display/n952 ;
  wire \u2_Display/n953 ;
  wire \u2_Display/n954 ;
  wire \u2_Display/n955 ;
  wire \u2_Display/n956 ;
  wire \u2_Display/n957 ;
  wire \u2_Display/n958 ;
  wire \u2_Display/n959 ;
  wire \u2_Display/n960 ;
  wire \u2_Display/n961 ;
  wire \u2_Display/n962 ;
  wire \u2_Display/n963 ;
  wire \u2_Display/n964 ;
  wire \u2_Display/n965 ;
  wire \u2_Display/n966 ;
  wire \u2_Display/n967 ;
  wire \u2_Display/n968 ;
  wire \u2_Display/n969 ;
  wire \u2_Display/n97 ;
  wire \u2_Display/n970 ;
  wire \u2_Display/n971 ;
  wire \u2_Display/n972 ;
  wire \u2_Display/n973 ;
  wire \u2_Display/n974 ;
  wire \u2_Display/n975 ;
  wire \u2_Display/n976 ;
  wire \u2_Display/n977 ;
  wire \u2_Display/n980 ;
  wire \u2_Display/n981 ;
  wire \u2_Display/n982 ;
  wire \u2_Display/n983 ;
  wire \u2_Display/n984 ;
  wire \u2_Display/n985 ;
  wire \u2_Display/n986 ;
  wire \u2_Display/n987 ;
  wire \u2_Display/n988 ;
  wire \u2_Display/n989 ;
  wire \u2_Display/n990 ;
  wire \u2_Display/n991 ;
  wire \u2_Display/n992 ;
  wire \u2_Display/n993 ;
  wire \u2_Display/n994 ;
  wire \u2_Display/n995 ;
  wire \u2_Display/n996 ;
  wire \u2_Display/n997 ;
  wire \u2_Display/n998 ;
  wire \u2_Display/n999 ;
  wire \u2_Display/sub0_2/c11 ;
  wire \u2_Display/sub0_2/c3 ;
  wire \u2_Display/sub0_2/c7 ;
  wire \u2_Display/sub1_2/c3 ;
  wire \u2_Display/sub1_2/c7 ;
  wire \u2_Display/sub2_2/c3 ;
  wire \u2_Display/sub2_2/c7 ;
  wire \u2_Display/sub3_2/c11 ;
  wire \u2_Display/sub3_2/c3 ;
  wire \u2_Display/sub3_2/c7 ;
  wire vga_clk_pad;  // source/rtl/VGA_Demo.v(9)
  wire vga_de_pad;  // source/rtl/VGA_Demo.v(13)
  wire vga_hs_pad;  // source/rtl/VGA_Demo.v(10)
  wire vga_vs_pad;  // source/rtl/VGA_Demo.v(11)

  initial $sdf_annotate("VGA_Demo.sdf");
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1000|_al_u1002  (
    .b({\u2_Display/n3928 [0],\u2_Display/n3928 [2]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3925 ,\u2_Display/n3923 }),
    .f({\u2_Display/n3960 ,\u2_Display/n3958 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1001|_al_u1004  (
    .b({\u2_Display/n3928 [1],\u2_Display/n3928 [4]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3924 ,\u2_Display/n3921 }),
    .f({\u2_Display/n3959 ,\u2_Display/n3956 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1003|_al_u1006  (
    .b({\u2_Display/n3928 [3],\u2_Display/n3928 [6]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3922 ,\u2_Display/n3919 }),
    .f({\u2_Display/n3957 ,\u2_Display/n3954 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1005|_al_u1008  (
    .b({\u2_Display/n3928 [5],\u2_Display/n3928 [8]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3920 ,\u2_Display/n3917 }),
    .f({\u2_Display/n3955 ,\u2_Display/n3952 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1007|_al_u1010  (
    .b({\u2_Display/n3928 [7],\u2_Display/n3928 [10]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3918 ,\u2_Display/n3915 }),
    .f({\u2_Display/n3953 ,\u2_Display/n3950 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1009|_al_u1013  (
    .b({\u2_Display/n3928 [9],\u2_Display/n3928 [13]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3916 ,\u2_Display/n3912 }),
    .f({\u2_Display/n3951 ,\u2_Display/n3947 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1011|_al_u1016  (
    .b({\u2_Display/n3928 [11],\u2_Display/n3928 [16]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3914 ,\u2_Display/n3909 }),
    .f({\u2_Display/n3949 ,\u2_Display/n3944 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1012|_al_u1014  (
    .b({\u2_Display/n3928 [12],\u2_Display/n3928 [14]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3913 ,\u2_Display/n3911 }),
    .f({\u2_Display/n3948 ,\u2_Display/n3946 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1015|_al_u1018  (
    .b({\u2_Display/n3928 [15],\u2_Display/n3928 [18]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3910 ,\u2_Display/n3907 }),
    .f({\u2_Display/n3945 ,\u2_Display/n3942 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1017|_al_u1020  (
    .b({\u2_Display/n3928 [17],\u2_Display/n3928 [20]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3908 ,\u2_Display/n3905 }),
    .f({\u2_Display/n3943 ,\u2_Display/n3940 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1019|_al_u1022  (
    .b({\u2_Display/n3928 [19],\u2_Display/n3928 [22]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3906 ,\u2_Display/n3903 }),
    .f({\u2_Display/n3941 ,\u2_Display/n3938 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1021|_al_u1024  (
    .b({\u2_Display/n3928 [21],\u2_Display/n3928 [24]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3904 ,\u2_Display/n3901 }),
    .f({\u2_Display/n3939 ,\u2_Display/n3936 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1023|_al_u1026  (
    .b({\u2_Display/n3928 [23],\u2_Display/n3928 [26]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3902 ,\u2_Display/n3899 }),
    .f({\u2_Display/n3937 ,\u2_Display/n3934 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1025|_al_u1029  (
    .b({\u2_Display/n3928 [25],\u2_Display/n3928 [29]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3900 ,\u2_Display/n3896 }),
    .f({\u2_Display/n3935 ,\u2_Display/n3931 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1027|_al_u1031  (
    .b({\u2_Display/n3928 [27],\u2_Display/n3928 [31]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3898 ,\u2_Display/n3894 }),
    .f({\u2_Display/n3933 ,\u2_Display/n3929 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1028|_al_u1030  (
    .b({\u2_Display/n3928 [28],\u2_Display/n3928 [30]}),
    .c({\u2_Display/n3926 ,\u2_Display/n3926 }),
    .d({\u2_Display/n3897 ,\u2_Display/n3895 }),
    .f({\u2_Display/n3932 ,\u2_Display/n3930 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1032|_al_u1034  (
    .b({\u2_Display/n5051 [0],\u2_Display/n5051 [2]}),
    .c({\u2_Display/n5049 ,\u2_Display/n5049 }),
    .d({\u2_Display/n6206 ,\u2_Display/n6204 }),
    .f({\u2_Display/n6241 ,\u2_Display/n6239 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .MODE("LOGIC"))
    _al_u1033 (
    .b({open_n408,\u2_Display/n5051 [1]}),
    .c({open_n409,\u2_Display/n5049 }),
    .d({open_n412,\u2_Display/n6205 }),
    .f({open_n426,\u2_Display/n6240 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1035|_al_u1036  (
    .b({\u2_Display/n5051 [3],\u2_Display/n5051 [4]}),
    .c({\u2_Display/n5049 ,\u2_Display/n5049 }),
    .d({\u2_Display/n6203 ,\u2_Display/n6202 }),
    .f({\u2_Display/n6238 ,\u2_Display/n6237 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1037|_al_u1038  (
    .b({\u2_Display/n5051 [5],\u2_Display/n5051 [6]}),
    .c({\u2_Display/n5049 ,\u2_Display/n5049 }),
    .d({\u2_Display/n6201 ,\u2_Display/n6200 }),
    .f({\u2_Display/n6236 ,\u2_Display/n6235 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1039|_al_u1040  (
    .b({\u2_Display/n5051 [7],\u2_Display/n5051 [8]}),
    .c({\u2_Display/n5049 ,\u2_Display/n5049 }),
    .d({\u2_Display/n6199 ,\u2_Display/n6198 }),
    .f({\u2_Display/n6234 ,\u2_Display/n6233 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u1041|_al_u1042  (
    .b({\u2_Display/n5049 ,\u2_Display/n5051 [10]}),
    .c({\u2_Display/n5051 [9],\u2_Display/n5049 }),
    .d({\u2_Display/n6197 ,\u2_Display/n6196 }),
    .f({\u2_Display/n6232 ,\u2_Display/n6231 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1043|_al_u1635  (
    .b({\u2_Display/n5051 [11],\u2_Display/n1787 [24]}),
    .c({\u2_Display/n5049 ,\u2_Display/n1785 }),
    .d({\u2_Display/n6195 ,\u2_Display/n1760 }),
    .f({\u2_Display/n6230 ,\u2_Display/n1795 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1044|_al_u1049  (
    .b({\u2_Display/n5051 [12],\u2_Display/n5051 [17]}),
    .c({\u2_Display/n5049 ,\u2_Display/n5049 }),
    .d({\u2_Display/n6194 ,\u2_Display/n6189 }),
    .f({\u2_Display/n6229 ,\u2_Display/n6224 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1045|_al_u1046  (
    .b({\u2_Display/n5051 [13],\u2_Display/n5051 [14]}),
    .c({\u2_Display/n5049 ,\u2_Display/n5049 }),
    .d({\u2_Display/n6193 ,\u2_Display/n6192 }),
    .f({\u2_Display/n6228 ,\u2_Display/n6227 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100101011001010),
    .MODE("LOGIC"))
    \_al_u1047|_al_u1053  (
    .a({\u2_Display/n5051 [15],open_n602}),
    .b({\u2_Display/n6191 ,\u2_Display/n5051 [21]}),
    .c({\u2_Display/n5049 ,\u2_Display/n5049 }),
    .d({open_n605,\u2_Display/n6185 }),
    .f({\u2_Display/n6226 ,\u2_Display/n6220 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1048|_al_u1050  (
    .b({\u2_Display/n5051 [16],\u2_Display/n5051 [18]}),
    .c({\u2_Display/n5049 ,\u2_Display/n5049 }),
    .d({\u2_Display/n6190 ,\u2_Display/n6188 }),
    .f({\u2_Display/n6225 ,\u2_Display/n6223 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1051|_al_u1057  (
    .b({\u2_Display/n5051 [19],\u2_Display/n5051 [25]}),
    .c({\u2_Display/n5049 ,\u2_Display/n5049 }),
    .d({\u2_Display/n6187 ,\u2_Display/n6181 }),
    .f({\u2_Display/n6222 ,\u2_Display/n6216 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1052|_al_u1054  (
    .b({\u2_Display/n5051 [20],\u2_Display/n5051 [22]}),
    .c({\u2_Display/n5049 ,\u2_Display/n5049 }),
    .d({\u2_Display/n6186 ,\u2_Display/n6184 }),
    .f({\u2_Display/n6221 ,\u2_Display/n6219 }));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1110111000100010),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1055|_al_u1061  (
    .a({open_n698,\u2_Display/n5051 [29]}),
    .b({\u2_Display/n5051 [23],\u2_Display/n5049 }),
    .c({\u2_Display/n5049 ,open_n699}),
    .d({\u2_Display/n6183 ,\u2_Display/n6177 }),
    .f({\u2_Display/n6218 ,\u2_Display/n6212 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1056|_al_u1058  (
    .b({\u2_Display/n5051 [24],\u2_Display/n5051 [26]}),
    .c({\u2_Display/n5049 ,\u2_Display/n5049 }),
    .d({\u2_Display/n6182 ,\u2_Display/n6180 }),
    .f({\u2_Display/n6217 ,\u2_Display/n6215 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1059|_al_u1063  (
    .b({\u2_Display/n5051 [27],\u2_Display/n5051 [31]}),
    .c({\u2_Display/n5049 ,\u2_Display/n5049 }),
    .d({\u2_Display/n6179 ,\u2_Display/n6175 }),
    .f({\u2_Display/n6214 ,\u2_Display/n6210 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1060|_al_u1062  (
    .b({\u2_Display/n5051 [28],\u2_Display/n5051 [30]}),
    .c({\u2_Display/n5049 ,\u2_Display/n5049 }),
    .d({\u2_Display/n6178 ,\u2_Display/n6176 }),
    .f({\u2_Display/n6213 ,\u2_Display/n6211 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1064|_al_u1068  (
    .b({\u2_Display/n559 [0],\u2_Display/n559 [4]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n556 ,\u2_Display/n552 }),
    .f({\u2_Display/n591 ,\u2_Display/n587 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u1065|_al_u1066  (
    .b({\u2_Display/n555 ,\u2_Display/n559 [2]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n559 [1],\u2_Display/n554 }),
    .f({\u2_Display/n590 ,\u2_Display/n589 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1067|_al_u1070  (
    .b({\u2_Display/n559 [3],\u2_Display/n559 [6]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n553 ,\u2_Display/n550 }),
    .f({\u2_Display/n588 ,\u2_Display/n585 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1069|_al_u1072  (
    .b({\u2_Display/n559 [5],\u2_Display/n559 [8]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n551 ,\u2_Display/n548 }),
    .f({\u2_Display/n586 ,\u2_Display/n583 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1071|_al_u1074  (
    .b({\u2_Display/n559 [7],\u2_Display/n559 [10]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n549 ,\u2_Display/n546 }),
    .f({\u2_Display/n584 ,\u2_Display/n581 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1073|_al_u1076  (
    .b({\u2_Display/n559 [9],\u2_Display/n559 [12]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n547 ,\u2_Display/n544 }),
    .f({\u2_Display/n582 ,\u2_Display/n579 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1075|_al_u1078  (
    .b({\u2_Display/n559 [11],\u2_Display/n559 [14]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n545 ,\u2_Display/n542 }),
    .f({\u2_Display/n580 ,\u2_Display/n577 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1077|_al_u1080  (
    .b({\u2_Display/n559 [13],\u2_Display/n559 [16]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n543 ,\u2_Display/n540 }),
    .f({\u2_Display/n578 ,\u2_Display/n575 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1079|_al_u1082  (
    .b({\u2_Display/n559 [15],\u2_Display/n559 [18]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n541 ,\u2_Display/n538 }),
    .f({\u2_Display/n576 ,\u2_Display/n573 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1081|_al_u1084  (
    .b({\u2_Display/n559 [17],\u2_Display/n559 [20]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n539 ,\u2_Display/n536 }),
    .f({\u2_Display/n574 ,\u2_Display/n571 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1083|_al_u1086  (
    .b({\u2_Display/n559 [19],\u2_Display/n559 [22]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n537 ,\u2_Display/n534 }),
    .f({\u2_Display/n572 ,\u2_Display/n569 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1085|_al_u1088  (
    .b({\u2_Display/n559 [21],\u2_Display/n559 [24]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n535 ,\u2_Display/n532 }),
    .f({\u2_Display/n570 ,\u2_Display/n567 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1087|_al_u1090  (
    .b({\u2_Display/n559 [23],\u2_Display/n559 [26]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n533 ,\u2_Display/n530 }),
    .f({\u2_Display/n568 ,\u2_Display/n565 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1089|_al_u1092  (
    .b({\u2_Display/n559 [25],\u2_Display/n559 [28]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n531 ,\u2_Display/n528 }),
    .f({\u2_Display/n566 ,\u2_Display/n563 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1091|_al_u1094  (
    .b({\u2_Display/n559 [27],\u2_Display/n559 [30]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n529 ,\u2_Display/n526 }),
    .f({\u2_Display/n564 ,\u2_Display/n561 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1093|_al_u1095  (
    .b({\u2_Display/n559 [29],\u2_Display/n559 [31]}),
    .c({\u2_Display/n557 ,\u2_Display/n557 }),
    .d({\u2_Display/n527 ,\u2_Display/n525 }),
    .f({\u2_Display/n562 ,\u2_Display/n560 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1096|_al_u1098  (
    .b({\u2_Display/n1682 [0],\u2_Display/n1682 [2]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1679 ,\u2_Display/n1677 }),
    .f({\u2_Display/n1714 ,\u2_Display/n1712 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1097|_al_u1100  (
    .b({\u2_Display/n1682 [1],\u2_Display/n1682 [4]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1678 ,\u2_Display/n1675 }),
    .f({\u2_Display/n1713 ,\u2_Display/n1710 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1099|_al_u1102  (
    .b({\u2_Display/n1682 [3],\u2_Display/n1682 [6]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1676 ,\u2_Display/n1673 }),
    .f({\u2_Display/n1711 ,\u2_Display/n1708 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1101|_al_u1104  (
    .b({\u2_Display/n1682 [5],\u2_Display/n1682 [8]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1674 ,\u2_Display/n1671 }),
    .f({\u2_Display/n1709 ,\u2_Display/n1706 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1103|_al_u1106  (
    .b({\u2_Display/n1682 [7],\u2_Display/n1682 [10]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1672 ,\u2_Display/n1669 }),
    .f({\u2_Display/n1707 ,\u2_Display/n1704 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u1105|_al_u1108  (
    .b({\u2_Display/n1680 ,\u2_Display/n1682 [12]}),
    .c({\u2_Display/n1682 [9],\u2_Display/n1680 }),
    .d({\u2_Display/n1670 ,\u2_Display/n1667 }),
    .f({\u2_Display/n1705 ,\u2_Display/n1702 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1107|_al_u1110  (
    .b({\u2_Display/n1682 [11],\u2_Display/n1682 [14]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1668 ,\u2_Display/n1665 }),
    .f({\u2_Display/n1703 ,\u2_Display/n1700 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1109|_al_u1112  (
    .b({\u2_Display/n1682 [13],\u2_Display/n1682 [16]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1666 ,\u2_Display/n1663 }),
    .f({\u2_Display/n1701 ,\u2_Display/n1698 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1111|_al_u1114  (
    .b({\u2_Display/n1682 [15],\u2_Display/n1682 [18]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1664 ,\u2_Display/n1661 }),
    .f({\u2_Display/n1699 ,\u2_Display/n1696 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u1113|_al_u1117  (
    .b({\u2_Display/n1662 ,\u2_Display/n1682 [21]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1682 [17],\u2_Display/n1658 }),
    .f({\u2_Display/n1697 ,\u2_Display/n1693 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1115|_al_u1120  (
    .b({\u2_Display/n1682 [19],\u2_Display/n1682 [24]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1660 ,\u2_Display/n1655 }),
    .f({\u2_Display/n1695 ,\u2_Display/n1690 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1116|_al_u1118  (
    .b({\u2_Display/n1682 [20],\u2_Display/n1682 [22]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1659 ,\u2_Display/n1657 }),
    .f({\u2_Display/n1694 ,\u2_Display/n1692 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1119|_al_u1122  (
    .b({\u2_Display/n1682 [23],\u2_Display/n1682 [26]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1656 ,\u2_Display/n1653 }),
    .f({\u2_Display/n1691 ,\u2_Display/n1688 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1121|_al_u1125  (
    .b({\u2_Display/n1682 [25],\u2_Display/n1682 [29]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1654 ,\u2_Display/n1650 }),
    .f({\u2_Display/n1689 ,\u2_Display/n1685 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1123|_al_u1127  (
    .b({\u2_Display/n1682 [27],\u2_Display/n1682 [31]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1652 ,\u2_Display/n1648 }),
    .f({\u2_Display/n1687 ,\u2_Display/n1683 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1124|_al_u1126  (
    .b({\u2_Display/n1682 [28],\u2_Display/n1682 [30]}),
    .c({\u2_Display/n1680 ,\u2_Display/n1680 }),
    .d({\u2_Display/n1651 ,\u2_Display/n1649 }),
    .f({\u2_Display/n1686 ,\u2_Display/n1684 }));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1100101011001010),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1128|_al_u1344  (
    .a({open_n1562,\u2_Display/n2840 [31]}),
    .b({\u2_Display/n2805 [0],\u2_Display/n2806 }),
    .c({\u2_Display/n2803 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2802 ,open_n1565}),
    .f({\u2_Display/n2837 ,\u2_Display/n2841 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1129|_al_u1132  (
    .b({\u2_Display/n2805 [1],\u2_Display/n2805 [4]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2801 ,\u2_Display/n2798 }),
    .f({\u2_Display/n2836 ,\u2_Display/n2833 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .MODE("LOGIC"))
    _al_u1130 (
    .b({open_n1608,\u2_Display/n2805 [2]}),
    .c({open_n1609,\u2_Display/n2803 }),
    .d({open_n1612,\u2_Display/n2800 }),
    .f({open_n1626,\u2_Display/n2835 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1131|_al_u1134  (
    .b({\u2_Display/n2805 [3],\u2_Display/n2805 [6]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2799 ,\u2_Display/n2796 }),
    .f({\u2_Display/n2834 ,\u2_Display/n2831 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1133|_al_u1136  (
    .b({\u2_Display/n2805 [5],\u2_Display/n2805 [8]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2797 ,\u2_Display/n2794 }),
    .f({\u2_Display/n2832 ,\u2_Display/n2829 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1135|_al_u1138  (
    .b({\u2_Display/n2805 [7],\u2_Display/n2805 [10]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2795 ,\u2_Display/n2792 }),
    .f({\u2_Display/n2830 ,\u2_Display/n2827 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1137|_al_u1140  (
    .b({\u2_Display/n2805 [9],\u2_Display/n2805 [12]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2793 ,\u2_Display/n2790 }),
    .f({\u2_Display/n2828 ,\u2_Display/n2825 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1139|_al_u1142  (
    .b({\u2_Display/n2805 [11],\u2_Display/n2805 [14]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2791 ,\u2_Display/n2788 }),
    .f({\u2_Display/n2826 ,\u2_Display/n2823 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1141|_al_u1145  (
    .b({\u2_Display/n2805 [13],\u2_Display/n2805 [17]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2789 ,\u2_Display/n2785 }),
    .f({\u2_Display/n2824 ,\u2_Display/n2820 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1143|_al_u1148  (
    .b({\u2_Display/n2805 [15],\u2_Display/n2805 [20]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2787 ,\u2_Display/n2782 }),
    .f({\u2_Display/n2822 ,\u2_Display/n2817 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1144|_al_u1146  (
    .b({\u2_Display/n2805 [16],\u2_Display/n2805 [18]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2786 ,\u2_Display/n2784 }),
    .f({\u2_Display/n2821 ,\u2_Display/n2819 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1147|_al_u1150  (
    .b({\u2_Display/n2805 [19],\u2_Display/n2805 [22]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2783 ,\u2_Display/n2780 }),
    .f({\u2_Display/n2818 ,\u2_Display/n2815 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1149|_al_u1153  (
    .b({\u2_Display/n2805 [21],\u2_Display/n2805 [25]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2781 ,\u2_Display/n2777 }),
    .f({\u2_Display/n2816 ,\u2_Display/n2812 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1151|_al_u1157  (
    .b({\u2_Display/n2805 [23],\u2_Display/n2805 [29]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2779 ,\u2_Display/n2773 }),
    .f({\u2_Display/n2814 ,\u2_Display/n2808 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1152|_al_u1154  (
    .b({\u2_Display/n2805 [24],\u2_Display/n2805 [26]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2778 ,\u2_Display/n2776 }),
    .f({\u2_Display/n2813 ,\u2_Display/n2811 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1155|_al_u1159  (
    .b({\u2_Display/n2805 [27],\u2_Display/n2805 [31]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2775 ,\u2_Display/n2771 }),
    .f({\u2_Display/n2810 ,\u2_Display/n2806 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1156|_al_u1158  (
    .b({\u2_Display/n2805 [28],\u2_Display/n2805 [30]}),
    .c({\u2_Display/n2803 ,\u2_Display/n2803 }),
    .d({\u2_Display/n2774 ,\u2_Display/n2772 }),
    .f({\u2_Display/n2809 ,\u2_Display/n2807 }));
  EG_PHY_LSLICE #(
    //.LUTF0("((A*~(~C*D))*~(B)*~(0)+(A*~(~C*D))*B*~(0)+~((A*~(~C*D)))*B*0+(A*~(~C*D))*B*0)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("((A*~(~C*D))*~(B)*~(1)+(A*~(~C*D))*B*~(1)+~((A*~(~C*D)))*B*1+(A*~(~C*D))*B*1)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1010000010101010),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1160|_al_u1166  (
    .a({open_n1972,\u2_Display/n145 }),
    .b({open_n1973,\u2_Display/n104 }),
    .c({on_off_pad[2],on_off_pad[4]}),
    .d({on_off_pad[3],\u2_Display/mux11_b0_sel_is_0_o }),
    .e({open_n1976,on_off_pad[1]}),
    .f({\u2_Display/mux11_b0_sel_is_0_o ,\u2_Display/n236 [0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    .INIT_LUT0(16'b0000000000001111),
    .MODE("LOGIC"))
    _al_u1161 (
    .c({open_n2001,on_off_pad[3]}),
    .d({open_n2004,on_off_pad[4]}),
    .f({open_n2018,\u2_Display/mux5_b0_sel_is_0_o }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTG0("(D*C*B*A)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u1162 (
    .a({open_n2024,\u2_Display/n141 }),
    .b({open_n2025,\u2_Display/n144 }),
    .c({open_n2026,\u2_Display/n136 }),
    .d({open_n2029,\u2_Display/n138 }),
    .f({open_n2047,\u2_Display/n145 }));
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~(A*B)*~(C*D))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("~(~(A*B)*~(C*D))"),
    //.LUTG1("(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111100010001000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111100010001000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1163|u2_Display/reg3_b10  (
    .a({open_n2053,\u2_Display/i [10]}),
    .b({open_n2054,_al_u1168_o}),
    .c({on_off_pad[0],on_off_pad[0]}),
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({on_off_pad[1],\u2_Display/n5668 }),
    .f({\u2_Display/mux19_b0_sel_is_0_o ,open_n2072}),
    .q({open_n2076,\u2_Display/i [10]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1164|u2_Display/reg1_b0  (
    .a({\u2_Display/n44 ,open_n2077}),
    .b({\u2_Display/n45 ,\u2_Display/n236 [0]}),
    .c({\u2_Display/n48 ,on_off_pad[0]}),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({\u2_Display/n50 ,\u2_Display/n51 }),
    .sr(rst_n_pad),
    .f({\u2_Display/n51 ,open_n2095}),
    .q({open_n2099,lcd_data[23]}));  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTG0("(D*C*B*A)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u1165 (
    .a({open_n2100,\u2_Display/n95 }),
    .b({open_n2101,\u2_Display/n97 }),
    .c({open_n2102,\u2_Display/n100 }),
    .d({open_n2105,\u2_Display/n103 }),
    .f({open_n2123,\u2_Display/n104 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTG0("(~C*B*D)"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTG0(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u1168 (
    .b({open_n2131,\u2_Display/mux19_b0_sel_is_0_o }),
    .c({open_n2132,on_off_pad[4]}),
    .d({open_n2135,\u2_Display/mux11_b0_sel_is_0_o }),
    .f({open_n2153,_al_u1168_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(1*D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1170|_al_u1172  (
    .a({\u1_Driver/vcnt [6],_al_u1171_o}),
    .b({\u1_Driver/vcnt [7],\u1_Driver/vcnt [1]}),
    .c({\u1_Driver/vcnt [8],\u1_Driver/vcnt [11]}),
    .d({\u1_Driver/vcnt [9],\u1_Driver/vcnt [3]}),
    .e({open_n2161,\u1_Driver/vcnt [5]}),
    .f({_al_u1170_o,\u1_Driver/n6_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1185|_al_u1189  (
    .b({\u2_Display/n3963 [0],\u2_Display/n3963 [4]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3960 ,\u2_Display/n3956 }),
    .f({\u2_Display/n3995 ,\u2_Display/n3991 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1186|_al_u1187  (
    .b({\u2_Display/n3963 [1],\u2_Display/n3963 [2]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3959 ,\u2_Display/n3958 }),
    .f({\u2_Display/n3994 ,\u2_Display/n3993 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1188|_al_u1191  (
    .b({\u2_Display/n3963 [3],\u2_Display/n3963 [6]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3957 ,\u2_Display/n3954 }),
    .f({\u2_Display/n3992 ,\u2_Display/n3989 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1190|_al_u1193  (
    .b({\u2_Display/n3963 [5],\u2_Display/n3963 [8]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3955 ,\u2_Display/n3952 }),
    .f({\u2_Display/n3990 ,\u2_Display/n3987 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1192|_al_u1195  (
    .b({\u2_Display/n3963 [7],\u2_Display/n3963 [10]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3953 ,\u2_Display/n3950 }),
    .f({\u2_Display/n3988 ,\u2_Display/n3985 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1194|_al_u1198  (
    .b({\u2_Display/n3963 [9],\u2_Display/n3963 [13]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3951 ,\u2_Display/n3947 }),
    .f({\u2_Display/n3986 ,\u2_Display/n3982 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1196|_al_u1201  (
    .b({\u2_Display/n3963 [11],\u2_Display/n3963 [16]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3949 ,\u2_Display/n3944 }),
    .f({\u2_Display/n3984 ,\u2_Display/n3979 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1197|_al_u1199  (
    .b({\u2_Display/n3963 [12],\u2_Display/n3963 [14]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3948 ,\u2_Display/n3946 }),
    .f({\u2_Display/n3983 ,\u2_Display/n3981 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1200|_al_u1203  (
    .b({\u2_Display/n3963 [15],\u2_Display/n3963 [18]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3945 ,\u2_Display/n3942 }),
    .f({\u2_Display/n3980 ,\u2_Display/n3977 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u1202|_al_u1205  (
    .b({\u2_Display/n3943 ,\u2_Display/n3963 [20]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3963 [17],\u2_Display/n3940 }),
    .f({\u2_Display/n3978 ,\u2_Display/n3975 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1204|_al_u1207  (
    .b({\u2_Display/n3963 [19],\u2_Display/n3963 [22]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3941 ,\u2_Display/n3938 }),
    .f({\u2_Display/n3976 ,\u2_Display/n3973 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1206|_al_u1209  (
    .b({\u2_Display/n3963 [21],\u2_Display/n3963 [24]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3939 ,\u2_Display/n3936 }),
    .f({\u2_Display/n3974 ,\u2_Display/n3971 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100101011001010),
    .MODE("LOGIC"))
    \_al_u1208|_al_u1211  (
    .a({\u2_Display/n3963 [23],open_n2470}),
    .b({\u2_Display/n3937 ,\u2_Display/n3963 [26]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({open_n2473,\u2_Display/n3934 }),
    .f({\u2_Display/n3972 ,\u2_Display/n3969 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1210|_al_u1213  (
    .b({\u2_Display/n3963 [25],\u2_Display/n3963 [28]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3935 ,\u2_Display/n3932 }),
    .f({\u2_Display/n3970 ,\u2_Display/n3967 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1212|_al_u1215  (
    .b({\u2_Display/n3963 [27],\u2_Display/n3963 [30]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3933 ,\u2_Display/n3930 }),
    .f({\u2_Display/n3968 ,\u2_Display/n3965 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1214|_al_u1216  (
    .b({\u2_Display/n3963 [29],\u2_Display/n3963 [31]}),
    .c({\u2_Display/n3961 ,\u2_Display/n3961 }),
    .d({\u2_Display/n3931 ,\u2_Display/n3929 }),
    .f({\u2_Display/n3966 ,\u2_Display/n3964 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1217|_al_u1418  (
    .b({\u2_Display/n5086 [0],\u2_Display/n5121 [31]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6241 ,\u2_Display/n6245 }),
    .f({\u2_Display/n6276 ,\u2_Display/n6280 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1218|_al_u1222  (
    .b({\u2_Display/n5086 [1],\u2_Display/n5086 [5]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6240 ,\u2_Display/n6236 }),
    .f({\u2_Display/n6275 ,\u2_Display/n6271 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .MODE("LOGIC"))
    _al_u1219 (
    .b({open_n2612,\u2_Display/n5086 [2]}),
    .c({open_n2613,\u2_Display/n5084 }),
    .d({open_n2616,\u2_Display/n6239 }),
    .f({open_n2630,\u2_Display/n6274 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1220|_al_u1226  (
    .b({\u2_Display/n5086 [3],\u2_Display/n5086 [9]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6238 ,\u2_Display/n6232 }),
    .f({\u2_Display/n6273 ,\u2_Display/n6267 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1221|_al_u1223  (
    .b({\u2_Display/n5086 [4],\u2_Display/n5086 [6]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6237 ,\u2_Display/n6235 }),
    .f({\u2_Display/n6272 ,\u2_Display/n6270 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1224|_al_u1230  (
    .b({\u2_Display/n5086 [7],\u2_Display/n5086 [13]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6234 ,\u2_Display/n6228 }),
    .f({\u2_Display/n6269 ,\u2_Display/n6263 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1225|_al_u1227  (
    .b({\u2_Display/n5086 [8],\u2_Display/n5086 [10]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6233 ,\u2_Display/n6231 }),
    .f({\u2_Display/n6268 ,\u2_Display/n6266 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1228|_al_u1234  (
    .b({\u2_Display/n5086 [11],\u2_Display/n5086 [17]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6230 ,\u2_Display/n6224 }),
    .f({\u2_Display/n6265 ,\u2_Display/n6259 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1229|_al_u1231  (
    .b({\u2_Display/n5086 [12],\u2_Display/n5086 [14]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6229 ,\u2_Display/n6227 }),
    .f({\u2_Display/n6264 ,\u2_Display/n6262 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1232|_al_u1237  (
    .b({\u2_Display/n5086 [15],\u2_Display/n5086 [20]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6226 ,\u2_Display/n6221 }),
    .f({\u2_Display/n6261 ,\u2_Display/n6256 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1233|_al_u1235  (
    .b({\u2_Display/n5086 [16],\u2_Display/n5086 [18]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6225 ,\u2_Display/n6223 }),
    .f({\u2_Display/n6260 ,\u2_Display/n6258 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1236|_al_u1239  (
    .b({\u2_Display/n5086 [19],\u2_Display/n5086 [22]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6222 ,\u2_Display/n6219 }),
    .f({\u2_Display/n6257 ,\u2_Display/n6254 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1238|_al_u1242  (
    .b({\u2_Display/n5086 [21],\u2_Display/n5086 [25]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6220 ,\u2_Display/n6216 }),
    .f({\u2_Display/n6255 ,\u2_Display/n6251 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1240|_al_u1245  (
    .b({\u2_Display/n5086 [23],\u2_Display/n5086 [28]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6218 ,\u2_Display/n6213 }),
    .f({\u2_Display/n6253 ,\u2_Display/n6248 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1241|_al_u1243  (
    .b({\u2_Display/n5086 [24],\u2_Display/n5086 [26]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6217 ,\u2_Display/n6215 }),
    .f({\u2_Display/n6252 ,\u2_Display/n6250 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1244|_al_u1246  (
    .b({\u2_Display/n5086 [27],\u2_Display/n5086 [29]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6214 ,\u2_Display/n6212 }),
    .f({\u2_Display/n6249 ,\u2_Display/n6247 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1247|_al_u1248  (
    .b({\u2_Display/n5086 [30],\u2_Display/n5086 [31]}),
    .c({\u2_Display/n5084 ,\u2_Display/n5084 }),
    .d({\u2_Display/n6211 ,\u2_Display/n6210 }),
    .f({\u2_Display/n6246 ,\u2_Display/n6245 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1249|_al_u1254  (
    .b({\u2_Display/n594 [0],\u2_Display/n594 [5]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n591 ,\u2_Display/n586 }),
    .f({\u2_Display/n626 ,\u2_Display/n621 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1250|_al_u1251  (
    .b({\u2_Display/n594 [1],\u2_Display/n594 [2]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n590 ,\u2_Display/n589 }),
    .f({\u2_Display/n625 ,\u2_Display/n624 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1252|_al_u1257  (
    .b({\u2_Display/n594 [3],\u2_Display/n594 [8]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n588 ,\u2_Display/n583 }),
    .f({\u2_Display/n623 ,\u2_Display/n618 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1253|_al_u1255  (
    .b({\u2_Display/n594 [4],\u2_Display/n594 [6]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n587 ,\u2_Display/n585 }),
    .f({\u2_Display/n622 ,\u2_Display/n620 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1256|_al_u1259  (
    .b({\u2_Display/n594 [7],\u2_Display/n594 [10]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n584 ,\u2_Display/n581 }),
    .f({\u2_Display/n619 ,\u2_Display/n616 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1258|_al_u1261  (
    .b({\u2_Display/n594 [9],\u2_Display/n594 [12]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n582 ,\u2_Display/n579 }),
    .f({\u2_Display/n617 ,\u2_Display/n614 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1260|_al_u1263  (
    .b({\u2_Display/n594 [11],\u2_Display/n594 [14]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n580 ,\u2_Display/n577 }),
    .f({\u2_Display/n615 ,\u2_Display/n612 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1262|_al_u1265  (
    .b({\u2_Display/n594 [13],\u2_Display/n594 [16]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n578 ,\u2_Display/n575 }),
    .f({\u2_Display/n613 ,\u2_Display/n610 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1264|_al_u1267  (
    .b({\u2_Display/n594 [15],\u2_Display/n594 [18]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n576 ,\u2_Display/n573 }),
    .f({\u2_Display/n611 ,\u2_Display/n608 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1266|_al_u1269  (
    .b({\u2_Display/n594 [17],\u2_Display/n594 [20]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n574 ,\u2_Display/n571 }),
    .f({\u2_Display/n609 ,\u2_Display/n606 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1268|_al_u1271  (
    .b({\u2_Display/n594 [19],\u2_Display/n594 [22]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n572 ,\u2_Display/n569 }),
    .f({\u2_Display/n607 ,\u2_Display/n604 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1270|_al_u1274  (
    .b({\u2_Display/n594 [21],\u2_Display/n594 [25]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n570 ,\u2_Display/n566 }),
    .f({\u2_Display/n605 ,\u2_Display/n601 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1272|_al_u1278  (
    .b({\u2_Display/n594 [23],\u2_Display/n594 [29]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n568 ,\u2_Display/n562 }),
    .f({\u2_Display/n603 ,\u2_Display/n597 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1273|_al_u1275  (
    .b({\u2_Display/n594 [24],\u2_Display/n594 [26]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n567 ,\u2_Display/n565 }),
    .f({\u2_Display/n602 ,\u2_Display/n600 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1276|_al_u1280  (
    .b({\u2_Display/n594 [27],\u2_Display/n594 [31]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n564 ,\u2_Display/n560 }),
    .f({\u2_Display/n599 ,\u2_Display/n595 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1277|_al_u1279  (
    .b({\u2_Display/n594 [28],\u2_Display/n594 [30]}),
    .c({\u2_Display/n592 ,\u2_Display/n592 }),
    .d({\u2_Display/n563 ,\u2_Display/n561 }),
    .f({\u2_Display/n598 ,\u2_Display/n596 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1281|_al_u1285  (
    .b({\u2_Display/n1717 [0],\u2_Display/n1717 [4]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1714 ,\u2_Display/n1710 }),
    .f({\u2_Display/n1749 ,\u2_Display/n1745 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1282|_al_u1283  (
    .b({\u2_Display/n1717 [1],\u2_Display/n1717 [2]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1713 ,\u2_Display/n1712 }),
    .f({\u2_Display/n1748 ,\u2_Display/n1747 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1284|_al_u1287  (
    .b({\u2_Display/n1717 [3],\u2_Display/n1717 [6]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1711 ,\u2_Display/n1708 }),
    .f({\u2_Display/n1746 ,\u2_Display/n1743 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1286|_al_u1289  (
    .b({\u2_Display/n1717 [5],\u2_Display/n1717 [8]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1709 ,\u2_Display/n1706 }),
    .f({\u2_Display/n1744 ,\u2_Display/n1741 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1288|_al_u1291  (
    .b({\u2_Display/n1717 [7],\u2_Display/n1717 [10]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1707 ,\u2_Display/n1704 }),
    .f({\u2_Display/n1742 ,\u2_Display/n1739 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1290|_al_u1293  (
    .b({\u2_Display/n1717 [9],\u2_Display/n1717 [12]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1705 ,\u2_Display/n1702 }),
    .f({\u2_Display/n1740 ,\u2_Display/n1737 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1292|_al_u1295  (
    .b({\u2_Display/n1717 [11],\u2_Display/n1717 [14]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1703 ,\u2_Display/n1700 }),
    .f({\u2_Display/n1738 ,\u2_Display/n1735 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1294|_al_u1297  (
    .b({\u2_Display/n1717 [13],\u2_Display/n1717 [16]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1701 ,\u2_Display/n1698 }),
    .f({\u2_Display/n1736 ,\u2_Display/n1733 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1296|_al_u1299  (
    .b({\u2_Display/n1717 [15],\u2_Display/n1717 [18]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1699 ,\u2_Display/n1696 }),
    .f({\u2_Display/n1734 ,\u2_Display/n1731 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1298|_al_u1302  (
    .b({\u2_Display/n1717 [17],\u2_Display/n1717 [21]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1697 ,\u2_Display/n1693 }),
    .f({\u2_Display/n1732 ,\u2_Display/n1728 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1300|_al_u1305  (
    .b({\u2_Display/n1717 [19],\u2_Display/n1717 [24]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1695 ,\u2_Display/n1690 }),
    .f({\u2_Display/n1730 ,\u2_Display/n1725 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1301|_al_u1303  (
    .b({\u2_Display/n1717 [20],\u2_Display/n1717 [22]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1694 ,\u2_Display/n1692 }),
    .f({\u2_Display/n1729 ,\u2_Display/n1727 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1304|_al_u1307  (
    .b({\u2_Display/n1717 [23],\u2_Display/n1717 [26]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1691 ,\u2_Display/n1688 }),
    .f({\u2_Display/n1726 ,\u2_Display/n1723 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1306|_al_u1310  (
    .b({\u2_Display/n1717 [25],\u2_Display/n1717 [29]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1689 ,\u2_Display/n1685 }),
    .f({\u2_Display/n1724 ,\u2_Display/n1720 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1308|_al_u1312  (
    .b({\u2_Display/n1717 [27],\u2_Display/n1717 [31]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1687 ,\u2_Display/n1683 }),
    .f({\u2_Display/n1722 ,\u2_Display/n1718 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1309|_al_u1311  (
    .b({\u2_Display/n1717 [28],\u2_Display/n1717 [30]}),
    .c({\u2_Display/n1715 ,\u2_Display/n1715 }),
    .d({\u2_Display/n1686 ,\u2_Display/n1684 }),
    .f({\u2_Display/n1721 ,\u2_Display/n1719 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1313|_al_u1315  (
    .b({\u2_Display/n2840 [0],\u2_Display/n2840 [2]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2837 ,\u2_Display/n2835 }),
    .f({\u2_Display/n2872 ,\u2_Display/n2870 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .MODE("LOGIC"))
    _al_u1314 (
    .b({open_n3768,\u2_Display/n2840 [1]}),
    .c({open_n3769,\u2_Display/n2838 }),
    .d({open_n3772,\u2_Display/n2836 }),
    .f({open_n3786,\u2_Display/n2871 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1316|_al_u1317  (
    .b({\u2_Display/n2840 [3],\u2_Display/n2840 [4]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2834 ,\u2_Display/n2833 }),
    .f({\u2_Display/n2869 ,\u2_Display/n2868 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1318|_al_u1319  (
    .b({\u2_Display/n2840 [5],\u2_Display/n2840 [6]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2832 ,\u2_Display/n2831 }),
    .f({\u2_Display/n2867 ,\u2_Display/n2866 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1320|_al_u1321  (
    .b({\u2_Display/n2840 [7],\u2_Display/n2840 [8]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2830 ,\u2_Display/n2829 }),
    .f({\u2_Display/n2865 ,\u2_Display/n2864 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1322|_al_u1323  (
    .b({\u2_Display/n2840 [9],\u2_Display/n2840 [10]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2828 ,\u2_Display/n2827 }),
    .f({\u2_Display/n2863 ,\u2_Display/n2862 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1324|_al_u1325  (
    .b({\u2_Display/n2840 [11],\u2_Display/n2840 [12]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2826 ,\u2_Display/n2825 }),
    .f({\u2_Display/n2861 ,\u2_Display/n2860 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1326|_al_u1327  (
    .b({\u2_Display/n2840 [13],\u2_Display/n2840 [14]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2824 ,\u2_Display/n2823 }),
    .f({\u2_Display/n2859 ,\u2_Display/n2858 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100101011001010),
    .MODE("LOGIC"))
    \_al_u1328|_al_u1331  (
    .a({\u2_Display/n2840 [15],open_n3940}),
    .b({\u2_Display/n2822 ,\u2_Display/n2840 [18]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({open_n3943,\u2_Display/n2819 }),
    .f({\u2_Display/n2857 ,\u2_Display/n2854 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000110000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1329|_al_u1330  (
    .b({\u2_Display/n2840 [16],\u2_Display/n2838 }),
    .c({\u2_Display/n2838 ,\u2_Display/n2840 [17]}),
    .d({\u2_Display/n2821 ,\u2_Display/n2820 }),
    .f({\u2_Display/n2856 ,\u2_Display/n2855 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1332|_al_u1333  (
    .b({\u2_Display/n2840 [19],\u2_Display/n2840 [20]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2818 ,\u2_Display/n2817 }),
    .f({\u2_Display/n2853 ,\u2_Display/n2852 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1334|_al_u1335  (
    .b({\u2_Display/n2840 [21],\u2_Display/n2840 [22]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2816 ,\u2_Display/n2815 }),
    .f({\u2_Display/n2851 ,\u2_Display/n2850 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111101000001010),
    .MODE("LOGIC"))
    \_al_u1336|_al_u1339  (
    .a({\u2_Display/n2840 [23],open_n4036}),
    .b({open_n4037,\u2_Display/n2840 [26]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2814 ,\u2_Display/n2811 }),
    .f({\u2_Display/n2849 ,\u2_Display/n2846 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1337|_al_u1338  (
    .b({\u2_Display/n2840 [24],\u2_Display/n2840 [25]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2813 ,\u2_Display/n2812 }),
    .f({\u2_Display/n2848 ,\u2_Display/n2847 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1340|_al_u1343  (
    .b({\u2_Display/n2840 [27],\u2_Display/n2840 [30]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2810 ,\u2_Display/n2807 }),
    .f({\u2_Display/n2845 ,\u2_Display/n2842 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1341|_al_u1342  (
    .b({\u2_Display/n2840 [28],\u2_Display/n2840 [29]}),
    .c({\u2_Display/n2838 ,\u2_Display/n2838 }),
    .d({\u2_Display/n2809 ,\u2_Display/n2808 }),
    .f({\u2_Display/n2844 ,\u2_Display/n2843 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1355|_al_u1357  (
    .b({\u2_Display/n3998 [0],\u2_Display/n3998 [2]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3995 ,\u2_Display/n3993 }),
    .f({\u2_Display/n4030 ,\u2_Display/n4028 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1356|_al_u1360  (
    .b({\u2_Display/n3998 [1],\u2_Display/n3998 [5]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3994 ,\u2_Display/n3990 }),
    .f({\u2_Display/n4029 ,\u2_Display/n4025 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u1358|_al_u1364  (
    .b({\u2_Display/n3992 ,\u2_Display/n3998 [9]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3998 [3],\u2_Display/n3986 }),
    .f({\u2_Display/n4027 ,\u2_Display/n4021 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1359|_al_u1361  (
    .b({\u2_Display/n3998 [4],\u2_Display/n3998 [6]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3991 ,\u2_Display/n3989 }),
    .f({\u2_Display/n4026 ,\u2_Display/n4024 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1362|_al_u1367  (
    .b({\u2_Display/n3998 [7],\u2_Display/n3998 [12]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3988 ,\u2_Display/n3983 }),
    .f({\u2_Display/n4023 ,\u2_Display/n4018 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1363|_al_u1365  (
    .b({\u2_Display/n3998 [8],\u2_Display/n3998 [10]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3987 ,\u2_Display/n3985 }),
    .f({\u2_Display/n4022 ,\u2_Display/n4020 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1366|_al_u1369  (
    .b({\u2_Display/n3998 [11],\u2_Display/n3998 [14]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3984 ,\u2_Display/n3981 }),
    .f({\u2_Display/n4019 ,\u2_Display/n4016 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1368|_al_u1371  (
    .b({\u2_Display/n3998 [13],\u2_Display/n3998 [16]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3982 ,\u2_Display/n3979 }),
    .f({\u2_Display/n4017 ,\u2_Display/n4014 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1370|_al_u1373  (
    .b({\u2_Display/n3998 [15],\u2_Display/n3998 [18]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3980 ,\u2_Display/n3977 }),
    .f({\u2_Display/n4015 ,\u2_Display/n4012 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1372|_al_u1376  (
    .b({\u2_Display/n3998 [17],\u2_Display/n3998 [21]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3978 ,\u2_Display/n3974 }),
    .f({\u2_Display/n4013 ,\u2_Display/n4009 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1374|_al_u1380  (
    .b({\u2_Display/n3998 [19],\u2_Display/n3998 [25]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3976 ,\u2_Display/n3970 }),
    .f({\u2_Display/n4011 ,\u2_Display/n4005 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1375|_al_u1377  (
    .b({\u2_Display/n3998 [20],\u2_Display/n3998 [22]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3975 ,\u2_Display/n3973 }),
    .f({\u2_Display/n4010 ,\u2_Display/n4008 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1378|_al_u1383  (
    .b({\u2_Display/n3998 [23],\u2_Display/n3998 [28]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3972 ,\u2_Display/n3967 }),
    .f({\u2_Display/n4007 ,\u2_Display/n4002 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1379|_al_u1381  (
    .b({\u2_Display/n3998 [24],\u2_Display/n3998 [26]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3971 ,\u2_Display/n3969 }),
    .f({\u2_Display/n4006 ,\u2_Display/n4004 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1382|_al_u1385  (
    .b({\u2_Display/n3998 [27],\u2_Display/n3998 [30]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3968 ,\u2_Display/n3965 }),
    .f({\u2_Display/n4003 ,\u2_Display/n4000 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1384|_al_u1386  (
    .b({\u2_Display/n3998 [29],\u2_Display/n3998 [31]}),
    .c({\u2_Display/n3996 ,\u2_Display/n3996 }),
    .d({\u2_Display/n3966 ,\u2_Display/n3964 }),
    .f({\u2_Display/n4001 ,\u2_Display/n3999 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .MODE("LOGIC"))
    _al_u1387 (
    .b({open_n4518,\u2_Display/n5121 [0]}),
    .c({open_n4519,\u2_Display/n5119 }),
    .d({open_n4522,\u2_Display/n6276 }),
    .f({open_n4536,\u2_Display/n6311 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1388|_al_u1389  (
    .b({\u2_Display/n5121 [1],\u2_Display/n5121 [2]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6275 ,\u2_Display/n6274 }),
    .f({\u2_Display/n6310 ,\u2_Display/n6309 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1390|_al_u1393  (
    .b({\u2_Display/n5121 [3],\u2_Display/n5121 [6]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6273 ,\u2_Display/n6270 }),
    .f({\u2_Display/n6308 ,\u2_Display/n6305 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1391|_al_u1392  (
    .b({\u2_Display/n5121 [4],\u2_Display/n5121 [5]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6272 ,\u2_Display/n6271 }),
    .f({\u2_Display/n6307 ,\u2_Display/n6306 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1394|_al_u1397  (
    .b({\u2_Display/n5121 [7],\u2_Display/n5121 [10]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6269 ,\u2_Display/n6266 }),
    .f({\u2_Display/n6304 ,\u2_Display/n6301 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1395|_al_u1396  (
    .b({\u2_Display/n5121 [8],\u2_Display/n5121 [9]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6268 ,\u2_Display/n6267 }),
    .f({\u2_Display/n6303 ,\u2_Display/n6302 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1398|_al_u1401  (
    .b({\u2_Display/n5121 [11],\u2_Display/n5121 [14]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6265 ,\u2_Display/n6262 }),
    .f({\u2_Display/n6300 ,\u2_Display/n6297 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1399|_al_u1400  (
    .b({\u2_Display/n5121 [12],\u2_Display/n5121 [13]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6264 ,\u2_Display/n6263 }),
    .f({\u2_Display/n6299 ,\u2_Display/n6298 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1402|_al_u1405  (
    .b({\u2_Display/n5121 [15],\u2_Display/n5121 [18]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6261 ,\u2_Display/n6258 }),
    .f({\u2_Display/n6296 ,\u2_Display/n6293 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1403|_al_u1404  (
    .b({\u2_Display/n5121 [16],\u2_Display/n5121 [17]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6260 ,\u2_Display/n6259 }),
    .f({\u2_Display/n6295 ,\u2_Display/n6294 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1406|_al_u1409  (
    .b({\u2_Display/n5121 [19],\u2_Display/n5121 [22]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6257 ,\u2_Display/n6254 }),
    .f({\u2_Display/n6292 ,\u2_Display/n6289 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1407|_al_u1408  (
    .b({\u2_Display/n5121 [20],\u2_Display/n5121 [21]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6256 ,\u2_Display/n6255 }),
    .f({\u2_Display/n6291 ,\u2_Display/n6290 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1410|_al_u1413  (
    .b({\u2_Display/n5121 [23],\u2_Display/n5121 [26]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6253 ,\u2_Display/n6250 }),
    .f({\u2_Display/n6288 ,\u2_Display/n6285 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1411|_al_u1412  (
    .b({\u2_Display/n5121 [24],\u2_Display/n5121 [25]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6252 ,\u2_Display/n6251 }),
    .f({\u2_Display/n6287 ,\u2_Display/n6286 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1414|_al_u1417  (
    .b({\u2_Display/n5121 [27],\u2_Display/n5121 [30]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6249 ,\u2_Display/n6246 }),
    .f({\u2_Display/n6284 ,\u2_Display/n6281 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1415|_al_u1416  (
    .b({\u2_Display/n5121 [28],\u2_Display/n5121 [29]}),
    .c({\u2_Display/n5119 ,\u2_Display/n5119 }),
    .d({\u2_Display/n6248 ,\u2_Display/n6247 }),
    .f({\u2_Display/n6283 ,\u2_Display/n6282 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1419|_al_u1424  (
    .b({\u2_Display/n629 [0],\u2_Display/n629 [5]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n626 ,\u2_Display/n621 }),
    .f({\u2_Display/n661 ,\u2_Display/n656 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1420|_al_u1421  (
    .b({\u2_Display/n629 [1],\u2_Display/n629 [2]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n625 ,\u2_Display/n624 }),
    .f({\u2_Display/n660 ,\u2_Display/n659 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1422|_al_u1428  (
    .b({\u2_Display/n629 [3],\u2_Display/n629 [9]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n623 ,\u2_Display/n617 }),
    .f({\u2_Display/n658 ,\u2_Display/n652 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1423|_al_u1425  (
    .b({\u2_Display/n629 [4],\u2_Display/n629 [6]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n622 ,\u2_Display/n620 }),
    .f({\u2_Display/n657 ,\u2_Display/n655 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1426|_al_u1431  (
    .b({\u2_Display/n629 [7],\u2_Display/n629 [12]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n619 ,\u2_Display/n614 }),
    .f({\u2_Display/n654 ,\u2_Display/n649 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1427|_al_u1429  (
    .b({\u2_Display/n629 [8],\u2_Display/n629 [10]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n618 ,\u2_Display/n616 }),
    .f({\u2_Display/n653 ,\u2_Display/n651 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1430|_al_u1433  (
    .b({\u2_Display/n629 [11],\u2_Display/n629 [14]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n615 ,\u2_Display/n612 }),
    .f({\u2_Display/n650 ,\u2_Display/n647 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1432|_al_u1436  (
    .b({\u2_Display/n629 [13],\u2_Display/n629 [17]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n613 ,\u2_Display/n609 }),
    .f({\u2_Display/n648 ,\u2_Display/n644 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1434|_al_u1440  (
    .b({\u2_Display/n629 [15],\u2_Display/n629 [21]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n611 ,\u2_Display/n605 }),
    .f({\u2_Display/n646 ,\u2_Display/n640 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1435|_al_u1437  (
    .b({\u2_Display/n629 [16],\u2_Display/n629 [18]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n610 ,\u2_Display/n608 }),
    .f({\u2_Display/n645 ,\u2_Display/n643 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1438|_al_u1444  (
    .b({\u2_Display/n629 [19],\u2_Display/n629 [25]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n607 ,\u2_Display/n601 }),
    .f({\u2_Display/n642 ,\u2_Display/n636 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1439|_al_u1441  (
    .b({\u2_Display/n629 [20],\u2_Display/n629 [22]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n606 ,\u2_Display/n604 }),
    .f({\u2_Display/n641 ,\u2_Display/n639 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1442|_al_u1447  (
    .b({\u2_Display/n629 [23],\u2_Display/n629 [28]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n603 ,\u2_Display/n598 }),
    .f({\u2_Display/n638 ,\u2_Display/n633 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1443|_al_u1445  (
    .b({\u2_Display/n629 [24],\u2_Display/n629 [26]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n602 ,\u2_Display/n600 }),
    .f({\u2_Display/n637 ,\u2_Display/n635 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1446|_al_u1449  (
    .b({\u2_Display/n629 [27],\u2_Display/n629 [30]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n599 ,\u2_Display/n596 }),
    .f({\u2_Display/n634 ,\u2_Display/n631 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1448|_al_u1450  (
    .b({\u2_Display/n629 [29],\u2_Display/n629 [31]}),
    .c({\u2_Display/n627 ,\u2_Display/n627 }),
    .d({\u2_Display/n597 ,\u2_Display/n595 }),
    .f({\u2_Display/n632 ,\u2_Display/n630 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1451|_al_u1456  (
    .b({\u2_Display/n1752 [0],\u2_Display/n1752 [5]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1749 ,\u2_Display/n1744 }),
    .f({\u2_Display/n1784 ,\u2_Display/n1779 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1452|_al_u1453  (
    .b({\u2_Display/n1752 [1],\u2_Display/n1752 [2]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1748 ,\u2_Display/n1747 }),
    .f({\u2_Display/n1783 ,\u2_Display/n1782 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u1454|_al_u1459  (
    .b({\u2_Display/n1750 ,\u2_Display/n1752 [8]}),
    .c({\u2_Display/n1752 [3],\u2_Display/n1750 }),
    .d({\u2_Display/n1746 ,\u2_Display/n1741 }),
    .f({\u2_Display/n1781 ,\u2_Display/n1776 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1455|_al_u1457  (
    .b({\u2_Display/n1752 [4],\u2_Display/n1752 [6]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1745 ,\u2_Display/n1743 }),
    .f({\u2_Display/n1780 ,\u2_Display/n1778 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1458|_al_u1461  (
    .b({\u2_Display/n1752 [7],\u2_Display/n1752 [10]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1742 ,\u2_Display/n1739 }),
    .f({\u2_Display/n1777 ,\u2_Display/n1774 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1460|_al_u1463  (
    .b({\u2_Display/n1752 [9],\u2_Display/n1752 [12]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1740 ,\u2_Display/n1737 }),
    .f({\u2_Display/n1775 ,\u2_Display/n1772 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u1462|_al_u1465  (
    .b({\u2_Display/n1738 ,\u2_Display/n1752 [14]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1752 [11],\u2_Display/n1735 }),
    .f({\u2_Display/n1773 ,\u2_Display/n1770 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1464|_al_u1467  (
    .b({\u2_Display/n1752 [13],\u2_Display/n1752 [16]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1736 ,\u2_Display/n1733 }),
    .f({\u2_Display/n1771 ,\u2_Display/n1768 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1466|_al_u902  (
    .b({\u2_Display/n1752 [15],\u2_Display/n524 [1]}),
    .c({\u2_Display/n1750 ,\u2_Display/n522 }),
    .d({\u2_Display/n1734 ,\u2_Display/n520 }),
    .f({\u2_Display/n1769 ,\u2_Display/n555 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1468|_al_u1469  (
    .b({\u2_Display/n1752 [17],\u2_Display/n1752 [18]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1732 ,\u2_Display/n1731 }),
    .f({\u2_Display/n1767 ,\u2_Display/n1766 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1470|_al_u1471  (
    .b({\u2_Display/n1752 [19],\u2_Display/n1752 [20]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1730 ,\u2_Display/n1729 }),
    .f({\u2_Display/n1765 ,\u2_Display/n1764 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1472|_al_u1473  (
    .b({\u2_Display/n1752 [21],\u2_Display/n1752 [22]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1728 ,\u2_Display/n1727 }),
    .f({\u2_Display/n1763 ,\u2_Display/n1762 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1474|_al_u1477  (
    .b({\u2_Display/n1752 [23],\u2_Display/n1752 [26]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1726 ,\u2_Display/n1723 }),
    .f({\u2_Display/n1761 ,\u2_Display/n1758 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1475|_al_u1476  (
    .b({\u2_Display/n1752 [24],\u2_Display/n1752 [25]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1725 ,\u2_Display/n1724 }),
    .f({\u2_Display/n1760 ,\u2_Display/n1759 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1478|_al_u1479  (
    .b({\u2_Display/n1752 [27],\u2_Display/n1752 [28]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1722 ,\u2_Display/n1721 }),
    .f({\u2_Display/n1757 ,\u2_Display/n1756 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1480|_al_u1481  (
    .b({\u2_Display/n1752 [29],\u2_Display/n1752 [30]}),
    .c({\u2_Display/n1750 ,\u2_Display/n1750 }),
    .d({\u2_Display/n1720 ,\u2_Display/n1719 }),
    .f({\u2_Display/n1755 ,\u2_Display/n1754 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1482|_al_u918  (
    .b({\u2_Display/n1752 [31],\u2_Display/n524 [17]}),
    .c({\u2_Display/n1750 ,\u2_Display/n522 }),
    .d({\u2_Display/n1718 ,\u2_Display/n504 }),
    .f({\u2_Display/n1753 ,\u2_Display/n539 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1483|_al_u1485  (
    .b({\u2_Display/n2875 [0],\u2_Display/n2875 [2]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2872 ,\u2_Display/n2870 }),
    .f({\u2_Display/n2907 ,\u2_Display/n2905 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .MODE("LOGIC"))
    _al_u1484 (
    .b({open_n5730,\u2_Display/n2875 [1]}),
    .c({open_n5731,\u2_Display/n2873 }),
    .d({open_n5734,\u2_Display/n2871 }),
    .f({open_n5748,\u2_Display/n2906 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1486|_al_u1489  (
    .b({\u2_Display/n2875 [3],\u2_Display/n2875 [6]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2869 ,\u2_Display/n2866 }),
    .f({\u2_Display/n2904 ,\u2_Display/n2901 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1487|_al_u1488  (
    .b({\u2_Display/n2875 [4],\u2_Display/n2875 [5]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2868 ,\u2_Display/n2867 }),
    .f({\u2_Display/n2903 ,\u2_Display/n2902 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1490|_al_u1493  (
    .b({\u2_Display/n2875 [7],\u2_Display/n2875 [10]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2865 ,\u2_Display/n2862 }),
    .f({\u2_Display/n2900 ,\u2_Display/n2897 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1491|_al_u1492  (
    .b({\u2_Display/n2875 [8],\u2_Display/n2875 [9]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2864 ,\u2_Display/n2863 }),
    .f({\u2_Display/n2899 ,\u2_Display/n2898 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1494|_al_u1497  (
    .b({\u2_Display/n2875 [11],\u2_Display/n2875 [14]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2861 ,\u2_Display/n2858 }),
    .f({\u2_Display/n2896 ,\u2_Display/n2893 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1495|_al_u1496  (
    .b({\u2_Display/n2875 [12],\u2_Display/n2875 [13]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2860 ,\u2_Display/n2859 }),
    .f({\u2_Display/n2895 ,\u2_Display/n2894 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1498|_al_u1499  (
    .b({\u2_Display/n2875 [15],\u2_Display/n2875 [16]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2857 ,\u2_Display/n2856 }),
    .f({\u2_Display/n2892 ,\u2_Display/n2891 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1500|_al_u1501  (
    .b({\u2_Display/n2875 [17],\u2_Display/n2875 [18]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2855 ,\u2_Display/n2854 }),
    .f({\u2_Display/n2890 ,\u2_Display/n2889 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1502|_al_u1505  (
    .b({\u2_Display/n2875 [19],\u2_Display/n2875 [22]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2853 ,\u2_Display/n2850 }),
    .f({\u2_Display/n2888 ,\u2_Display/n2885 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1503|_al_u1504  (
    .b({\u2_Display/n2875 [20],\u2_Display/n2875 [21]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2852 ,\u2_Display/n2851 }),
    .f({\u2_Display/n2887 ,\u2_Display/n2886 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1506|_al_u1509  (
    .b({\u2_Display/n2875 [23],\u2_Display/n2875 [26]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2849 ,\u2_Display/n2846 }),
    .f({\u2_Display/n2884 ,\u2_Display/n2881 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1507|_al_u1508  (
    .b({\u2_Display/n2875 [24],\u2_Display/n2875 [25]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2848 ,\u2_Display/n2847 }),
    .f({\u2_Display/n2883 ,\u2_Display/n2882 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1510|_al_u1511  (
    .b({\u2_Display/n2875 [27],\u2_Display/n2875 [28]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2845 ,\u2_Display/n2844 }),
    .f({\u2_Display/n2880 ,\u2_Display/n2879 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1512|_al_u1513  (
    .b({\u2_Display/n2875 [29],\u2_Display/n2875 [30]}),
    .c({\u2_Display/n2873 ,\u2_Display/n2873 }),
    .d({\u2_Display/n2843 ,\u2_Display/n2842 }),
    .f({\u2_Display/n2878 ,\u2_Display/n2877 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(~D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000000011111111),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0000000011111111),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1514|_al_u4000  (
    .b({\u2_Display/n2875 [31],open_n6092}),
    .c({\u2_Display/n2873 ,open_n6093}),
    .d({\u2_Display/n2841 ,clk_vga}),
    .f({\u2_Display/n2876 ,vga_clk_pad}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1515|_al_u1519  (
    .b({\u2_Display/n4033 [0],\u2_Display/n4033 [4]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4030 ,\u2_Display/n4026 }),
    .f({\u2_Display/n4065 ,\u2_Display/n4061 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1516|_al_u1517  (
    .b({\u2_Display/n4033 [1],\u2_Display/n4033 [2]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4029 ,\u2_Display/n4028 }),
    .f({\u2_Display/n4064 ,\u2_Display/n4063 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1518|_al_u1521  (
    .b({\u2_Display/n4033 [3],\u2_Display/n4033 [6]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4027 ,\u2_Display/n4024 }),
    .f({\u2_Display/n4062 ,\u2_Display/n4059 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1520|_al_u1524  (
    .b({\u2_Display/n4033 [5],\u2_Display/n4033 [9]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4025 ,\u2_Display/n4021 }),
    .f({\u2_Display/n4060 ,\u2_Display/n4056 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1522|_al_u1528  (
    .b({\u2_Display/n4033 [7],\u2_Display/n4033 [13]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4023 ,\u2_Display/n4017 }),
    .f({\u2_Display/n4058 ,\u2_Display/n4052 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1523|_al_u1525  (
    .b({\u2_Display/n4033 [8],\u2_Display/n4033 [10]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4022 ,\u2_Display/n4020 }),
    .f({\u2_Display/n4057 ,\u2_Display/n4055 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1526|_al_u1531  (
    .b({\u2_Display/n4033 [11],\u2_Display/n4033 [16]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4019 ,\u2_Display/n4014 }),
    .f({\u2_Display/n4054 ,\u2_Display/n4049 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1527|_al_u1529  (
    .b({\u2_Display/n4033 [12],\u2_Display/n4033 [14]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4018 ,\u2_Display/n4016 }),
    .f({\u2_Display/n4053 ,\u2_Display/n4051 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1530|_al_u1533  (
    .b({\u2_Display/n4033 [15],\u2_Display/n4033 [18]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4015 ,\u2_Display/n4012 }),
    .f({\u2_Display/n4050 ,\u2_Display/n4047 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1532|_al_u1535  (
    .b({\u2_Display/n4033 [17],\u2_Display/n4033 [20]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4013 ,\u2_Display/n4010 }),
    .f({\u2_Display/n4048 ,\u2_Display/n4045 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1534|_al_u1537  (
    .b({\u2_Display/n4033 [19],\u2_Display/n4033 [22]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4011 ,\u2_Display/n4008 }),
    .f({\u2_Display/n4046 ,\u2_Display/n4043 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1536|_al_u1539  (
    .b({\u2_Display/n4033 [21],\u2_Display/n4033 [24]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4009 ,\u2_Display/n4006 }),
    .f({\u2_Display/n4044 ,\u2_Display/n4041 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1538|_al_u1541  (
    .b({\u2_Display/n4033 [23],\u2_Display/n4033 [26]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4007 ,\u2_Display/n4004 }),
    .f({\u2_Display/n4042 ,\u2_Display/n4039 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1540|_al_u1543  (
    .b({\u2_Display/n4033 [25],\u2_Display/n4033 [28]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4005 ,\u2_Display/n4002 }),
    .f({\u2_Display/n4040 ,\u2_Display/n4037 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1542|_al_u1545  (
    .b({\u2_Display/n4033 [27],\u2_Display/n4033 [30]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4003 ,\u2_Display/n4000 }),
    .f({\u2_Display/n4038 ,\u2_Display/n4035 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1544|_al_u1546  (
    .b({\u2_Display/n4033 [29],\u2_Display/n4033 [31]}),
    .c({\u2_Display/n4031 ,\u2_Display/n4031 }),
    .d({\u2_Display/n4001 ,\u2_Display/n3999 }),
    .f({\u2_Display/n4036 ,\u2_Display/n4034 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1547|_al_u1549  (
    .b({\u2_Display/n5156 [0],\u2_Display/n5156 [2]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6311 ,\u2_Display/n6309 }),
    .f({\u2_Display/n6346 ,\u2_Display/n6344 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1548|_al_u1552  (
    .b({\u2_Display/n5156 [1],\u2_Display/n5156 [5]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6310 ,\u2_Display/n6306 }),
    .f({\u2_Display/n6345 ,\u2_Display/n6341 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1550|_al_u1556  (
    .b({\u2_Display/n5156 [3],\u2_Display/n5156 [9]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6308 ,\u2_Display/n6302 }),
    .f({\u2_Display/n6343 ,\u2_Display/n6337 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1551|_al_u1553  (
    .b({\u2_Display/n5156 [4],\u2_Display/n5156 [6]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6307 ,\u2_Display/n6305 }),
    .f({\u2_Display/n6342 ,\u2_Display/n6340 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1554|_al_u1559  (
    .b({\u2_Display/n5156 [7],\u2_Display/n5156 [12]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6304 ,\u2_Display/n6299 }),
    .f({\u2_Display/n6339 ,\u2_Display/n6334 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1555|_al_u1557  (
    .b({\u2_Display/n5156 [8],\u2_Display/n5156 [10]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6303 ,\u2_Display/n6301 }),
    .f({\u2_Display/n6338 ,\u2_Display/n6336 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1558|_al_u1561  (
    .b({\u2_Display/n5156 [11],\u2_Display/n5156 [14]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6300 ,\u2_Display/n6297 }),
    .f({\u2_Display/n6335 ,\u2_Display/n6332 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100101011001010),
    .MODE("LOGIC"))
    \_al_u1560|_al_u1564  (
    .a({\u2_Display/n5156 [13],open_n6672}),
    .b({\u2_Display/n6298 ,\u2_Display/n5156 [17]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({open_n6675,\u2_Display/n6294 }),
    .f({\u2_Display/n6333 ,\u2_Display/n6329 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1562|_al_u1567  (
    .b({\u2_Display/n5156 [15],\u2_Display/n5156 [20]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6296 ,\u2_Display/n6291 }),
    .f({\u2_Display/n6331 ,\u2_Display/n6326 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1563|_al_u1565  (
    .b({\u2_Display/n5156 [16],\u2_Display/n5156 [18]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6295 ,\u2_Display/n6293 }),
    .f({\u2_Display/n6330 ,\u2_Display/n6328 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1566|_al_u1569  (
    .b({\u2_Display/n5156 [19],\u2_Display/n5156 [22]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6292 ,\u2_Display/n6289 }),
    .f({\u2_Display/n6327 ,\u2_Display/n6324 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1568|_al_u1571  (
    .b({\u2_Display/n5156 [21],\u2_Display/n5156 [24]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6290 ,\u2_Display/n6287 }),
    .f({\u2_Display/n6325 ,\u2_Display/n6322 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1570|_al_u1573  (
    .b({\u2_Display/n5156 [23],\u2_Display/n5156 [26]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6288 ,\u2_Display/n6285 }),
    .f({\u2_Display/n6323 ,\u2_Display/n6320 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1572|_al_u1575  (
    .b({\u2_Display/n5156 [25],\u2_Display/n5156 [28]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6286 ,\u2_Display/n6283 }),
    .f({\u2_Display/n6321 ,\u2_Display/n6318 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1574|_al_u1577  (
    .b({\u2_Display/n5156 [27],\u2_Display/n5156 [30]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6284 ,\u2_Display/n6281 }),
    .f({\u2_Display/n6319 ,\u2_Display/n6316 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1576|_al_u1578  (
    .b({\u2_Display/n5156 [29],\u2_Display/n5156 [31]}),
    .c({\u2_Display/n5154 ,\u2_Display/n5154 }),
    .d({\u2_Display/n6282 ,\u2_Display/n6280 }),
    .f({\u2_Display/n6317 ,\u2_Display/n6315 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1579|_al_u1581  (
    .b({\u2_Display/n664 [0],\u2_Display/n664 [2]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n661 ,\u2_Display/n659 }),
    .f({\u2_Display/n696 ,\u2_Display/n694 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1580|_al_u1584  (
    .b({\u2_Display/n664 [1],\u2_Display/n664 [5]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n660 ,\u2_Display/n656 }),
    .f({\u2_Display/n695 ,\u2_Display/n691 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u1582|_al_u1588  (
    .b({\u2_Display/n658 ,\u2_Display/n664 [9]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n664 [3],\u2_Display/n652 }),
    .f({\u2_Display/n693 ,\u2_Display/n687 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1583|_al_u1585  (
    .b({\u2_Display/n664 [4],\u2_Display/n664 [6]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n657 ,\u2_Display/n655 }),
    .f({\u2_Display/n692 ,\u2_Display/n690 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1586|_al_u1592  (
    .b({\u2_Display/n664 [7],\u2_Display/n664 [13]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n654 ,\u2_Display/n648 }),
    .f({\u2_Display/n689 ,\u2_Display/n683 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1587|_al_u1589  (
    .b({\u2_Display/n664 [8],\u2_Display/n664 [10]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n653 ,\u2_Display/n651 }),
    .f({\u2_Display/n688 ,\u2_Display/n686 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u1590|_al_u1596  (
    .b({\u2_Display/n662 ,\u2_Display/n664 [17]}),
    .c({\u2_Display/n664 [11],\u2_Display/n662 }),
    .d({\u2_Display/n650 ,\u2_Display/n644 }),
    .f({\u2_Display/n685 ,\u2_Display/n679 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1591|_al_u1593  (
    .b({\u2_Display/n664 [12],\u2_Display/n664 [14]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n649 ,\u2_Display/n647 }),
    .f({\u2_Display/n684 ,\u2_Display/n682 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1594|_al_u1600  (
    .b({\u2_Display/n664 [15],\u2_Display/n664 [21]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n646 ,\u2_Display/n640 }),
    .f({\u2_Display/n681 ,\u2_Display/n675 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1595|_al_u1597  (
    .b({\u2_Display/n664 [16],\u2_Display/n664 [18]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n645 ,\u2_Display/n643 }),
    .f({\u2_Display/n680 ,\u2_Display/n678 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u1598|_al_u1604  (
    .b({\u2_Display/n662 ,\u2_Display/n664 [25]}),
    .c({\u2_Display/n664 [19],\u2_Display/n662 }),
    .d({\u2_Display/n642 ,\u2_Display/n636 }),
    .f({\u2_Display/n677 ,\u2_Display/n671 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1599|_al_u1601  (
    .b({\u2_Display/n664 [20],\u2_Display/n664 [22]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n641 ,\u2_Display/n639 }),
    .f({\u2_Display/n676 ,\u2_Display/n674 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1602|_al_u1608  (
    .b({\u2_Display/n664 [23],\u2_Display/n664 [29]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n638 ,\u2_Display/n632 }),
    .f({\u2_Display/n673 ,\u2_Display/n667 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1603|_al_u1605  (
    .b({\u2_Display/n664 [24],\u2_Display/n664 [26]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n637 ,\u2_Display/n635 }),
    .f({\u2_Display/n672 ,\u2_Display/n670 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1606|_al_u1610  (
    .b({\u2_Display/n664 [27],\u2_Display/n664 [31]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n634 ,\u2_Display/n630 }),
    .f({\u2_Display/n669 ,\u2_Display/n665 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1607|_al_u1609  (
    .b({\u2_Display/n664 [28],\u2_Display/n664 [30]}),
    .c({\u2_Display/n662 ,\u2_Display/n662 }),
    .d({\u2_Display/n633 ,\u2_Display/n631 }),
    .f({\u2_Display/n668 ,\u2_Display/n666 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .MODE("LOGIC"))
    _al_u1611 (
    .b({open_n7272,\u2_Display/n1787 [0]}),
    .c({open_n7273,\u2_Display/n1785 }),
    .d({open_n7276,\u2_Display/n1784 }),
    .f({open_n7290,\u2_Display/n1819 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1612|_al_u1613  (
    .b({\u2_Display/n1787 [1],\u2_Display/n1787 [2]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1783 ,\u2_Display/n1782 }),
    .f({\u2_Display/n1818 ,\u2_Display/n1817 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1614|_al_u1615  (
    .b({\u2_Display/n1787 [3],\u2_Display/n1787 [4]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1781 ,\u2_Display/n1780 }),
    .f({\u2_Display/n1816 ,\u2_Display/n1815 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1616|_al_u1617  (
    .b({\u2_Display/n1787 [5],\u2_Display/n1787 [6]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1779 ,\u2_Display/n1778 }),
    .f({\u2_Display/n1814 ,\u2_Display/n1813 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1618|_al_u1621  (
    .b({\u2_Display/n1787 [7],\u2_Display/n1787 [10]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1777 ,\u2_Display/n1774 }),
    .f({\u2_Display/n1812 ,\u2_Display/n1809 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1619|_al_u1620  (
    .b({\u2_Display/n1787 [8],\u2_Display/n1787 [9]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1776 ,\u2_Display/n1775 }),
    .f({\u2_Display/n1811 ,\u2_Display/n1810 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1622|_al_u1625  (
    .b({\u2_Display/n1787 [11],\u2_Display/n1787 [14]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1773 ,\u2_Display/n1770 }),
    .f({\u2_Display/n1808 ,\u2_Display/n1805 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1623|_al_u1624  (
    .b({\u2_Display/n1787 [12],\u2_Display/n1787 [13]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1772 ,\u2_Display/n1771 }),
    .f({\u2_Display/n1807 ,\u2_Display/n1806 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1626|_al_u1629  (
    .b({\u2_Display/n1787 [15],\u2_Display/n1787 [18]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1769 ,\u2_Display/n1766 }),
    .f({\u2_Display/n1804 ,\u2_Display/n1801 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1627|_al_u1628  (
    .b({\u2_Display/n1787 [16],\u2_Display/n1787 [17]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1768 ,\u2_Display/n1767 }),
    .f({\u2_Display/n1803 ,\u2_Display/n1802 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1630|_al_u1631  (
    .b({\u2_Display/n1787 [19],\u2_Display/n1787 [20]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1765 ,\u2_Display/n1764 }),
    .f({\u2_Display/n1800 ,\u2_Display/n1799 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1632|_al_u1633  (
    .b({\u2_Display/n1787 [21],\u2_Display/n1787 [22]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1763 ,\u2_Display/n1762 }),
    .f({\u2_Display/n1798 ,\u2_Display/n1797 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1634|_al_u1637  (
    .b({\u2_Display/n1787 [23],\u2_Display/n1787 [26]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1761 ,\u2_Display/n1758 }),
    .f({\u2_Display/n1796 ,\u2_Display/n1793 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1636|_al_u1639  (
    .b({\u2_Display/n1787 [25],\u2_Display/n1787 [28]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1759 ,\u2_Display/n1756 }),
    .f({\u2_Display/n1794 ,\u2_Display/n1791 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1638|_al_u1641  (
    .b({\u2_Display/n1787 [27],\u2_Display/n1787 [30]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1757 ,\u2_Display/n1754 }),
    .f({\u2_Display/n1792 ,\u2_Display/n1789 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1640|_al_u1642  (
    .b({\u2_Display/n1787 [29],\u2_Display/n1787 [31]}),
    .c({\u2_Display/n1785 ,\u2_Display/n1785 }),
    .d({\u2_Display/n1755 ,\u2_Display/n1753 }),
    .f({\u2_Display/n1790 ,\u2_Display/n1788 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1643|_al_u1645  (
    .b({\u2_Display/n2910 [0],\u2_Display/n2910 [2]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2907 ,\u2_Display/n2905 }),
    .f({\u2_Display/n2942 ,\u2_Display/n2940 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1644|_al_u1648  (
    .b({\u2_Display/n2910 [1],\u2_Display/n2910 [5]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2906 ,\u2_Display/n2902 }),
    .f({\u2_Display/n2941 ,\u2_Display/n2937 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1646|_al_u1651  (
    .b({\u2_Display/n2910 [3],\u2_Display/n2910 [8]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2904 ,\u2_Display/n2899 }),
    .f({\u2_Display/n2939 ,\u2_Display/n2934 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1647|_al_u1649  (
    .b({\u2_Display/n2910 [4],\u2_Display/n2910 [6]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2903 ,\u2_Display/n2901 }),
    .f({\u2_Display/n2938 ,\u2_Display/n2936 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1650|_al_u1653  (
    .b({\u2_Display/n2910 [7],\u2_Display/n2910 [10]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2900 ,\u2_Display/n2897 }),
    .f({\u2_Display/n2935 ,\u2_Display/n2932 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1652|_al_u1655  (
    .b({\u2_Display/n2910 [9],\u2_Display/n2910 [12]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2898 ,\u2_Display/n2895 }),
    .f({\u2_Display/n2933 ,\u2_Display/n2930 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1654|_al_u1657  (
    .b({\u2_Display/n2910 [11],\u2_Display/n2910 [14]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2896 ,\u2_Display/n2893 }),
    .f({\u2_Display/n2931 ,\u2_Display/n2928 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1656|_al_u1659  (
    .b({\u2_Display/n2910 [13],\u2_Display/n2910 [16]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2894 ,\u2_Display/n2891 }),
    .f({\u2_Display/n2929 ,\u2_Display/n2926 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1658|_al_u1661  (
    .b({\u2_Display/n2910 [15],\u2_Display/n2910 [18]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2892 ,\u2_Display/n2889 }),
    .f({\u2_Display/n2927 ,\u2_Display/n2924 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1660|_al_u1664  (
    .b({\u2_Display/n2910 [17],\u2_Display/n2910 [21]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2890 ,\u2_Display/n2886 }),
    .f({\u2_Display/n2925 ,\u2_Display/n2921 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1662|_al_u1668  (
    .b({\u2_Display/n2910 [19],\u2_Display/n2910 [25]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2888 ,\u2_Display/n2882 }),
    .f({\u2_Display/n2923 ,\u2_Display/n2917 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1663|_al_u1665  (
    .b({\u2_Display/n2910 [20],\u2_Display/n2910 [22]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2887 ,\u2_Display/n2885 }),
    .f({\u2_Display/n2922 ,\u2_Display/n2920 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1666|_al_u1672  (
    .b({\u2_Display/n2910 [23],\u2_Display/n2910 [29]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2884 ,\u2_Display/n2878 }),
    .f({\u2_Display/n2919 ,\u2_Display/n2913 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1667|_al_u1669  (
    .b({\u2_Display/n2910 [24],\u2_Display/n2910 [26]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2883 ,\u2_Display/n2881 }),
    .f({\u2_Display/n2918 ,\u2_Display/n2916 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1670|_al_u1674  (
    .b({\u2_Display/n2910 [27],\u2_Display/n2910 [31]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2880 ,\u2_Display/n2876 }),
    .f({\u2_Display/n2915 ,\u2_Display/n2911 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1671|_al_u1673  (
    .b({\u2_Display/n2910 [28],\u2_Display/n2910 [30]}),
    .c({\u2_Display/n2908 ,\u2_Display/n2908 }),
    .d({\u2_Display/n2879 ,\u2_Display/n2877 }),
    .f({\u2_Display/n2914 ,\u2_Display/n2912 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u1675 (
    .b({open_n8044,\u2_Display/n4068 [0]}),
    .c({open_n8045,\u2_Display/n4066 }),
    .d({open_n8048,\u2_Display/n4065 }),
    .f({open_n8066,\u2_Display/n4100 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1676|_al_u1677  (
    .b({\u2_Display/n4068 [1],\u2_Display/n4068 [2]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4064 ,\u2_Display/n4063 }),
    .f({\u2_Display/n4099 ,\u2_Display/n4098 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1678|_al_u1681  (
    .b({\u2_Display/n4068 [3],\u2_Display/n4068 [6]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4062 ,\u2_Display/n4059 }),
    .f({\u2_Display/n4097 ,\u2_Display/n4094 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1679|_al_u1680  (
    .b({\u2_Display/n4068 [4],\u2_Display/n4068 [5]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4061 ,\u2_Display/n4060 }),
    .f({\u2_Display/n4096 ,\u2_Display/n4095 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1682|_al_u1683  (
    .b({\u2_Display/n4068 [7],\u2_Display/n4068 [8]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4058 ,\u2_Display/n4057 }),
    .f({\u2_Display/n4093 ,\u2_Display/n4092 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1684|_al_u1685  (
    .b({\u2_Display/n4068 [9],\u2_Display/n4068 [10]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4056 ,\u2_Display/n4055 }),
    .f({\u2_Display/n4091 ,\u2_Display/n4090 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1686|_al_u1687  (
    .b({\u2_Display/n4068 [11],\u2_Display/n4068 [12]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4054 ,\u2_Display/n4053 }),
    .f({\u2_Display/n4089 ,\u2_Display/n4088 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1688|_al_u1689  (
    .b({\u2_Display/n4068 [13],\u2_Display/n4068 [14]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4052 ,\u2_Display/n4051 }),
    .f({\u2_Display/n4087 ,\u2_Display/n4086 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1690|_al_u1691  (
    .b({\u2_Display/n4068 [15],\u2_Display/n4068 [16]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4050 ,\u2_Display/n4049 }),
    .f({\u2_Display/n4085 ,\u2_Display/n4084 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1692|_al_u1693  (
    .b({\u2_Display/n4068 [17],\u2_Display/n4068 [18]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4048 ,\u2_Display/n4047 }),
    .f({\u2_Display/n4083 ,\u2_Display/n4082 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1694|_al_u1695  (
    .b({\u2_Display/n4068 [19],\u2_Display/n4068 [20]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4046 ,\u2_Display/n4045 }),
    .f({\u2_Display/n4081 ,\u2_Display/n4080 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1696|_al_u1697  (
    .b({\u2_Display/n4068 [21],\u2_Display/n4068 [22]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4044 ,\u2_Display/n4043 }),
    .f({\u2_Display/n4079 ,\u2_Display/n4078 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1698|_al_u1701  (
    .b({\u2_Display/n4068 [23],\u2_Display/n4068 [26]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4042 ,\u2_Display/n4039 }),
    .f({\u2_Display/n4077 ,\u2_Display/n4074 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u1699 (
    .b({open_n8362,\u2_Display/n4068 [24]}),
    .c({open_n8363,\u2_Display/n4066 }),
    .d({open_n8366,\u2_Display/n4041 }),
    .f({open_n8384,\u2_Display/n4076 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1700|_al_u1704  (
    .b({\u2_Display/n4068 [25],\u2_Display/n4068 [29]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4040 ,\u2_Display/n4036 }),
    .f({\u2_Display/n4075 ,\u2_Display/n4071 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1702|_al_u1706  (
    .b({\u2_Display/n4068 [27],\u2_Display/n4068 [31]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4038 ,\u2_Display/n4034 }),
    .f({\u2_Display/n4073 ,\u2_Display/n4069 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1703|_al_u1705  (
    .b({\u2_Display/n4068 [28],\u2_Display/n4068 [30]}),
    .c({\u2_Display/n4066 ,\u2_Display/n4066 }),
    .d({\u2_Display/n4037 ,\u2_Display/n4035 }),
    .f({\u2_Display/n4072 ,\u2_Display/n4070 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1707|_al_u1709  (
    .b({\u2_Display/n5191 [0],\u2_Display/n5191 [2]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6346 ,\u2_Display/n6344 }),
    .f({\u2_Display/n5223 ,\u2_Display/n5221 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u1708 (
    .b({open_n8484,\u2_Display/n5191 [1]}),
    .c({open_n8485,\u2_Display/n5189 }),
    .d({open_n8488,\u2_Display/n6345 }),
    .f({open_n8506,\u2_Display/n5222 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1710|_al_u1713  (
    .b({\u2_Display/n5191 [3],\u2_Display/n5191 [6]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6343 ,\u2_Display/n6340 }),
    .f({\u2_Display/n5220 ,\u2_Display/n5217 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1711|_al_u1712  (
    .b({\u2_Display/n5191 [4],\u2_Display/n5191 [5]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6342 ,\u2_Display/n6341 }),
    .f({\u2_Display/n5219 ,\u2_Display/n5218 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1714|_al_u1717  (
    .b({\u2_Display/n5191 [7],\u2_Display/n5191 [10]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6339 ,\u2_Display/n6336 }),
    .f({\u2_Display/n5216 ,\u2_Display/n5213 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1715|_al_u1716  (
    .b({\u2_Display/n5191 [8],\u2_Display/n5191 [9]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6338 ,\u2_Display/n6337 }),
    .f({\u2_Display/n5215 ,\u2_Display/n5214 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1718|_al_u1721  (
    .b({\u2_Display/n5191 [11],\u2_Display/n5191 [14]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6335 ,\u2_Display/n6332 }),
    .f({\u2_Display/n5212 ,\u2_Display/n5209 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1719|_al_u1720  (
    .b({\u2_Display/n5191 [12],\u2_Display/n5191 [13]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6334 ,\u2_Display/n6333 }),
    .f({\u2_Display/n5211 ,\u2_Display/n5210 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1722|_al_u1723  (
    .b({\u2_Display/n5191 [15],\u2_Display/n5191 [16]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6331 ,\u2_Display/n6330 }),
    .f({\u2_Display/n5208 ,\u2_Display/n5207 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1724|_al_u1725  (
    .b({\u2_Display/n5191 [17],\u2_Display/n5191 [18]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6329 ,\u2_Display/n6328 }),
    .f({\u2_Display/n5206 ,\u2_Display/n5205 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1726|_al_u1727  (
    .b({\u2_Display/n5191 [19],\u2_Display/n5191 [20]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6327 ,\u2_Display/n6326 }),
    .f({\u2_Display/n5204 ,\u2_Display/n5203 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1728|_al_u1729  (
    .b({\u2_Display/n5191 [21],\u2_Display/n5191 [22]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6325 ,\u2_Display/n6324 }),
    .f({\u2_Display/n5202 ,\u2_Display/n5201 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1730|_al_u1735  (
    .b({\u2_Display/n5191 [23],\u2_Display/n5191 [28]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6323 ,\u2_Display/n6318 }),
    .f({\u2_Display/n5200 ,\u2_Display/n6353 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1731|_al_u1733  (
    .b({\u2_Display/n5191 [24],\u2_Display/n5191 [26]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6322 ,\u2_Display/n6320 }),
    .f({\u2_Display/n5199 ,\u2_Display/n5197 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u1732 (
    .b({open_n8798,\u2_Display/n5191 [25]}),
    .c({open_n8799,\u2_Display/n5189 }),
    .d({open_n8802,\u2_Display/n6321 }),
    .f({open_n8820,\u2_Display/n5198 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1734|_al_u1737  (
    .b({\u2_Display/n5191 [27],\u2_Display/n5191 [30]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6319 ,\u2_Display/n6316 }),
    .f({\u2_Display/n5196 ,\u2_Display/n6351 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1736|_al_u1738  (
    .b({\u2_Display/n5191 [29],\u2_Display/n5191 [31]}),
    .c({\u2_Display/n5189 ,\u2_Display/n5189 }),
    .d({\u2_Display/n6317 ,\u2_Display/n6315 }),
    .f({\u2_Display/n6352 ,\u2_Display/n6350 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1739|_al_u1741  (
    .b({\u2_Display/n699 [0],\u2_Display/n699 [2]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n696 ,\u2_Display/n694 }),
    .f({\u2_Display/n731 ,\u2_Display/n729 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1740|_al_u1743  (
    .b({\u2_Display/n699 [1],\u2_Display/n699 [4]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n695 ,\u2_Display/n692 }),
    .f({\u2_Display/n730 ,\u2_Display/n727 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1742|_al_u1745  (
    .b({\u2_Display/n699 [3],\u2_Display/n699 [6]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n693 ,\u2_Display/n690 }),
    .f({\u2_Display/n728 ,\u2_Display/n725 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1744|_al_u1747  (
    .b({\u2_Display/n699 [5],\u2_Display/n699 [8]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n691 ,\u2_Display/n688 }),
    .f({\u2_Display/n726 ,\u2_Display/n723 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1746|_al_u1749  (
    .b({\u2_Display/n699 [7],\u2_Display/n699 [10]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n689 ,\u2_Display/n686 }),
    .f({\u2_Display/n724 ,\u2_Display/n721 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1748|_al_u1752  (
    .b({\u2_Display/n699 [9],\u2_Display/n699 [13]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n687 ,\u2_Display/n683 }),
    .f({\u2_Display/n722 ,\u2_Display/n718 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1750|_al_u1756  (
    .b({\u2_Display/n699 [11],\u2_Display/n699 [17]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n685 ,\u2_Display/n679 }),
    .f({\u2_Display/n720 ,\u2_Display/n714 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1751|_al_u1753  (
    .b({\u2_Display/n699 [12],\u2_Display/n699 [14]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n684 ,\u2_Display/n682 }),
    .f({\u2_Display/n719 ,\u2_Display/n717 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1754|_al_u1760  (
    .b({\u2_Display/n699 [15],\u2_Display/n699 [21]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n681 ,\u2_Display/n675 }),
    .f({\u2_Display/n716 ,\u2_Display/n710 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1755|_al_u1757  (
    .b({\u2_Display/n699 [16],\u2_Display/n699 [18]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n680 ,\u2_Display/n678 }),
    .f({\u2_Display/n715 ,\u2_Display/n713 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1758|_al_u1763  (
    .b({\u2_Display/n699 [19],\u2_Display/n699 [24]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n677 ,\u2_Display/n672 }),
    .f({\u2_Display/n712 ,\u2_Display/n707 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1759|_al_u1761  (
    .b({\u2_Display/n699 [20],\u2_Display/n699 [22]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n676 ,\u2_Display/n674 }),
    .f({\u2_Display/n711 ,\u2_Display/n709 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1762|_al_u1765  (
    .b({\u2_Display/n699 [23],\u2_Display/n699 [26]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n673 ,\u2_Display/n670 }),
    .f({\u2_Display/n708 ,\u2_Display/n705 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1764|_al_u1767  (
    .b({\u2_Display/n699 [25],\u2_Display/n699 [28]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n671 ,\u2_Display/n668 }),
    .f({\u2_Display/n706 ,\u2_Display/n703 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1766|_al_u1769  (
    .b({\u2_Display/n699 [27],\u2_Display/n699 [30]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n669 ,\u2_Display/n666 }),
    .f({\u2_Display/n704 ,\u2_Display/n701 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1768|_al_u1770  (
    .b({\u2_Display/n699 [29],\u2_Display/n699 [31]}),
    .c({\u2_Display/n697 ,\u2_Display/n697 }),
    .d({\u2_Display/n667 ,\u2_Display/n665 }),
    .f({\u2_Display/n702 ,\u2_Display/n700 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1771|_al_u1775  (
    .b({\u2_Display/n1822 [0],\u2_Display/n1822 [4]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1819 ,\u2_Display/n1815 }),
    .f({\u2_Display/n1854 ,\u2_Display/n1850 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u1772|_al_u1773  (
    .b({\u2_Display/n1818 ,\u2_Display/n1822 [2]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1822 [1],\u2_Display/n1817 }),
    .f({\u2_Display/n1853 ,\u2_Display/n1852 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1774|_al_u1777  (
    .b({\u2_Display/n1822 [3],\u2_Display/n1822 [6]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1816 ,\u2_Display/n1813 }),
    .f({\u2_Display/n1851 ,\u2_Display/n1848 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1776|_al_u1780  (
    .b({\u2_Display/n1822 [5],\u2_Display/n1822 [9]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1814 ,\u2_Display/n1810 }),
    .f({\u2_Display/n1849 ,\u2_Display/n1845 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1778|_al_u1784  (
    .b({\u2_Display/n1822 [7],\u2_Display/n1822 [13]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1812 ,\u2_Display/n1806 }),
    .f({\u2_Display/n1847 ,\u2_Display/n1841 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1779|_al_u1781  (
    .b({\u2_Display/n1822 [8],\u2_Display/n1822 [10]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1811 ,\u2_Display/n1809 }),
    .f({\u2_Display/n1846 ,\u2_Display/n1844 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1782|_al_u1787  (
    .b({\u2_Display/n1822 [11],\u2_Display/n1822 [16]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1808 ,\u2_Display/n1803 }),
    .f({\u2_Display/n1843 ,\u2_Display/n1838 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1783|_al_u1785  (
    .b({\u2_Display/n1822 [12],\u2_Display/n1822 [14]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1807 ,\u2_Display/n1805 }),
    .f({\u2_Display/n1842 ,\u2_Display/n1840 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1786|_al_u1791  (
    .b({\u2_Display/n1822 [15],\u2_Display/n1822 [20]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1804 ,\u2_Display/n1799 }),
    .f({\u2_Display/n1839 ,\u2_Display/n1834 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1788|_al_u1789  (
    .b({\u2_Display/n1822 [17],\u2_Display/n1822 [18]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1802 ,\u2_Display/n1801 }),
    .f({\u2_Display/n1837 ,\u2_Display/n1836 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1790|_al_u1793  (
    .b({\u2_Display/n1822 [19],\u2_Display/n1822 [22]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1800 ,\u2_Display/n1797 }),
    .f({\u2_Display/n1835 ,\u2_Display/n1832 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1792|_al_u1795  (
    .b({\u2_Display/n1822 [21],\u2_Display/n1822 [24]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1798 ,\u2_Display/n1795 }),
    .f({\u2_Display/n1833 ,\u2_Display/n1830 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1794|_al_u1797  (
    .b({\u2_Display/n1822 [23],\u2_Display/n1822 [26]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1796 ,\u2_Display/n1793 }),
    .f({\u2_Display/n1831 ,\u2_Display/n1828 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1796|_al_u1799  (
    .b({\u2_Display/n1822 [25],\u2_Display/n1822 [28]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1794 ,\u2_Display/n1791 }),
    .f({\u2_Display/n1829 ,\u2_Display/n1826 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1798|_al_u1801  (
    .b({\u2_Display/n1822 [27],\u2_Display/n1822 [30]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1792 ,\u2_Display/n1789 }),
    .f({\u2_Display/n1827 ,\u2_Display/n1824 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1800|_al_u1802  (
    .b({\u2_Display/n1822 [29],\u2_Display/n1822 [31]}),
    .c({\u2_Display/n1820 ,\u2_Display/n1820 }),
    .d({\u2_Display/n1790 ,\u2_Display/n1788 }),
    .f({\u2_Display/n1825 ,\u2_Display/n1823 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .MODE("LOGIC"))
    _al_u1803 (
    .b({open_n9648,\u2_Display/n2945 [0]}),
    .c({open_n9649,\u2_Display/n2943 }),
    .d({open_n9652,\u2_Display/n2942 }),
    .f({open_n9666,\u2_Display/n2977 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1804|_al_u1805  (
    .b({\u2_Display/n2945 [1],\u2_Display/n2945 [2]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2941 ,\u2_Display/n2940 }),
    .f({\u2_Display/n2976 ,\u2_Display/n2975 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1806|_al_u1994  (
    .b({\u2_Display/n2945 [3],\u2_Display/n2980 [31]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2939 ,\u2_Display/n2946 }),
    .f({\u2_Display/n2974 ,\u2_Display/n2981 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1807|_al_u1809  (
    .b({\u2_Display/n2945 [4],\u2_Display/n2945 [6]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2938 ,\u2_Display/n2936 }),
    .f({\u2_Display/n2973 ,\u2_Display/n2971 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1808|_al_u1812  (
    .b({\u2_Display/n2945 [5],\u2_Display/n2945 [9]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2937 ,\u2_Display/n2933 }),
    .f({\u2_Display/n2972 ,\u2_Display/n2968 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1810|_al_u1816  (
    .b({\u2_Display/n2945 [7],\u2_Display/n2945 [13]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2935 ,\u2_Display/n2929 }),
    .f({\u2_Display/n2970 ,\u2_Display/n2964 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1811|_al_u1813  (
    .b({\u2_Display/n2945 [8],\u2_Display/n2945 [10]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2934 ,\u2_Display/n2932 }),
    .f({\u2_Display/n2969 ,\u2_Display/n2967 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1814|_al_u1819  (
    .b({\u2_Display/n2945 [11],\u2_Display/n2945 [16]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2931 ,\u2_Display/n2926 }),
    .f({\u2_Display/n2966 ,\u2_Display/n2961 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1815|_al_u1817  (
    .b({\u2_Display/n2945 [12],\u2_Display/n2945 [14]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2930 ,\u2_Display/n2928 }),
    .f({\u2_Display/n2965 ,\u2_Display/n2963 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1818|_al_u1821  (
    .b({\u2_Display/n2945 [15],\u2_Display/n2945 [18]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2927 ,\u2_Display/n2924 }),
    .f({\u2_Display/n2962 ,\u2_Display/n2959 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1820|_al_u1823  (
    .b({\u2_Display/n2945 [17],\u2_Display/n2945 [20]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2925 ,\u2_Display/n2922 }),
    .f({\u2_Display/n2960 ,\u2_Display/n2957 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1822|_al_u1825  (
    .b({\u2_Display/n2945 [19],\u2_Display/n2945 [22]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2923 ,\u2_Display/n2920 }),
    .f({\u2_Display/n2958 ,\u2_Display/n2955 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1824|_al_u1828  (
    .b({\u2_Display/n2945 [21],\u2_Display/n2945 [25]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2921 ,\u2_Display/n2917 }),
    .f({\u2_Display/n2956 ,\u2_Display/n2952 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1826|_al_u1831  (
    .b({\u2_Display/n2945 [23],\u2_Display/n2945 [28]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2919 ,\u2_Display/n2914 }),
    .f({\u2_Display/n2954 ,\u2_Display/n2949 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1827|_al_u1829  (
    .b({\u2_Display/n2945 [24],\u2_Display/n2945 [26]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2918 ,\u2_Display/n2916 }),
    .f({\u2_Display/n2953 ,\u2_Display/n2951 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1830|_al_u1833  (
    .b({\u2_Display/n2945 [27],\u2_Display/n2945 [30]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2915 ,\u2_Display/n2912 }),
    .f({\u2_Display/n2950 ,\u2_Display/n2947 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1832|_al_u1834  (
    .b({\u2_Display/n2945 [29],\u2_Display/n2945 [31]}),
    .c({\u2_Display/n2943 ,\u2_Display/n2943 }),
    .d({\u2_Display/n2913 ,\u2_Display/n2911 }),
    .f({\u2_Display/n2948 ,\u2_Display/n2946 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1835|_al_u1837  (
    .b({\u2_Display/n4103 [0],\u2_Display/n4103 [2]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4100 ,\u2_Display/n4098 }),
    .f({\u2_Display/n4135 ,\u2_Display/n4133 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u1836|_al_u1839  (
    .b({\u2_Display/n4101 ,\u2_Display/n4103 [4]}),
    .c({\u2_Display/n4103 [1],\u2_Display/n4101 }),
    .d({\u2_Display/n4099 ,\u2_Display/n4096 }),
    .f({\u2_Display/n4134 ,\u2_Display/n4131 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1838|_al_u1841  (
    .b({\u2_Display/n4103 [3],\u2_Display/n4103 [6]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4097 ,\u2_Display/n4094 }),
    .f({\u2_Display/n4132 ,\u2_Display/n4129 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1840|_al_u1843  (
    .b({\u2_Display/n4103 [5],\u2_Display/n4103 [8]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4095 ,\u2_Display/n4092 }),
    .f({\u2_Display/n4130 ,\u2_Display/n4127 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1842|_al_u1845  (
    .b({\u2_Display/n4103 [7],\u2_Display/n4103 [10]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4093 ,\u2_Display/n4090 }),
    .f({\u2_Display/n4128 ,\u2_Display/n4125 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u1844|_al_u1847  (
    .b({\u2_Display/n4091 ,\u2_Display/n4103 [12]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4103 [9],\u2_Display/n4088 }),
    .f({\u2_Display/n4126 ,\u2_Display/n4123 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1846|_al_u1848  (
    .b({\u2_Display/n4103 [11],\u2_Display/n4103 [13]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4089 ,\u2_Display/n4087 }),
    .f({\u2_Display/n4124 ,\u2_Display/n4122 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1849|_al_u1851  (
    .b({\u2_Display/n4103 [14],\u2_Display/n4103 [16]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4086 ,\u2_Display/n4084 }),
    .f({\u2_Display/n4121 ,\u2_Display/n4119 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1850|_al_u1853  (
    .b({\u2_Display/n4103 [15],\u2_Display/n4103 [18]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4085 ,\u2_Display/n4082 }),
    .f({\u2_Display/n4120 ,\u2_Display/n4117 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1852|_al_u1855  (
    .b({\u2_Display/n4103 [17],\u2_Display/n4103 [20]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4083 ,\u2_Display/n4080 }),
    .f({\u2_Display/n4118 ,\u2_Display/n4115 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1854|_al_u1857  (
    .b({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .c({\u2_Display/n4103 [19],\u2_Display/n4103 [22]}),
    .d({\u2_Display/n4081 ,\u2_Display/n4078 }),
    .f({\u2_Display/n4116 ,\u2_Display/n4113 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1856|_al_u1860  (
    .b({\u2_Display/n4103 [21],\u2_Display/n4103 [25]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4079 ,\u2_Display/n4075 }),
    .f({\u2_Display/n4114 ,\u2_Display/n4110 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1858|_al_u1864  (
    .b({\u2_Display/n4103 [23],\u2_Display/n4103 [29]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4077 ,\u2_Display/n4071 }),
    .f({\u2_Display/n4112 ,\u2_Display/n4106 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1859|_al_u1861  (
    .b({\u2_Display/n4103 [24],\u2_Display/n4103 [26]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4076 ,\u2_Display/n4074 }),
    .f({\u2_Display/n4111 ,\u2_Display/n4109 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1862|_al_u1866  (
    .b({\u2_Display/n4103 [27],\u2_Display/n4103 [31]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4073 ,\u2_Display/n4069 }),
    .f({\u2_Display/n4108 ,\u2_Display/n4104 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1863|_al_u1865  (
    .b({\u2_Display/n4103 [28],\u2_Display/n4103 [30]}),
    .c({\u2_Display/n4101 ,\u2_Display/n4101 }),
    .d({\u2_Display/n4072 ,\u2_Display/n4070 }),
    .f({\u2_Display/n4107 ,\u2_Display/n4105 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1867|_al_u1871  (
    .b({\u2_Display/n5226 [0],\u2_Display/n5226 [4]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5223 ,\u2_Display/n5219 }),
    .f({\u2_Display/n5258 ,\u2_Display/n5254 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u1868|_al_u1869  (
    .b({\u2_Display/n5224 ,\u2_Display/n5226 [2]}),
    .c({\u2_Display/n5226 [1],\u2_Display/n5224 }),
    .d({\u2_Display/n5222 ,\u2_Display/n5221 }),
    .f({\u2_Display/n5257 ,\u2_Display/n5256 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1870|_al_u1873  (
    .b({\u2_Display/n5226 [3],\u2_Display/n5226 [6]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5220 ,\u2_Display/n5217 }),
    .f({\u2_Display/n5255 ,\u2_Display/n5252 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1872|_al_u1875  (
    .b({\u2_Display/n5226 [5],\u2_Display/n5226 [8]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5218 ,\u2_Display/n5215 }),
    .f({\u2_Display/n5253 ,\u2_Display/n5250 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1874|_al_u1877  (
    .b({\u2_Display/n5226 [7],\u2_Display/n5226 [10]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5216 ,\u2_Display/n5213 }),
    .f({\u2_Display/n5251 ,\u2_Display/n5248 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u1876|_al_u1880  (
    .b({\u2_Display/n5214 ,\u2_Display/n5226 [13]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5226 [9],\u2_Display/n5210 }),
    .f({\u2_Display/n5249 ,\u2_Display/n5245 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1878|_al_u1883  (
    .b({\u2_Display/n5226 [11],\u2_Display/n5226 [16]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5212 ,\u2_Display/n5207 }),
    .f({\u2_Display/n5247 ,\u2_Display/n5242 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1879|_al_u1881  (
    .b({\u2_Display/n5226 [12],\u2_Display/n5226 [14]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5211 ,\u2_Display/n5209 }),
    .f({\u2_Display/n5246 ,\u2_Display/n5244 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1882|_al_u1885  (
    .b({\u2_Display/n5226 [15],\u2_Display/n5226 [18]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5208 ,\u2_Display/n5205 }),
    .f({\u2_Display/n5243 ,\u2_Display/n5240 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u1884|_al_u1887  (
    .b({\u2_Display/n5206 ,\u2_Display/n5226 [20]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5226 [17],\u2_Display/n5203 }),
    .f({\u2_Display/n5241 ,\u2_Display/n5238 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1886|_al_u1889  (
    .b({\u2_Display/n5226 [19],\u2_Display/n5226 [22]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5204 ,\u2_Display/n5201 }),
    .f({\u2_Display/n5239 ,\u2_Display/n5236 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1888|_al_u1891  (
    .b({\u2_Display/n5226 [21],\u2_Display/n5226 [24]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5202 ,\u2_Display/n5199 }),
    .f({\u2_Display/n5237 ,\u2_Display/n5234 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1890|_al_u1893  (
    .b({\u2_Display/n5226 [23],\u2_Display/n5226 [26]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5200 ,\u2_Display/n5197 }),
    .f({\u2_Display/n5235 ,\u2_Display/n5232 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1892|_al_u1895  (
    .b({\u2_Display/n5226 [25],\u2_Display/n5226 [28]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5198 ,\u2_Display/n6353 }),
    .f({\u2_Display/n5233 ,\u2_Display/n5230 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1894|_al_u1897  (
    .b({\u2_Display/n5226 [27],\u2_Display/n5226 [30]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n5196 ,\u2_Display/n6351 }),
    .f({\u2_Display/n5231 ,\u2_Display/n5228 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1896|_al_u1898  (
    .b({\u2_Display/n5226 [29],\u2_Display/n5226 [31]}),
    .c({\u2_Display/n5224 ,\u2_Display/n5224 }),
    .d({\u2_Display/n6352 ,\u2_Display/n6350 }),
    .f({\u2_Display/n5229 ,\u2_Display/n5227 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1899|_al_u1901  (
    .b({\u2_Display/n734 [0],\u2_Display/n734 [2]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n731 ,\u2_Display/n729 }),
    .f({\u2_Display/n766 ,\u2_Display/n764 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .MODE("LOGIC"))
    _al_u1900 (
    .b({open_n10848,\u2_Display/n734 [1]}),
    .c({open_n10849,\u2_Display/n732 }),
    .d({open_n10852,\u2_Display/n730 }),
    .f({open_n10866,\u2_Display/n765 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1902|_al_u1905  (
    .b({\u2_Display/n734 [3],\u2_Display/n734 [6]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n728 ,\u2_Display/n725 }),
    .f({\u2_Display/n763 ,\u2_Display/n760 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1903|_al_u1904  (
    .b({\u2_Display/n734 [4],\u2_Display/n734 [5]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n727 ,\u2_Display/n726 }),
    .f({\u2_Display/n762 ,\u2_Display/n761 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1906|_al_u1909  (
    .b({\u2_Display/n734 [7],\u2_Display/n734 [10]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n724 ,\u2_Display/n721 }),
    .f({\u2_Display/n759 ,\u2_Display/n756 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1907|_al_u1908  (
    .b({\u2_Display/n734 [8],\u2_Display/n734 [9]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n723 ,\u2_Display/n722 }),
    .f({\u2_Display/n758 ,\u2_Display/n757 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1910|_al_u1913  (
    .b({\u2_Display/n734 [11],\u2_Display/n734 [14]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n720 ,\u2_Display/n717 }),
    .f({\u2_Display/n755 ,\u2_Display/n752 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1911|_al_u1912  (
    .b({\u2_Display/n734 [12],\u2_Display/n734 [13]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n719 ,\u2_Display/n718 }),
    .f({\u2_Display/n754 ,\u2_Display/n753 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1914|_al_u1915  (
    .b({\u2_Display/n734 [15],\u2_Display/n734 [16]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n716 ,\u2_Display/n715 }),
    .f({\u2_Display/n751 ,\u2_Display/n750 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1916|_al_u1917  (
    .b({\u2_Display/n734 [17],\u2_Display/n734 [18]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n714 ,\u2_Display/n713 }),
    .f({\u2_Display/n749 ,\u2_Display/n748 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1918|_al_u1919  (
    .b({\u2_Display/n734 [19],\u2_Display/n734 [20]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n712 ,\u2_Display/n711 }),
    .f({\u2_Display/n747 ,\u2_Display/n746 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1920|_al_u1921  (
    .b({\u2_Display/n734 [21],\u2_Display/n734 [22]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n710 ,\u2_Display/n709 }),
    .f({\u2_Display/n745 ,\u2_Display/n744 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1922|_al_u1925  (
    .b({\u2_Display/n734 [23],\u2_Display/n734 [26]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n708 ,\u2_Display/n705 }),
    .f({\u2_Display/n743 ,\u2_Display/n740 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .MODE("LOGIC"))
    _al_u1923 (
    .b({open_n11140,\u2_Display/n734 [24]}),
    .c({open_n11141,\u2_Display/n732 }),
    .d({open_n11144,\u2_Display/n707 }),
    .f({open_n11158,\u2_Display/n742 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1924|_al_u1927  (
    .b({\u2_Display/n734 [25],\u2_Display/n734 [28]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n706 ,\u2_Display/n703 }),
    .f({\u2_Display/n741 ,\u2_Display/n738 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1926|_al_u1929  (
    .b({\u2_Display/n734 [27],\u2_Display/n734 [30]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n704 ,\u2_Display/n701 }),
    .f({\u2_Display/n739 ,\u2_Display/n736 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1928|_al_u1930  (
    .b({\u2_Display/n734 [29],\u2_Display/n734 [31]}),
    .c({\u2_Display/n732 ,\u2_Display/n732 }),
    .d({\u2_Display/n702 ,\u2_Display/n700 }),
    .f({\u2_Display/n737 ,\u2_Display/n735 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1931|_al_u1935  (
    .b({\u2_Display/n1857 [0],\u2_Display/n1857 [4]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1854 ,\u2_Display/n1850 }),
    .f({\u2_Display/n1889 ,\u2_Display/n1885 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1932|_al_u1933  (
    .b({\u2_Display/n1857 [1],\u2_Display/n1857 [2]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1853 ,\u2_Display/n1852 }),
    .f({\u2_Display/n1888 ,\u2_Display/n1887 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1934|_al_u1937  (
    .b({\u2_Display/n1857 [3],\u2_Display/n1857 [6]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1851 ,\u2_Display/n1848 }),
    .f({\u2_Display/n1886 ,\u2_Display/n1883 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1936|_al_u1940  (
    .b({\u2_Display/n1857 [5],\u2_Display/n1857 [9]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1849 ,\u2_Display/n1845 }),
    .f({\u2_Display/n1884 ,\u2_Display/n1880 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1938|_al_u1943  (
    .b({\u2_Display/n1857 [7],\u2_Display/n1857 [12]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1847 ,\u2_Display/n1842 }),
    .f({\u2_Display/n1882 ,\u2_Display/n1877 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1939|_al_u1941  (
    .b({\u2_Display/n1857 [8],\u2_Display/n1857 [10]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1846 ,\u2_Display/n1844 }),
    .f({\u2_Display/n1881 ,\u2_Display/n1879 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1942|_al_u1945  (
    .b({\u2_Display/n1857 [11],\u2_Display/n1857 [14]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1843 ,\u2_Display/n1840 }),
    .f({\u2_Display/n1878 ,\u2_Display/n1875 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1944|_al_u1947  (
    .b({\u2_Display/n1857 [13],\u2_Display/n1857 [16]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1841 ,\u2_Display/n1838 }),
    .f({\u2_Display/n1876 ,\u2_Display/n1873 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1946|_al_u1949  (
    .b({\u2_Display/n1857 [15],\u2_Display/n1857 [18]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1839 ,\u2_Display/n1836 }),
    .f({\u2_Display/n1874 ,\u2_Display/n1871 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1948|_al_u1952  (
    .b({\u2_Display/n1857 [17],\u2_Display/n1857 [21]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1837 ,\u2_Display/n1833 }),
    .f({\u2_Display/n1872 ,\u2_Display/n1868 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1950|_al_u1955  (
    .b({\u2_Display/n1857 [19],\u2_Display/n1857 [24]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1835 ,\u2_Display/n1830 }),
    .f({\u2_Display/n1870 ,\u2_Display/n1865 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1951|_al_u1953  (
    .b({\u2_Display/n1857 [20],\u2_Display/n1857 [22]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1834 ,\u2_Display/n1832 }),
    .f({\u2_Display/n1869 ,\u2_Display/n1867 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1954|_al_u1957  (
    .b({\u2_Display/n1857 [23],\u2_Display/n1857 [26]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1831 ,\u2_Display/n1828 }),
    .f({\u2_Display/n1866 ,\u2_Display/n1863 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1956|_al_u1960  (
    .b({\u2_Display/n1857 [25],\u2_Display/n1857 [29]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1829 ,\u2_Display/n1825 }),
    .f({\u2_Display/n1864 ,\u2_Display/n1860 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1958|_al_u1962  (
    .b({\u2_Display/n1857 [27],\u2_Display/n1857 [31]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1827 ,\u2_Display/n1823 }),
    .f({\u2_Display/n1862 ,\u2_Display/n1858 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1959|_al_u1961  (
    .b({\u2_Display/n1857 [28],\u2_Display/n1857 [30]}),
    .c({\u2_Display/n1855 ,\u2_Display/n1855 }),
    .d({\u2_Display/n1826 ,\u2_Display/n1824 }),
    .f({\u2_Display/n1861 ,\u2_Display/n1859 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1963|_al_u1965  (
    .b({\u2_Display/n2980 [0],\u2_Display/n2980 [2]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2977 ,\u2_Display/n2975 }),
    .f({\u2_Display/n3012 ,\u2_Display/n3010 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .MODE("LOGIC"))
    _al_u1964 (
    .b({open_n11650,\u2_Display/n2980 [1]}),
    .c({open_n11651,\u2_Display/n2978 }),
    .d({open_n11654,\u2_Display/n2976 }),
    .f({open_n11668,\u2_Display/n3011 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1966|_al_u1967  (
    .b({\u2_Display/n2980 [3],\u2_Display/n2980 [4]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2974 ,\u2_Display/n2973 }),
    .f({\u2_Display/n3009 ,\u2_Display/n3008 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1968|_al_u1969  (
    .b({\u2_Display/n2980 [5],\u2_Display/n2980 [6]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2972 ,\u2_Display/n2971 }),
    .f({\u2_Display/n3007 ,\u2_Display/n3006 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1970|_al_u1971  (
    .b({\u2_Display/n2980 [7],\u2_Display/n2980 [8]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2970 ,\u2_Display/n2969 }),
    .f({\u2_Display/n3005 ,\u2_Display/n3004 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1972|_al_u1973  (
    .b({\u2_Display/n2980 [9],\u2_Display/n2980 [10]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2968 ,\u2_Display/n2967 }),
    .f({\u2_Display/n3003 ,\u2_Display/n3002 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1974|_al_u1975  (
    .b({\u2_Display/n2980 [11],\u2_Display/n2980 [12]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2966 ,\u2_Display/n2965 }),
    .f({\u2_Display/n3001 ,\u2_Display/n3000 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1976|_al_u1977  (
    .b({\u2_Display/n2980 [13],\u2_Display/n2980 [14]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2964 ,\u2_Display/n2963 }),
    .f({\u2_Display/n2999 ,\u2_Display/n2998 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1978|_al_u1979  (
    .b({\u2_Display/n2980 [15],\u2_Display/n2980 [16]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2962 ,\u2_Display/n2961 }),
    .f({\u2_Display/n2997 ,\u2_Display/n2996 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1980|_al_u1981  (
    .b({\u2_Display/n2980 [17],\u2_Display/n2980 [18]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2960 ,\u2_Display/n2959 }),
    .f({\u2_Display/n2995 ,\u2_Display/n2994 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1982|_al_u1985  (
    .b({\u2_Display/n2980 [19],\u2_Display/n2980 [22]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2958 ,\u2_Display/n2955 }),
    .f({\u2_Display/n2993 ,\u2_Display/n2990 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1983|_al_u1984  (
    .b({\u2_Display/n2980 [20],\u2_Display/n2980 [21]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2957 ,\u2_Display/n2956 }),
    .f({\u2_Display/n2992 ,\u2_Display/n2991 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1986|_al_u1987  (
    .b({\u2_Display/n2980 [23],\u2_Display/n2980 [24]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2954 ,\u2_Display/n2953 }),
    .f({\u2_Display/n2989 ,\u2_Display/n2988 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1988|_al_u1989  (
    .b({\u2_Display/n2980 [25],\u2_Display/n2980 [26]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2952 ,\u2_Display/n2951 }),
    .f({\u2_Display/n2987 ,\u2_Display/n2986 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1990|_al_u1993  (
    .b({\u2_Display/n2980 [27],\u2_Display/n2980 [30]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2950 ,\u2_Display/n2947 }),
    .f({\u2_Display/n2985 ,\u2_Display/n2982 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1991|_al_u1992  (
    .b({\u2_Display/n2980 [28],\u2_Display/n2980 [29]}),
    .c({\u2_Display/n2978 ,\u2_Display/n2978 }),
    .d({\u2_Display/n2949 ,\u2_Display/n2948 }),
    .f({\u2_Display/n2984 ,\u2_Display/n2983 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1995|_al_u1997  (
    .b({\u2_Display/n4138 [0],\u2_Display/n4138 [2]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4135 ,\u2_Display/n4133 }),
    .f({\u2_Display/n4170 ,\u2_Display/n4168 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1996|_al_u1999  (
    .b({\u2_Display/n4138 [1],\u2_Display/n4138 [4]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4134 ,\u2_Display/n4131 }),
    .f({\u2_Display/n4169 ,\u2_Display/n4166 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u1998|_al_u2001  (
    .b({\u2_Display/n4138 [3],\u2_Display/n4138 [6]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4132 ,\u2_Display/n4129 }),
    .f({\u2_Display/n4167 ,\u2_Display/n4164 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2000|_al_u2003  (
    .b({\u2_Display/n4138 [5],\u2_Display/n4138 [8]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4130 ,\u2_Display/n4127 }),
    .f({\u2_Display/n4165 ,\u2_Display/n4162 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2002|_al_u2005  (
    .b({\u2_Display/n4138 [7],\u2_Display/n4138 [10]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4128 ,\u2_Display/n4125 }),
    .f({\u2_Display/n4163 ,\u2_Display/n4160 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2004|_al_u2007  (
    .b({\u2_Display/n4138 [9],\u2_Display/n4138 [12]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4126 ,\u2_Display/n4123 }),
    .f({\u2_Display/n4161 ,\u2_Display/n4158 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2006|_al_u2009  (
    .b({\u2_Display/n4138 [11],\u2_Display/n4138 [14]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4124 ,\u2_Display/n4121 }),
    .f({\u2_Display/n4159 ,\u2_Display/n4156 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2008|_al_u2012  (
    .b({\u2_Display/n4138 [13],\u2_Display/n4138 [17]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4122 ,\u2_Display/n4118 }),
    .f({\u2_Display/n4157 ,\u2_Display/n4153 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2010|_al_u2015  (
    .b({\u2_Display/n4138 [15],\u2_Display/n4138 [20]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4120 ,\u2_Display/n4115 }),
    .f({\u2_Display/n4155 ,\u2_Display/n4150 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2011|_al_u2013  (
    .b({\u2_Display/n4138 [16],\u2_Display/n4138 [18]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4119 ,\u2_Display/n4117 }),
    .f({\u2_Display/n4154 ,\u2_Display/n4152 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2014|_al_u2017  (
    .b({\u2_Display/n4138 [19],\u2_Display/n4138 [22]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4116 ,\u2_Display/n4113 }),
    .f({\u2_Display/n4151 ,\u2_Display/n4148 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2016|_al_u2019  (
    .b({\u2_Display/n4138 [21],\u2_Display/n4138 [24]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4114 ,\u2_Display/n4111 }),
    .f({\u2_Display/n4149 ,\u2_Display/n4146 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2018|_al_u2021  (
    .b({\u2_Display/n4138 [23],\u2_Display/n4138 [26]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4112 ,\u2_Display/n4109 }),
    .f({\u2_Display/n4147 ,\u2_Display/n4144 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2020|_al_u2024  (
    .b({\u2_Display/n4138 [25],\u2_Display/n4138 [29]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4110 ,\u2_Display/n4106 }),
    .f({\u2_Display/n4145 ,\u2_Display/n4141 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2022|_al_u2026  (
    .b({\u2_Display/n4138 [27],\u2_Display/n4138 [31]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4108 ,\u2_Display/n4104 }),
    .f({\u2_Display/n4143 ,\u2_Display/n4139 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2023|_al_u2025  (
    .b({\u2_Display/n4138 [28],\u2_Display/n4138 [30]}),
    .c({\u2_Display/n4136 ,\u2_Display/n4136 }),
    .d({\u2_Display/n4107 ,\u2_Display/n4105 }),
    .f({\u2_Display/n4142 ,\u2_Display/n4140 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2027|_al_u2029  (
    .b({\u2_Display/n5261 [0],\u2_Display/n5261 [2]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5258 ,\u2_Display/n5256 }),
    .f({\u2_Display/n5293 ,\u2_Display/n5291 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u2028 (
    .b({open_n12422,\u2_Display/n5261 [1]}),
    .c({open_n12423,\u2_Display/n5259 }),
    .d({open_n12426,\u2_Display/n5257 }),
    .f({open_n12444,\u2_Display/n5292 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2030|_al_u2033  (
    .b({\u2_Display/n5261 [3],\u2_Display/n5261 [6]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5255 ,\u2_Display/n5252 }),
    .f({\u2_Display/n5290 ,\u2_Display/n5287 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2031|_al_u2032  (
    .b({\u2_Display/n5261 [4],\u2_Display/n5261 [5]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5254 ,\u2_Display/n5253 }),
    .f({\u2_Display/n5289 ,\u2_Display/n5288 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2034|_al_u2035  (
    .b({\u2_Display/n5261 [7],\u2_Display/n5261 [8]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5251 ,\u2_Display/n5250 }),
    .f({\u2_Display/n5286 ,\u2_Display/n5285 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2036|_al_u2037  (
    .b({\u2_Display/n5261 [9],\u2_Display/n5261 [10]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5249 ,\u2_Display/n5248 }),
    .f({\u2_Display/n5284 ,\u2_Display/n5283 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2038|_al_u2039  (
    .b({\u2_Display/n5261 [11],\u2_Display/n5261 [12]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5247 ,\u2_Display/n5246 }),
    .f({\u2_Display/n5282 ,\u2_Display/n5281 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2040|_al_u2041  (
    .b({\u2_Display/n5261 [13],\u2_Display/n5261 [14]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5245 ,\u2_Display/n5244 }),
    .f({\u2_Display/n5280 ,\u2_Display/n5279 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2042|_al_u2045  (
    .b({\u2_Display/n5261 [15],\u2_Display/n5261 [18]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5243 ,\u2_Display/n5240 }),
    .f({\u2_Display/n5278 ,\u2_Display/n5275 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2043|_al_u2044  (
    .b({\u2_Display/n5261 [16],\u2_Display/n5261 [17]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5242 ,\u2_Display/n5241 }),
    .f({\u2_Display/n5277 ,\u2_Display/n5276 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2046|_al_u2047  (
    .b({\u2_Display/n5261 [19],\u2_Display/n5261 [20]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5239 ,\u2_Display/n5238 }),
    .f({\u2_Display/n5274 ,\u2_Display/n5273 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2048|_al_u2049  (
    .b({\u2_Display/n5261 [21],\u2_Display/n5261 [22]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5237 ,\u2_Display/n5236 }),
    .f({\u2_Display/n5272 ,\u2_Display/n5271 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2050|_al_u2053  (
    .b({\u2_Display/n5261 [23],\u2_Display/n5261 [26]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5235 ,\u2_Display/n5232 }),
    .f({\u2_Display/n5270 ,\u2_Display/n5267 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2051|_al_u2052  (
    .b({\u2_Display/n5261 [24],\u2_Display/n5261 [25]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5234 ,\u2_Display/n5233 }),
    .f({\u2_Display/n5269 ,\u2_Display/n5268 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2054|_al_u2057  (
    .b({\u2_Display/n5261 [27],\u2_Display/n5261 [30]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5231 ,\u2_Display/n5228 }),
    .f({\u2_Display/n5266 ,\u2_Display/n5263 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2055|_al_u2056  (
    .b({\u2_Display/n5261 [28],\u2_Display/n5261 [29]}),
    .c({\u2_Display/n5259 ,\u2_Display/n5259 }),
    .d({\u2_Display/n5230 ,\u2_Display/n5229 }),
    .f({\u2_Display/n5265 ,\u2_Display/n5264 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(~D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000000011111111),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0000000011111111),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2058|_al_u3999  (
    .b({\u2_Display/n5261 [31],open_n12784}),
    .c({\u2_Display/n5259 ,open_n12785}),
    .d({\u2_Display/n5227 ,rst_n_pad}),
    .f({\u2_Display/n5262 ,\u0_PLL/n0 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u2059 (
    .b({open_n12812,\u2_Display/n769 [0]}),
    .c({open_n12813,\u2_Display/n767 }),
    .d({open_n12816,\u2_Display/n766 }),
    .f({open_n12834,\u2_Display/n801 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2060|_al_u2061  (
    .b({\u2_Display/n769 [1],\u2_Display/n769 [2]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n765 ,\u2_Display/n764 }),
    .f({\u2_Display/n800 ,\u2_Display/n799 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2062|_al_u2063  (
    .b({\u2_Display/n769 [3],\u2_Display/n769 [4]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n763 ,\u2_Display/n762 }),
    .f({\u2_Display/n798 ,\u2_Display/n797 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2064|_al_u2065  (
    .b({\u2_Display/n769 [5],\u2_Display/n769 [6]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n761 ,\u2_Display/n760 }),
    .f({\u2_Display/n796 ,\u2_Display/n795 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2066|_al_u2069  (
    .b({\u2_Display/n769 [7],\u2_Display/n769 [10]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n759 ,\u2_Display/n756 }),
    .f({\u2_Display/n794 ,\u2_Display/n791 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2067|_al_u2068  (
    .b({\u2_Display/n769 [8],\u2_Display/n769 [9]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n758 ,\u2_Display/n757 }),
    .f({\u2_Display/n793 ,\u2_Display/n792 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2070|_al_u2071  (
    .b({\u2_Display/n769 [11],\u2_Display/n769 [12]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n755 ,\u2_Display/n754 }),
    .f({\u2_Display/n790 ,\u2_Display/n789 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2072|_al_u2073  (
    .b({\u2_Display/n769 [13],\u2_Display/n769 [14]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n753 ,\u2_Display/n752 }),
    .f({\u2_Display/n788 ,\u2_Display/n787 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2074|_al_u2075  (
    .b({\u2_Display/n769 [15],\u2_Display/n769 [16]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n751 ,\u2_Display/n750 }),
    .f({\u2_Display/n786 ,\u2_Display/n785 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2076|_al_u2077  (
    .b({\u2_Display/n769 [17],\u2_Display/n769 [18]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n749 ,\u2_Display/n748 }),
    .f({\u2_Display/n784 ,\u2_Display/n783 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2078|_al_u2079  (
    .b({\u2_Display/n769 [19],\u2_Display/n769 [20]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n747 ,\u2_Display/n746 }),
    .f({\u2_Display/n782 ,\u2_Display/n781 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2080|_al_u2081  (
    .b({\u2_Display/n769 [21],\u2_Display/n769 [22]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n745 ,\u2_Display/n744 }),
    .f({\u2_Display/n780 ,\u2_Display/n779 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2082|_al_u2085  (
    .b({\u2_Display/n769 [23],\u2_Display/n769 [26]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n743 ,\u2_Display/n740 }),
    .f({\u2_Display/n778 ,\u2_Display/n775 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u2083 (
    .b({open_n13130,\u2_Display/n769 [24]}),
    .c({open_n13131,\u2_Display/n767 }),
    .d({open_n13134,\u2_Display/n742 }),
    .f({open_n13152,\u2_Display/n777 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2084|_al_u2088  (
    .b({\u2_Display/n769 [25],\u2_Display/n769 [29]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n741 ,\u2_Display/n737 }),
    .f({\u2_Display/n776 ,\u2_Display/n772 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2086|_al_u2090  (
    .b({\u2_Display/n769 [27],\u2_Display/n769 [31]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n739 ,\u2_Display/n735 }),
    .f({\u2_Display/n774 ,\u2_Display/n770 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2087|_al_u2089  (
    .b({\u2_Display/n769 [28],\u2_Display/n769 [30]}),
    .c({\u2_Display/n767 ,\u2_Display/n767 }),
    .d({\u2_Display/n738 ,\u2_Display/n736 }),
    .f({\u2_Display/n773 ,\u2_Display/n771 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2091|_al_u2093  (
    .b({\u2_Display/n1892 [0],\u2_Display/n1892 [2]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1889 ,\u2_Display/n1887 }),
    .f({\u2_Display/n1924 ,\u2_Display/n1922 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2092|_al_u2096  (
    .b({\u2_Display/n1892 [1],\u2_Display/n1892 [5]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1888 ,\u2_Display/n1884 }),
    .f({\u2_Display/n1923 ,\u2_Display/n1919 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2094|_al_u2099  (
    .b({\u2_Display/n1892 [3],\u2_Display/n1892 [8]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1886 ,\u2_Display/n1881 }),
    .f({\u2_Display/n1921 ,\u2_Display/n1916 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2095|_al_u2097  (
    .b({\u2_Display/n1892 [4],\u2_Display/n1892 [6]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1885 ,\u2_Display/n1883 }),
    .f({\u2_Display/n1920 ,\u2_Display/n1918 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2098|_al_u2101  (
    .b({\u2_Display/n1892 [7],\u2_Display/n1892 [10]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1882 ,\u2_Display/n1879 }),
    .f({\u2_Display/n1917 ,\u2_Display/n1914 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2100|_al_u2104  (
    .b({\u2_Display/n1892 [9],\u2_Display/n1892 [13]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1880 ,\u2_Display/n1876 }),
    .f({\u2_Display/n1915 ,\u2_Display/n1911 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2102|_al_u2108  (
    .b({\u2_Display/n1892 [11],\u2_Display/n1892 [17]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1878 ,\u2_Display/n1872 }),
    .f({\u2_Display/n1913 ,\u2_Display/n1907 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2103|_al_u2105  (
    .b({\u2_Display/n1892 [12],\u2_Display/n1892 [14]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1877 ,\u2_Display/n1875 }),
    .f({\u2_Display/n1912 ,\u2_Display/n1910 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2106|_al_u2111  (
    .b({\u2_Display/n1892 [15],\u2_Display/n1892 [20]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1874 ,\u2_Display/n1869 }),
    .f({\u2_Display/n1909 ,\u2_Display/n1904 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2107|_al_u2109  (
    .b({\u2_Display/n1892 [16],\u2_Display/n1892 [18]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1873 ,\u2_Display/n1871 }),
    .f({\u2_Display/n1908 ,\u2_Display/n1906 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2110|_al_u2113  (
    .b({\u2_Display/n1892 [19],\u2_Display/n1892 [22]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1870 ,\u2_Display/n1867 }),
    .f({\u2_Display/n1905 ,\u2_Display/n1902 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2112|_al_u2116  (
    .b({\u2_Display/n1892 [21],\u2_Display/n1892 [25]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1868 ,\u2_Display/n1864 }),
    .f({\u2_Display/n1903 ,\u2_Display/n1899 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2114|_al_u2120  (
    .b({\u2_Display/n1892 [23],\u2_Display/n1892 [29]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1866 ,\u2_Display/n1860 }),
    .f({\u2_Display/n1901 ,\u2_Display/n1895 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2115|_al_u2117  (
    .b({\u2_Display/n1892 [24],\u2_Display/n1892 [26]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1865 ,\u2_Display/n1863 }),
    .f({\u2_Display/n1900 ,\u2_Display/n1898 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2118|_al_u2252  (
    .b({\u2_Display/n1892 [27],\u2_Display/n1927 [1]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1862 ,\u2_Display/n1923 }),
    .f({\u2_Display/n1897 ,\u2_Display/n1958 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2119|_al_u2121  (
    .b({\u2_Display/n1892 [28],\u2_Display/n1892 [30]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1890 }),
    .d({\u2_Display/n1861 ,\u2_Display/n1859 }),
    .f({\u2_Display/n1896 ,\u2_Display/n1894 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2122|_al_u2255  (
    .b({\u2_Display/n1892 [31],\u2_Display/n1927 [4]}),
    .c({\u2_Display/n1890 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1858 ,\u2_Display/n1920 }),
    .f({\u2_Display/n1893 ,\u2_Display/n1955 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2123|_al_u2125  (
    .b({\u2_Display/n3015 [0],\u2_Display/n3015 [2]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n3012 ,\u2_Display/n3010 }),
    .f({\u2_Display/n3047 ,\u2_Display/n3045 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2124|_al_u2128  (
    .b({\u2_Display/n3015 [1],\u2_Display/n3015 [5]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n3011 ,\u2_Display/n3007 }),
    .f({\u2_Display/n3046 ,\u2_Display/n3042 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2126|_al_u2131  (
    .b({\u2_Display/n3015 [3],\u2_Display/n3015 [8]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n3009 ,\u2_Display/n3004 }),
    .f({\u2_Display/n3044 ,\u2_Display/n3039 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2127|_al_u2129  (
    .b({\u2_Display/n3015 [4],\u2_Display/n3015 [6]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n3008 ,\u2_Display/n3006 }),
    .f({\u2_Display/n3043 ,\u2_Display/n3041 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2130|_al_u2133  (
    .b({\u2_Display/n3015 [7],\u2_Display/n3015 [10]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n3005 ,\u2_Display/n3002 }),
    .f({\u2_Display/n3040 ,\u2_Display/n3037 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2132|_al_u2136  (
    .b({\u2_Display/n3015 [9],\u2_Display/n3015 [13]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n3003 ,\u2_Display/n2999 }),
    .f({\u2_Display/n3038 ,\u2_Display/n3034 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2134|_al_u2139  (
    .b({\u2_Display/n3015 [11],\u2_Display/n3015 [16]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n3001 ,\u2_Display/n2996 }),
    .f({\u2_Display/n3036 ,\u2_Display/n3031 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2135|_al_u2137  (
    .b({\u2_Display/n3015 [12],\u2_Display/n3015 [14]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n3000 ,\u2_Display/n2998 }),
    .f({\u2_Display/n3035 ,\u2_Display/n3033 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2138|_al_u2141  (
    .b({\u2_Display/n3015 [15],\u2_Display/n3015 [18]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n2997 ,\u2_Display/n2994 }),
    .f({\u2_Display/n3032 ,\u2_Display/n3029 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2140|_al_u2144  (
    .b({\u2_Display/n3015 [17],\u2_Display/n3015 [21]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n2995 ,\u2_Display/n2991 }),
    .f({\u2_Display/n3030 ,\u2_Display/n3026 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2142|_al_u2147  (
    .b({\u2_Display/n3015 [19],\u2_Display/n3015 [24]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n2993 ,\u2_Display/n2988 }),
    .f({\u2_Display/n3028 ,\u2_Display/n3023 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2143|_al_u2145  (
    .b({\u2_Display/n3015 [20],\u2_Display/n3015 [22]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n2992 ,\u2_Display/n2990 }),
    .f({\u2_Display/n3027 ,\u2_Display/n3025 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2146|_al_u2149  (
    .b({\u2_Display/n3015 [23],\u2_Display/n3015 [26]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n2989 ,\u2_Display/n2986 }),
    .f({\u2_Display/n3024 ,\u2_Display/n3021 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2148|_al_u2151  (
    .b({\u2_Display/n3015 [25],\u2_Display/n3015 [28]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n2987 ,\u2_Display/n2984 }),
    .f({\u2_Display/n3022 ,\u2_Display/n3019 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2150|_al_u2153  (
    .b({\u2_Display/n3015 [27],\u2_Display/n3015 [30]}),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n2985 ,\u2_Display/n2982 }),
    .f({\u2_Display/n3020 ,\u2_Display/n3017 }));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1100101011001010),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2152|_al_u2154  (
    .a({open_n13996,\u2_Display/n3015 [31]}),
    .b({\u2_Display/n3015 [29],\u2_Display/n2981 }),
    .c({\u2_Display/n3013 ,\u2_Display/n3013 }),
    .d({\u2_Display/n2983 ,open_n13999}),
    .f({\u2_Display/n3018 ,\u2_Display/n3016 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2155|_al_u2160  (
    .b({\u2_Display/n4173 [0],\u2_Display/n4173 [5]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4170 ,\u2_Display/n4165 }),
    .f({\u2_Display/n4205 ,\u2_Display/n4200 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2156|_al_u2157  (
    .b({\u2_Display/n4173 [1],\u2_Display/n4173 [2]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4169 ,\u2_Display/n4168 }),
    .f({\u2_Display/n4204 ,\u2_Display/n4203 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2158|_al_u2163  (
    .b({\u2_Display/n4173 [3],\u2_Display/n4173 [8]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4167 ,\u2_Display/n4162 }),
    .f({\u2_Display/n4202 ,\u2_Display/n4197 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2159|_al_u2161  (
    .b({\u2_Display/n4173 [4],\u2_Display/n4173 [6]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4166 ,\u2_Display/n4164 }),
    .f({\u2_Display/n4201 ,\u2_Display/n4199 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2162|_al_u2165  (
    .b({\u2_Display/n4173 [7],\u2_Display/n4173 [10]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4163 ,\u2_Display/n4160 }),
    .f({\u2_Display/n4198 ,\u2_Display/n4195 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2164|_al_u2167  (
    .b({\u2_Display/n4173 [9],\u2_Display/n4173 [12]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4161 ,\u2_Display/n4158 }),
    .f({\u2_Display/n4196 ,\u2_Display/n4193 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2166|_al_u2169  (
    .b({\u2_Display/n4173 [11],\u2_Display/n4173 [14]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4159 ,\u2_Display/n4156 }),
    .f({\u2_Display/n4194 ,\u2_Display/n4191 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2168|_al_u2172  (
    .b({\u2_Display/n4173 [13],\u2_Display/n4153 }),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4157 ,\u2_Display/n4173 [17]}),
    .f({\u2_Display/n4192 ,\u2_Display/n4188 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2170|_al_u2176  (
    .b({\u2_Display/n4173 [15],\u2_Display/n4173 [21]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4155 ,\u2_Display/n4149 }),
    .f({\u2_Display/n4190 ,\u2_Display/n4184 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2171|_al_u2173  (
    .b({\u2_Display/n4173 [16],\u2_Display/n4173 [18]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4154 ,\u2_Display/n4152 }),
    .f({\u2_Display/n4189 ,\u2_Display/n4187 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2174|_al_u2179  (
    .b({\u2_Display/n4173 [19],\u2_Display/n4173 [24]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4151 ,\u2_Display/n4146 }),
    .f({\u2_Display/n4186 ,\u2_Display/n4181 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2175|_al_u2177  (
    .b({\u2_Display/n4173 [20],\u2_Display/n4173 [22]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4150 ,\u2_Display/n4148 }),
    .f({\u2_Display/n4185 ,\u2_Display/n4183 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2178|_al_u2181  (
    .b({\u2_Display/n4173 [23],\u2_Display/n4173 [26]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4147 ,\u2_Display/n4144 }),
    .f({\u2_Display/n4182 ,\u2_Display/n4179 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2180|_al_u2183  (
    .b({\u2_Display/n4173 [25],\u2_Display/n4173 [28]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4145 ,\u2_Display/n4142 }),
    .f({\u2_Display/n4180 ,\u2_Display/n4177 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2182|_al_u2185  (
    .b({\u2_Display/n4173 [27],\u2_Display/n4173 [30]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4143 ,\u2_Display/n4140 }),
    .f({\u2_Display/n4178 ,\u2_Display/n4175 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2184|_al_u2186  (
    .b({\u2_Display/n4173 [29],\u2_Display/n4173 [31]}),
    .c({\u2_Display/n4171 ,\u2_Display/n4171 }),
    .d({\u2_Display/n4141 ,\u2_Display/n4139 }),
    .f({\u2_Display/n4176 ,\u2_Display/n4174 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2187|_al_u2191  (
    .b({\u2_Display/n5296 [0],\u2_Display/n5296 [4]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5293 ,\u2_Display/n5289 }),
    .f({\u2_Display/n5328 ,\u2_Display/n5324 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2188|_al_u2189  (
    .b({\u2_Display/n5296 [1],\u2_Display/n5296 [2]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5292 ,\u2_Display/n5291 }),
    .f({\u2_Display/n5327 ,\u2_Display/n5326 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2190|_al_u2193  (
    .b({\u2_Display/n5296 [3],\u2_Display/n5296 [6]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5290 ,\u2_Display/n5287 }),
    .f({\u2_Display/n5325 ,\u2_Display/n5322 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2192|_al_u2196  (
    .b({\u2_Display/n5296 [5],\u2_Display/n5296 [9]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5288 ,\u2_Display/n5284 }),
    .f({\u2_Display/n5323 ,\u2_Display/n5319 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2194|_al_u2199  (
    .b({\u2_Display/n5296 [7],\u2_Display/n5296 [12]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5286 ,\u2_Display/n5281 }),
    .f({\u2_Display/n5321 ,\u2_Display/n5316 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2195|_al_u2197  (
    .b({\u2_Display/n5296 [8],\u2_Display/n5296 [10]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5285 ,\u2_Display/n5283 }),
    .f({\u2_Display/n5320 ,\u2_Display/n5318 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2198|_al_u2201  (
    .b({\u2_Display/n5296 [11],\u2_Display/n5296 [14]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5282 ,\u2_Display/n5279 }),
    .f({\u2_Display/n5317 ,\u2_Display/n5314 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2200|_al_u2204  (
    .b({\u2_Display/n5296 [13],\u2_Display/n5296 [17]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5280 ,\u2_Display/n5276 }),
    .f({\u2_Display/n5315 ,\u2_Display/n5311 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2202|_al_u2207  (
    .b({\u2_Display/n5296 [15],\u2_Display/n5296 [20]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5278 ,\u2_Display/n5273 }),
    .f({\u2_Display/n5313 ,\u2_Display/n5308 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2203|_al_u2205  (
    .b({\u2_Display/n5296 [16],\u2_Display/n5296 [18]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5277 ,\u2_Display/n5275 }),
    .f({\u2_Display/n5312 ,\u2_Display/n5310 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2206|_al_u2211  (
    .b({\u2_Display/n5296 [19],\u2_Display/n5296 [24]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5274 ,\u2_Display/n5269 }),
    .f({\u2_Display/n5309 ,\u2_Display/n5304 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2208|_al_u2209  (
    .b({\u2_Display/n5296 [21],\u2_Display/n5296 [22]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5272 ,\u2_Display/n5271 }),
    .f({\u2_Display/n5307 ,\u2_Display/n5306 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2210|_al_u2213  (
    .b({\u2_Display/n5296 [23],\u2_Display/n5296 [26]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5270 ,\u2_Display/n5267 }),
    .f({\u2_Display/n5305 ,\u2_Display/n5302 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2212|_al_u2348  (
    .b({\u2_Display/n5296 [25],\u2_Display/n5331 [1]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5268 ,\u2_Display/n5327 }),
    .f({\u2_Display/n5303 ,\u2_Display/n5362 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2214|_al_u2215  (
    .b({\u2_Display/n5296 [27],\u2_Display/n5296 [28]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5266 ,\u2_Display/n5265 }),
    .f({\u2_Display/n5301 ,\u2_Display/n5300 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2216|_al_u2217  (
    .b({\u2_Display/n5296 [29],\u2_Display/n5296 [30]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5294 }),
    .d({\u2_Display/n5264 ,\u2_Display/n5263 }),
    .f({\u2_Display/n5299 ,\u2_Display/n5298 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2218|_al_u2356  (
    .b({\u2_Display/n5296 [31],\u2_Display/n5331 [9]}),
    .c({\u2_Display/n5294 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5262 ,\u2_Display/n5319 }),
    .f({\u2_Display/n5297 ,\u2_Display/n5354 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2219|_al_u2224  (
    .b({\u2_Display/n804 [0],\u2_Display/n804 [5]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n801 ,\u2_Display/n796 }),
    .f({\u2_Display/n836 ,\u2_Display/n831 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2220|_al_u2221  (
    .b({\u2_Display/n804 [1],\u2_Display/n804 [2]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n800 ,\u2_Display/n799 }),
    .f({\u2_Display/n835 ,\u2_Display/n834 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2222|_al_u2227  (
    .b({\u2_Display/n804 [3],\u2_Display/n804 [8]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n798 ,\u2_Display/n793 }),
    .f({\u2_Display/n833 ,\u2_Display/n828 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2223|_al_u2225  (
    .b({\u2_Display/n804 [4],\u2_Display/n804 [6]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n797 ,\u2_Display/n795 }),
    .f({\u2_Display/n832 ,\u2_Display/n830 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2226|_al_u2229  (
    .b({\u2_Display/n804 [7],\u2_Display/n804 [10]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n794 ,\u2_Display/n791 }),
    .f({\u2_Display/n829 ,\u2_Display/n826 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2228|_al_u2231  (
    .b({\u2_Display/n804 [9],\u2_Display/n804 [12]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n792 ,\u2_Display/n789 }),
    .f({\u2_Display/n827 ,\u2_Display/n824 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2230|_al_u2233  (
    .b({\u2_Display/n804 [11],\u2_Display/n804 [14]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n790 ,\u2_Display/n787 }),
    .f({\u2_Display/n825 ,\u2_Display/n822 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2232|_al_u2235  (
    .b({\u2_Display/n804 [13],\u2_Display/n804 [16]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n788 ,\u2_Display/n785 }),
    .f({\u2_Display/n823 ,\u2_Display/n820 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2234|_al_u2237  (
    .b({\u2_Display/n804 [15],\u2_Display/n804 [18]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n786 ,\u2_Display/n783 }),
    .f({\u2_Display/n821 ,\u2_Display/n818 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2236|_al_u2239  (
    .b({\u2_Display/n804 [17],\u2_Display/n804 [20]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n784 ,\u2_Display/n781 }),
    .f({\u2_Display/n819 ,\u2_Display/n816 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2238|_al_u2241  (
    .b({\u2_Display/n804 [19],\u2_Display/n804 [22]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n782 ,\u2_Display/n779 }),
    .f({\u2_Display/n817 ,\u2_Display/n814 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2240|_al_u2244  (
    .b({\u2_Display/n804 [21],\u2_Display/n804 [25]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n780 ,\u2_Display/n776 }),
    .f({\u2_Display/n815 ,\u2_Display/n811 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2242|_al_u2247  (
    .b({\u2_Display/n804 [23],\u2_Display/n804 [28]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n778 ,\u2_Display/n773 }),
    .f({\u2_Display/n813 ,\u2_Display/n808 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2243|_al_u2245  (
    .b({\u2_Display/n804 [24],\u2_Display/n804 [26]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n777 ,\u2_Display/n775 }),
    .f({\u2_Display/n812 ,\u2_Display/n810 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2246|_al_u2249  (
    .b({\u2_Display/n804 [27],\u2_Display/n804 [30]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n774 ,\u2_Display/n771 }),
    .f({\u2_Display/n809 ,\u2_Display/n806 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2248|_al_u2250  (
    .b({\u2_Display/n804 [29],\u2_Display/n804 [31]}),
    .c({\u2_Display/n802 ,\u2_Display/n802 }),
    .d({\u2_Display/n772 ,\u2_Display/n770 }),
    .f({\u2_Display/n807 ,\u2_Display/n805 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2251|_al_u2253  (
    .b({\u2_Display/n1927 [0],\u2_Display/n1927 [2]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1924 ,\u2_Display/n1922 }),
    .f({\u2_Display/n1959 ,\u2_Display/n1957 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2254|_al_u2257  (
    .b({\u2_Display/n1927 [3],\u2_Display/n1927 [6]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1921 ,\u2_Display/n1918 }),
    .f({\u2_Display/n1956 ,\u2_Display/n1953 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2256|_al_u2259  (
    .b({\u2_Display/n1927 [5],\u2_Display/n1927 [8]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1919 ,\u2_Display/n1916 }),
    .f({\u2_Display/n1954 ,\u2_Display/n1951 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2258|_al_u2261  (
    .b({\u2_Display/n1927 [7],\u2_Display/n1927 [10]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1917 ,\u2_Display/n1914 }),
    .f({\u2_Display/n1952 ,\u2_Display/n1949 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2260|_al_u2263  (
    .b({\u2_Display/n1927 [9],\u2_Display/n1927 [12]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1915 ,\u2_Display/n1912 }),
    .f({\u2_Display/n1950 ,\u2_Display/n1947 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2262|_al_u2265  (
    .b({\u2_Display/n1927 [11],\u2_Display/n1927 [14]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1913 ,\u2_Display/n1910 }),
    .f({\u2_Display/n1948 ,\u2_Display/n1945 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2264|_al_u2267  (
    .b({\u2_Display/n1927 [13],\u2_Display/n1927 [16]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1911 ,\u2_Display/n1908 }),
    .f({\u2_Display/n1946 ,\u2_Display/n1943 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2266|_al_u2269  (
    .b({\u2_Display/n1927 [15],\u2_Display/n1927 [18]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1909 ,\u2_Display/n1906 }),
    .f({\u2_Display/n1944 ,\u2_Display/n1941 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2268|_al_u2271  (
    .b({\u2_Display/n1927 [17],\u2_Display/n1927 [20]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1907 ,\u2_Display/n1904 }),
    .f({\u2_Display/n1942 ,\u2_Display/n1939 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2270|_al_u2273  (
    .b({\u2_Display/n1927 [19],\u2_Display/n1927 [22]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1905 ,\u2_Display/n1902 }),
    .f({\u2_Display/n1940 ,\u2_Display/n1937 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2272|_al_u2275  (
    .b({\u2_Display/n1927 [21],\u2_Display/n1927 [24]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1903 ,\u2_Display/n1900 }),
    .f({\u2_Display/n1938 ,\u2_Display/n1935 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2274|_al_u2277  (
    .b({\u2_Display/n1927 [23],\u2_Display/n1927 [26]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1901 ,\u2_Display/n1898 }),
    .f({\u2_Display/n1936 ,\u2_Display/n1933 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2276|_al_u2279  (
    .b({\u2_Display/n1927 [25],\u2_Display/n1927 [28]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1899 ,\u2_Display/n1896 }),
    .f({\u2_Display/n1934 ,\u2_Display/n1931 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2278|_al_u2281  (
    .b({\u2_Display/n1927 [27],\u2_Display/n1927 [30]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1897 ,\u2_Display/n1894 }),
    .f({\u2_Display/n1932 ,\u2_Display/n1929 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2280|_al_u2282  (
    .b({\u2_Display/n1927 [29],\u2_Display/n1927 [31]}),
    .c({\u2_Display/n1925 ,\u2_Display/n1925 }),
    .d({\u2_Display/n1895 ,\u2_Display/n1893 }),
    .f({\u2_Display/n1930 ,\u2_Display/n1928 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2283|_al_u2288  (
    .b({\u2_Display/n3050 [0],\u2_Display/n3050 [5]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3047 ,\u2_Display/n3042 }),
    .f({\u2_Display/n3082 ,\u2_Display/n3077 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2284|_al_u2285  (
    .b({\u2_Display/n3050 [1],\u2_Display/n3050 [2]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3046 ,\u2_Display/n3045 }),
    .f({\u2_Display/n3081 ,\u2_Display/n3080 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u2286|_al_u2291  (
    .b({\u2_Display/n3048 ,\u2_Display/n3050 [8]}),
    .c({\u2_Display/n3050 [3],\u2_Display/n3048 }),
    .d({\u2_Display/n3044 ,\u2_Display/n3039 }),
    .f({\u2_Display/n3079 ,\u2_Display/n3074 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2287|_al_u2289  (
    .b({\u2_Display/n3050 [4],\u2_Display/n3050 [6]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3043 ,\u2_Display/n3041 }),
    .f({\u2_Display/n3078 ,\u2_Display/n3076 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2290|_al_u2293  (
    .b({\u2_Display/n3050 [7],\u2_Display/n3050 [10]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3040 ,\u2_Display/n3037 }),
    .f({\u2_Display/n3075 ,\u2_Display/n3072 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2292|_al_u2296  (
    .b({\u2_Display/n3050 [9],\u2_Display/n3050 [13]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3038 ,\u2_Display/n3034 }),
    .f({\u2_Display/n3073 ,\u2_Display/n3069 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2294|_al_u2300  (
    .b({\u2_Display/n3050 [11],\u2_Display/n3030 }),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3036 ,\u2_Display/n3050 [17]}),
    .f({\u2_Display/n3071 ,\u2_Display/n3065 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2295|_al_u2297  (
    .b({\u2_Display/n3050 [12],\u2_Display/n3050 [14]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3035 ,\u2_Display/n3033 }),
    .f({\u2_Display/n3070 ,\u2_Display/n3068 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2298|_al_u2303  (
    .b({\u2_Display/n3050 [15],\u2_Display/n3050 [20]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3032 ,\u2_Display/n3027 }),
    .f({\u2_Display/n3067 ,\u2_Display/n3062 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2299|_al_u2301  (
    .b({\u2_Display/n3050 [16],\u2_Display/n3050 [18]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3031 ,\u2_Display/n3029 }),
    .f({\u2_Display/n3066 ,\u2_Display/n3064 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2302|_al_u2305  (
    .b({\u2_Display/n3050 [19],\u2_Display/n3050 [22]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3028 ,\u2_Display/n3025 }),
    .f({\u2_Display/n3063 ,\u2_Display/n3060 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2304|_al_u2308  (
    .b({\u2_Display/n3050 [21],\u2_Display/n3050 [25]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3026 ,\u2_Display/n3022 }),
    .f({\u2_Display/n3061 ,\u2_Display/n3057 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2306|_al_u2312  (
    .b({\u2_Display/n3050 [23],\u2_Display/n3050 [29]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3024 ,\u2_Display/n3018 }),
    .f({\u2_Display/n3059 ,\u2_Display/n3053 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2307|_al_u2309  (
    .b({\u2_Display/n3050 [24],\u2_Display/n3050 [26]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3023 ,\u2_Display/n3021 }),
    .f({\u2_Display/n3058 ,\u2_Display/n3056 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2310|_al_u2314  (
    .b({\u2_Display/n3050 [27],\u2_Display/n3050 [31]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3020 ,\u2_Display/n3016 }),
    .f({\u2_Display/n3055 ,\u2_Display/n3051 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2311|_al_u2313  (
    .b({\u2_Display/n3050 [28],\u2_Display/n3050 [30]}),
    .c({\u2_Display/n3048 ,\u2_Display/n3048 }),
    .d({\u2_Display/n3019 ,\u2_Display/n3017 }),
    .f({\u2_Display/n3054 ,\u2_Display/n3052 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2315|_al_u2317  (
    .b({\u2_Display/n4208 [0],\u2_Display/n4208 [2]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4205 ,\u2_Display/n4203 }),
    .f({\u2_Display/n4240 ,\u2_Display/n4238 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2316|_al_u2319  (
    .b({\u2_Display/n4208 [1],\u2_Display/n4208 [4]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4204 ,\u2_Display/n4201 }),
    .f({\u2_Display/n4239 ,\u2_Display/n4236 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2318|_al_u2321  (
    .b({\u2_Display/n4208 [3],\u2_Display/n4208 [6]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4202 ,\u2_Display/n4199 }),
    .f({\u2_Display/n4237 ,\u2_Display/n4234 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2320|_al_u2324  (
    .b({\u2_Display/n4208 [5],\u2_Display/n4208 [9]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4200 ,\u2_Display/n4196 }),
    .f({\u2_Display/n4235 ,\u2_Display/n4231 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2322|_al_u2327  (
    .b({\u2_Display/n4208 [7],\u2_Display/n4208 [12]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4198 ,\u2_Display/n4193 }),
    .f({\u2_Display/n4233 ,\u2_Display/n4228 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2323|_al_u2325  (
    .b({\u2_Display/n4208 [8],\u2_Display/n4208 [10]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4197 ,\u2_Display/n4195 }),
    .f({\u2_Display/n4232 ,\u2_Display/n4230 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2326|_al_u2329  (
    .b({\u2_Display/n4208 [11],\u2_Display/n4208 [14]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4194 ,\u2_Display/n4191 }),
    .f({\u2_Display/n4229 ,\u2_Display/n4226 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2328|_al_u2331  (
    .b({\u2_Display/n4208 [13],\u2_Display/n4208 [16]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4192 ,\u2_Display/n4189 }),
    .f({\u2_Display/n4227 ,\u2_Display/n4224 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2330|_al_u2333  (
    .b({\u2_Display/n4208 [15],\u2_Display/n4208 [18]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4190 ,\u2_Display/n4187 }),
    .f({\u2_Display/n4225 ,\u2_Display/n4222 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2332|_al_u2336  (
    .b({\u2_Display/n4208 [17],\u2_Display/n4208 [21]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4188 ,\u2_Display/n4184 }),
    .f({\u2_Display/n4223 ,\u2_Display/n4219 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2334|_al_u2340  (
    .b({\u2_Display/n4208 [19],\u2_Display/n4208 [25]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4186 ,\u2_Display/n4180 }),
    .f({\u2_Display/n4221 ,\u2_Display/n4215 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2335|_al_u2337  (
    .b({\u2_Display/n4208 [20],\u2_Display/n4208 [22]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4185 ,\u2_Display/n4183 }),
    .f({\u2_Display/n4220 ,\u2_Display/n4218 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2338|_al_u2344  (
    .b({\u2_Display/n4208 [23],\u2_Display/n4208 [29]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4182 ,\u2_Display/n4176 }),
    .f({\u2_Display/n4217 ,\u2_Display/n4211 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2339|_al_u2341  (
    .b({\u2_Display/n4208 [24],\u2_Display/n4208 [26]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4181 ,\u2_Display/n4179 }),
    .f({\u2_Display/n4216 ,\u2_Display/n4214 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2342|_al_u2476  (
    .b({\u2_Display/n4208 [27],\u2_Display/n4243 [1]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4178 ,\u2_Display/n4239 }),
    .f({\u2_Display/n4213 ,\u2_Display/n4274 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2343|_al_u2345  (
    .b({\u2_Display/n4208 [28],\u2_Display/n4208 [30]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4206 }),
    .d({\u2_Display/n4177 ,\u2_Display/n4175 }),
    .f({\u2_Display/n4212 ,\u2_Display/n4210 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2346|_al_u2484  (
    .b({\u2_Display/n4208 [31],\u2_Display/n4243 [9]}),
    .c({\u2_Display/n4206 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4174 ,\u2_Display/n4231 }),
    .f({\u2_Display/n4209 ,\u2_Display/n4266 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2347|_al_u2349  (
    .b({\u2_Display/n5331 [0],\u2_Display/n5331 [2]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5328 ,\u2_Display/n5326 }),
    .f({\u2_Display/n5363 ,\u2_Display/n5361 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2350|_al_u2353  (
    .b({\u2_Display/n5331 [3],\u2_Display/n5331 [6]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5325 ,\u2_Display/n5322 }),
    .f({\u2_Display/n5360 ,\u2_Display/n5357 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2351|_al_u2352  (
    .b({\u2_Display/n5331 [4],\u2_Display/n5331 [5]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5324 ,\u2_Display/n5323 }),
    .f({\u2_Display/n5359 ,\u2_Display/n5358 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2354|_al_u2360  (
    .b({\u2_Display/n5331 [7],\u2_Display/n5331 [13]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5321 ,\u2_Display/n5315 }),
    .f({\u2_Display/n5356 ,\u2_Display/n5350 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2355|_al_u2357  (
    .b({\u2_Display/n5331 [8],\u2_Display/n5331 [10]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5320 ,\u2_Display/n5318 }),
    .f({\u2_Display/n5355 ,\u2_Display/n5353 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2358|_al_u2364  (
    .b({\u2_Display/n5331 [11],\u2_Display/n5331 [17]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5317 ,\u2_Display/n5311 }),
    .f({\u2_Display/n5352 ,\u2_Display/n5346 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2359|_al_u2361  (
    .b({\u2_Display/n5331 [12],\u2_Display/n5331 [14]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5316 ,\u2_Display/n5314 }),
    .f({\u2_Display/n5351 ,\u2_Display/n5349 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2362|_al_u2367  (
    .b({\u2_Display/n5331 [15],\u2_Display/n5331 [20]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5313 ,\u2_Display/n5308 }),
    .f({\u2_Display/n5348 ,\u2_Display/n5343 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2363|_al_u2365  (
    .b({\u2_Display/n5331 [16],\u2_Display/n5331 [18]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5312 ,\u2_Display/n5310 }),
    .f({\u2_Display/n5347 ,\u2_Display/n5345 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2366|_al_u2369  (
    .b({\u2_Display/n5331 [19],\u2_Display/n5331 [22]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5309 ,\u2_Display/n5306 }),
    .f({\u2_Display/n5344 ,\u2_Display/n5341 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2368|_al_u2372  (
    .b({\u2_Display/n5331 [21],\u2_Display/n5331 [25]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5307 ,\u2_Display/n5303 }),
    .f({\u2_Display/n5342 ,\u2_Display/n5338 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2370|_al_u2376  (
    .b({\u2_Display/n5331 [23],\u2_Display/n5331 [29]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5305 ,\u2_Display/n5299 }),
    .f({\u2_Display/n5340 ,\u2_Display/n5334 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2371|_al_u2373  (
    .b({\u2_Display/n5331 [24],\u2_Display/n5331 [26]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5304 ,\u2_Display/n5302 }),
    .f({\u2_Display/n5339 ,\u2_Display/n5337 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2374|_al_u2378  (
    .b({\u2_Display/n5331 [27],\u2_Display/n5331 [31]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5301 ,\u2_Display/n5297 }),
    .f({\u2_Display/n5336 ,\u2_Display/n5332 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2375|_al_u2377  (
    .b({\u2_Display/n5331 [28],\u2_Display/n5331 [30]}),
    .c({\u2_Display/n5329 ,\u2_Display/n5329 }),
    .d({\u2_Display/n5300 ,\u2_Display/n5298 }),
    .f({\u2_Display/n5335 ,\u2_Display/n5333 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2379|_al_u2381  (
    .b({\u2_Display/n839 [0],\u2_Display/n839 [2]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n836 ,\u2_Display/n834 }),
    .f({\u2_Display/n871 ,\u2_Display/n869 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u2380 (
    .b({open_n16738,\u2_Display/n839 [1]}),
    .c({open_n16739,\u2_Display/n837 }),
    .d({open_n16742,\u2_Display/n835 }),
    .f({open_n16760,\u2_Display/n870 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2382|_al_u2385  (
    .b({\u2_Display/n839 [3],\u2_Display/n839 [6]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n833 ,\u2_Display/n830 }),
    .f({\u2_Display/n868 ,\u2_Display/n865 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2383|_al_u2384  (
    .b({\u2_Display/n839 [4],\u2_Display/n839 [5]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n832 ,\u2_Display/n831 }),
    .f({\u2_Display/n867 ,\u2_Display/n866 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2386|_al_u2387  (
    .b({\u2_Display/n839 [7],\u2_Display/n839 [8]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n829 ,\u2_Display/n828 }),
    .f({\u2_Display/n864 ,\u2_Display/n863 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2388|_al_u2389  (
    .b({\u2_Display/n839 [9],\u2_Display/n839 [10]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n827 ,\u2_Display/n826 }),
    .f({\u2_Display/n862 ,\u2_Display/n861 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2390|_al_u2391  (
    .b({\u2_Display/n839 [11],\u2_Display/n839 [12]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n825 ,\u2_Display/n824 }),
    .f({\u2_Display/n860 ,\u2_Display/n859 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2392|_al_u2393  (
    .b({\u2_Display/n839 [13],\u2_Display/n839 [14]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n823 ,\u2_Display/n822 }),
    .f({\u2_Display/n858 ,\u2_Display/n857 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2394|_al_u2395  (
    .b({\u2_Display/n839 [15],\u2_Display/n839 [16]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n821 ,\u2_Display/n820 }),
    .f({\u2_Display/n856 ,\u2_Display/n855 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2396|_al_u2397  (
    .b({\u2_Display/n839 [17],\u2_Display/n839 [18]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n819 ,\u2_Display/n818 }),
    .f({\u2_Display/n854 ,\u2_Display/n853 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2398|_al_u2399  (
    .b({\u2_Display/n839 [19],\u2_Display/n839 [20]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n817 ,\u2_Display/n816 }),
    .f({\u2_Display/n852 ,\u2_Display/n851 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2400|_al_u2401  (
    .b({\u2_Display/n839 [21],\u2_Display/n839 [22]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n815 ,\u2_Display/n814 }),
    .f({\u2_Display/n850 ,\u2_Display/n849 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2402|_al_u2408  (
    .b({\u2_Display/n839 [23],\u2_Display/n839 [29]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n813 ,\u2_Display/n807 }),
    .f({\u2_Display/n848 ,\u2_Display/n842 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2403|_al_u2405  (
    .b({\u2_Display/n839 [24],\u2_Display/n839 [26]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n812 ,\u2_Display/n810 }),
    .f({\u2_Display/n847 ,\u2_Display/n845 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u2404 (
    .b({open_n17052,\u2_Display/n839 [25]}),
    .c({open_n17053,\u2_Display/n837 }),
    .d({open_n17056,\u2_Display/n811 }),
    .f({open_n17074,\u2_Display/n846 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2406|_al_u2410  (
    .b({\u2_Display/n839 [27],\u2_Display/n839 [31]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n809 ,\u2_Display/n805 }),
    .f({\u2_Display/n844 ,\u2_Display/n840 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2407|_al_u2409  (
    .b({\u2_Display/n839 [28],\u2_Display/n839 [30]}),
    .c({\u2_Display/n837 ,\u2_Display/n837 }),
    .d({\u2_Display/n808 ,\u2_Display/n806 }),
    .f({\u2_Display/n843 ,\u2_Display/n841 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2411|_al_u2413  (
    .b({\u2_Display/n1962 [0],\u2_Display/n1962 [2]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1959 ,\u2_Display/n1957 }),
    .f({\u2_Display/n1994 ,\u2_Display/n1992 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2412|_al_u2415  (
    .b({\u2_Display/n1962 [1],\u2_Display/n1962 [4]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1958 ,\u2_Display/n1955 }),
    .f({\u2_Display/n1993 ,\u2_Display/n1990 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2414|_al_u2417  (
    .b({\u2_Display/n1962 [3],\u2_Display/n1962 [6]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1956 ,\u2_Display/n1953 }),
    .f({\u2_Display/n1991 ,\u2_Display/n1988 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2416|_al_u2419  (
    .b({\u2_Display/n1962 [5],\u2_Display/n1962 [8]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1954 ,\u2_Display/n1951 }),
    .f({\u2_Display/n1989 ,\u2_Display/n1986 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2418|_al_u2421  (
    .b({\u2_Display/n1962 [7],\u2_Display/n1962 [10]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1952 ,\u2_Display/n1949 }),
    .f({\u2_Display/n1987 ,\u2_Display/n1984 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2420|_al_u2423  (
    .b({\u2_Display/n1962 [9],\u2_Display/n1962 [12]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1950 ,\u2_Display/n1947 }),
    .f({\u2_Display/n1985 ,\u2_Display/n1982 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2422|_al_u2425  (
    .b({\u2_Display/n1962 [11],\u2_Display/n1962 [14]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1948 ,\u2_Display/n1945 }),
    .f({\u2_Display/n1983 ,\u2_Display/n1980 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2424|_al_u2428  (
    .b({\u2_Display/n1962 [13],\u2_Display/n1962 [17]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1946 ,\u2_Display/n1942 }),
    .f({\u2_Display/n1981 ,\u2_Display/n1977 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2426|_al_u2432  (
    .b({\u2_Display/n1962 [15],\u2_Display/n1962 [21]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1944 ,\u2_Display/n1938 }),
    .f({\u2_Display/n1979 ,\u2_Display/n1973 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2427|_al_u2429  (
    .b({\u2_Display/n1962 [16],\u2_Display/n1962 [18]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1943 ,\u2_Display/n1941 }),
    .f({\u2_Display/n1978 ,\u2_Display/n1976 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2430|_al_u2436  (
    .b({\u2_Display/n1962 [19],\u2_Display/n1962 [25]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1940 ,\u2_Display/n1934 }),
    .f({\u2_Display/n1975 ,\u2_Display/n1969 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2431|_al_u2433  (
    .b({\u2_Display/n1962 [20],\u2_Display/n1962 [22]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1939 ,\u2_Display/n1937 }),
    .f({\u2_Display/n1974 ,\u2_Display/n1972 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2434|_al_u2440  (
    .b({\u2_Display/n1962 [23],\u2_Display/n1962 [29]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1936 ,\u2_Display/n1930 }),
    .f({\u2_Display/n1971 ,\u2_Display/n1965 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2435|_al_u2437  (
    .b({\u2_Display/n1962 [24],\u2_Display/n1962 [26]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1935 ,\u2_Display/n1933 }),
    .f({\u2_Display/n1970 ,\u2_Display/n1968 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2438|_al_u2572  (
    .b({\u2_Display/n1962 [27],\u2_Display/n1997 [1]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1932 ,\u2_Display/n1993 }),
    .f({\u2_Display/n1967 ,\u2_Display/n2028 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2439|_al_u2441  (
    .b({\u2_Display/n1962 [28],\u2_Display/n1962 [30]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1960 }),
    .d({\u2_Display/n1931 ,\u2_Display/n1929 }),
    .f({\u2_Display/n1966 ,\u2_Display/n1964 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2442|_al_u2580  (
    .b({\u2_Display/n1962 [31],\u2_Display/n1997 [9]}),
    .c({\u2_Display/n1960 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1928 ,\u2_Display/n1985 }),
    .f({\u2_Display/n1963 ,\u2_Display/n2020 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2443|_al_u2445  (
    .b({\u2_Display/n3085 [0],\u2_Display/n3085 [2]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3082 ,\u2_Display/n3080 }),
    .f({\u2_Display/n3117 ,\u2_Display/n3115 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2444|_al_u2447  (
    .b({\u2_Display/n3085 [1],\u2_Display/n3085 [4]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3081 ,\u2_Display/n3078 }),
    .f({\u2_Display/n3116 ,\u2_Display/n3113 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2446|_al_u2449  (
    .b({\u2_Display/n3085 [3],\u2_Display/n3085 [6]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3079 ,\u2_Display/n3076 }),
    .f({\u2_Display/n3114 ,\u2_Display/n3111 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2448|_al_u2451  (
    .b({\u2_Display/n3085 [5],\u2_Display/n3085 [8]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3077 ,\u2_Display/n3074 }),
    .f({\u2_Display/n3112 ,\u2_Display/n3109 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2450|_al_u2453  (
    .b({\u2_Display/n3085 [7],\u2_Display/n3085 [10]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3075 ,\u2_Display/n3072 }),
    .f({\u2_Display/n3110 ,\u2_Display/n3107 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2452|_al_u2456  (
    .b({\u2_Display/n3085 [9],\u2_Display/n3085 [13]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3073 ,\u2_Display/n3069 }),
    .f({\u2_Display/n3108 ,\u2_Display/n3104 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2454|_al_u2459  (
    .b({\u2_Display/n3085 [11],\u2_Display/n3085 [16]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3071 ,\u2_Display/n3066 }),
    .f({\u2_Display/n3106 ,\u2_Display/n3101 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2455|_al_u2457  (
    .b({\u2_Display/n3085 [12],\u2_Display/n3085 [14]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3070 ,\u2_Display/n3068 }),
    .f({\u2_Display/n3105 ,\u2_Display/n3103 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2458|_al_u2461  (
    .b({\u2_Display/n3085 [15],\u2_Display/n3085 [18]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3067 ,\u2_Display/n3064 }),
    .f({\u2_Display/n3102 ,\u2_Display/n3099 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2460|_al_u2464  (
    .b({\u2_Display/n3085 [17],\u2_Display/n3085 [21]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3065 ,\u2_Display/n3061 }),
    .f({\u2_Display/n3100 ,\u2_Display/n3096 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2462|_al_u2468  (
    .b({\u2_Display/n3085 [19],\u2_Display/n3085 [25]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3063 ,\u2_Display/n3057 }),
    .f({\u2_Display/n3098 ,\u2_Display/n3092 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2463|_al_u2465  (
    .b({\u2_Display/n3085 [20],\u2_Display/n3085 [22]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3062 ,\u2_Display/n3060 }),
    .f({\u2_Display/n3097 ,\u2_Display/n3095 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2466|_al_u2471  (
    .b({\u2_Display/n3085 [23],\u2_Display/n3085 [28]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3059 ,\u2_Display/n3054 }),
    .f({\u2_Display/n3094 ,\u2_Display/n3089 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2467|_al_u2469  (
    .b({\u2_Display/n3085 [24],\u2_Display/n3085 [26]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3058 ,\u2_Display/n3056 }),
    .f({\u2_Display/n3093 ,\u2_Display/n3091 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2470|_al_u2473  (
    .b({\u2_Display/n3085 [27],\u2_Display/n3085 [30]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3055 ,\u2_Display/n3052 }),
    .f({\u2_Display/n3090 ,\u2_Display/n3087 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2472|_al_u2474  (
    .b({\u2_Display/n3085 [29],\u2_Display/n3085 [31]}),
    .c({\u2_Display/n3083 ,\u2_Display/n3083 }),
    .d({\u2_Display/n3053 ,\u2_Display/n3051 }),
    .f({\u2_Display/n3088 ,\u2_Display/n3086 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2475|_al_u2477  (
    .b({\u2_Display/n4243 [0],\u2_Display/n4243 [2]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4240 ,\u2_Display/n4238 }),
    .f({\u2_Display/n4275 ,\u2_Display/n4273 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2478|_al_u2479  (
    .b({\u2_Display/n4243 [3],\u2_Display/n4243 [4]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4237 ,\u2_Display/n4236 }),
    .f({\u2_Display/n4272 ,\u2_Display/n4271 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2480|_al_u2481  (
    .b({\u2_Display/n4243 [5],\u2_Display/n4243 [6]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4235 ,\u2_Display/n4234 }),
    .f({\u2_Display/n4270 ,\u2_Display/n4269 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2482|_al_u2488  (
    .b({\u2_Display/n4243 [7],\u2_Display/n4243 [13]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4233 ,\u2_Display/n4227 }),
    .f({\u2_Display/n4268 ,\u2_Display/n4262 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2483|_al_u2485  (
    .b({\u2_Display/n4243 [8],\u2_Display/n4243 [10]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4232 ,\u2_Display/n4230 }),
    .f({\u2_Display/n4267 ,\u2_Display/n4265 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2486|_al_u2492  (
    .b({\u2_Display/n4243 [11],\u2_Display/n4243 [17]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4229 ,\u2_Display/n4223 }),
    .f({\u2_Display/n4264 ,\u2_Display/n4258 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2487|_al_u2489  (
    .b({\u2_Display/n4243 [12],\u2_Display/n4243 [14]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4228 ,\u2_Display/n4226 }),
    .f({\u2_Display/n4263 ,\u2_Display/n4261 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2490|_al_u2496  (
    .b({\u2_Display/n4243 [15],\u2_Display/n4243 [21]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4225 ,\u2_Display/n4219 }),
    .f({\u2_Display/n4260 ,\u2_Display/n4254 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2491|_al_u2493  (
    .b({\u2_Display/n4243 [16],\u2_Display/n4243 [18]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4224 ,\u2_Display/n4222 }),
    .f({\u2_Display/n4259 ,\u2_Display/n4257 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2494|_al_u2500  (
    .b({\u2_Display/n4243 [19],\u2_Display/n4243 [25]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4221 ,\u2_Display/n4215 }),
    .f({\u2_Display/n4256 ,\u2_Display/n4250 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2495|_al_u2497  (
    .b({\u2_Display/n4243 [20],\u2_Display/n4243 [22]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4220 ,\u2_Display/n4218 }),
    .f({\u2_Display/n4255 ,\u2_Display/n4253 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2498|_al_u2504  (
    .b({\u2_Display/n4243 [23],\u2_Display/n4243 [29]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4217 ,\u2_Display/n4211 }),
    .f({\u2_Display/n4252 ,\u2_Display/n4246 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2499|_al_u2501  (
    .b({\u2_Display/n4243 [24],\u2_Display/n4243 [26]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4216 ,\u2_Display/n4214 }),
    .f({\u2_Display/n4251 ,\u2_Display/n4249 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2502|_al_u2506  (
    .b({\u2_Display/n4243 [27],\u2_Display/n4243 [31]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4213 ,\u2_Display/n4209 }),
    .f({\u2_Display/n4248 ,\u2_Display/n4244 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2503|_al_u2505  (
    .b({\u2_Display/n4243 [28],\u2_Display/n4243 [30]}),
    .c({\u2_Display/n4241 ,\u2_Display/n4241 }),
    .d({\u2_Display/n4212 ,\u2_Display/n4210 }),
    .f({\u2_Display/n4247 ,\u2_Display/n4245 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2507|_al_u2509  (
    .b({\u2_Display/n5366 [0],\u2_Display/n5366 [2]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5363 ,\u2_Display/n5361 }),
    .f({\u2_Display/n5398 ,\u2_Display/n5396 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2508|_al_u2511  (
    .b({\u2_Display/n5366 [1],\u2_Display/n5366 [4]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5362 ,\u2_Display/n5359 }),
    .f({\u2_Display/n5397 ,\u2_Display/n5394 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2510|_al_u2513  (
    .b({\u2_Display/n5366 [3],\u2_Display/n5366 [6]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5360 ,\u2_Display/n5357 }),
    .f({\u2_Display/n5395 ,\u2_Display/n5392 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2512|_al_u2515  (
    .b({\u2_Display/n5366 [5],\u2_Display/n5366 [8]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5358 ,\u2_Display/n5355 }),
    .f({\u2_Display/n5393 ,\u2_Display/n5390 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2514|_al_u2517  (
    .b({\u2_Display/n5366 [7],\u2_Display/n5366 [10]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5356 ,\u2_Display/n5353 }),
    .f({\u2_Display/n5391 ,\u2_Display/n5388 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2516|_al_u2520  (
    .b({\u2_Display/n5366 [9],\u2_Display/n5366 [13]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5354 ,\u2_Display/n5350 }),
    .f({\u2_Display/n5389 ,\u2_Display/n5385 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2518|_al_u2524  (
    .b({\u2_Display/n5366 [11],\u2_Display/n5366 [17]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5352 ,\u2_Display/n5346 }),
    .f({\u2_Display/n5387 ,\u2_Display/n5381 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2519|_al_u2521  (
    .b({\u2_Display/n5366 [12],\u2_Display/n5366 [14]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5351 ,\u2_Display/n5349 }),
    .f({\u2_Display/n5386 ,\u2_Display/n5384 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2522|_al_u2528  (
    .b({\u2_Display/n5366 [15],\u2_Display/n5366 [21]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5348 ,\u2_Display/n5342 }),
    .f({\u2_Display/n5383 ,\u2_Display/n5377 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2523|_al_u2525  (
    .b({\u2_Display/n5366 [16],\u2_Display/n5366 [18]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5347 ,\u2_Display/n5345 }),
    .f({\u2_Display/n5382 ,\u2_Display/n5380 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2526|_al_u2532  (
    .b({\u2_Display/n5366 [19],\u2_Display/n5366 [25]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5344 ,\u2_Display/n5338 }),
    .f({\u2_Display/n5379 ,\u2_Display/n5373 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2527|_al_u2529  (
    .b({\u2_Display/n5366 [20],\u2_Display/n5366 [22]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5343 ,\u2_Display/n5341 }),
    .f({\u2_Display/n5378 ,\u2_Display/n5376 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2530|_al_u2535  (
    .b({\u2_Display/n5366 [23],\u2_Display/n5366 [28]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5340 ,\u2_Display/n5335 }),
    .f({\u2_Display/n5375 ,\u2_Display/n5370 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2531|_al_u2533  (
    .b({\u2_Display/n5366 [24],\u2_Display/n5366 [26]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5339 ,\u2_Display/n5337 }),
    .f({\u2_Display/n5374 ,\u2_Display/n5372 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2534|_al_u2537  (
    .b({\u2_Display/n5366 [27],\u2_Display/n5366 [30]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5336 ,\u2_Display/n5333 }),
    .f({\u2_Display/n5371 ,\u2_Display/n5368 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2536|_al_u2538  (
    .b({\u2_Display/n5366 [29],\u2_Display/n5366 [31]}),
    .c({\u2_Display/n5364 ,\u2_Display/n5364 }),
    .d({\u2_Display/n5334 ,\u2_Display/n5332 }),
    .f({\u2_Display/n5369 ,\u2_Display/n5367 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2539|_al_u2541  (
    .b({\u2_Display/n874 [0],\u2_Display/n874 [2]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n871 ,\u2_Display/n869 }),
    .f({\u2_Display/n906 ,\u2_Display/n904 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u2540 (
    .b({open_n18732,\u2_Display/n874 [1]}),
    .c({open_n18733,\u2_Display/n872 }),
    .d({open_n18736,\u2_Display/n870 }),
    .f({open_n18754,\u2_Display/n905 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2542|_al_u2543  (
    .b({\u2_Display/n874 [3],\u2_Display/n874 [4]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n868 ,\u2_Display/n867 }),
    .f({\u2_Display/n903 ,\u2_Display/n902 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2544|_al_u2545  (
    .b({\u2_Display/n874 [5],\u2_Display/n874 [6]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n866 ,\u2_Display/n865 }),
    .f({\u2_Display/n901 ,\u2_Display/n900 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2546|_al_u2547  (
    .b({\u2_Display/n874 [7],\u2_Display/n874 [8]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n864 ,\u2_Display/n863 }),
    .f({\u2_Display/n899 ,\u2_Display/n898 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2548|_al_u2549  (
    .b({\u2_Display/n874 [9],\u2_Display/n874 [10]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n862 ,\u2_Display/n861 }),
    .f({\u2_Display/n897 ,\u2_Display/n896 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2550|_al_u2553  (
    .b({\u2_Display/n874 [11],\u2_Display/n874 [14]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n860 ,\u2_Display/n857 }),
    .f({\u2_Display/n895 ,\u2_Display/n892 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2551|_al_u2552  (
    .b({\u2_Display/n874 [12],\u2_Display/n874 [13]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n859 ,\u2_Display/n858 }),
    .f({\u2_Display/n894 ,\u2_Display/n893 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2554|_al_u2555  (
    .b({\u2_Display/n874 [15],\u2_Display/n874 [16]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n856 ,\u2_Display/n855 }),
    .f({\u2_Display/n891 ,\u2_Display/n890 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2556|_al_u2557  (
    .b({\u2_Display/n874 [17],\u2_Display/n874 [18]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n854 ,\u2_Display/n853 }),
    .f({\u2_Display/n889 ,\u2_Display/n888 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2558|_al_u2559  (
    .b({\u2_Display/n874 [19],\u2_Display/n874 [20]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n852 ,\u2_Display/n851 }),
    .f({\u2_Display/n887 ,\u2_Display/n886 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2560|_al_u2561  (
    .b({\u2_Display/n874 [21],\u2_Display/n874 [22]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n850 ,\u2_Display/n849 }),
    .f({\u2_Display/n885 ,\u2_Display/n884 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2562|_al_u2565  (
    .b({\u2_Display/n874 [23],\u2_Display/n874 [26]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n848 ,\u2_Display/n845 }),
    .f({\u2_Display/n883 ,\u2_Display/n880 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u2563 (
    .b({open_n19048,\u2_Display/n874 [24]}),
    .c({open_n19049,\u2_Display/n872 }),
    .d({open_n19052,\u2_Display/n847 }),
    .f({open_n19070,\u2_Display/n882 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2564|_al_u2567  (
    .b({\u2_Display/n874 [25],\u2_Display/n874 [28]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n846 ,\u2_Display/n843 }),
    .f({\u2_Display/n881 ,\u2_Display/n878 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2566|_al_u2569  (
    .b({\u2_Display/n874 [27],\u2_Display/n874 [30]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n844 ,\u2_Display/n841 }),
    .f({\u2_Display/n879 ,\u2_Display/n876 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2568|_al_u2570  (
    .b({\u2_Display/n874 [29],\u2_Display/n874 [31]}),
    .c({\u2_Display/n872 ,\u2_Display/n872 }),
    .d({\u2_Display/n842 ,\u2_Display/n840 }),
    .f({\u2_Display/n877 ,\u2_Display/n875 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2571|_al_u2573  (
    .b({\u2_Display/n1997 [0],\u2_Display/n1997 [2]}),
    .c({\u2_Display/n1995 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1994 ,\u2_Display/n1992 }),
    .f({\u2_Display/n2029 ,\u2_Display/n2027 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2574|_al_u2577  (
    .b({\u2_Display/n1997 [3],\u2_Display/n1997 [6]}),
    .c({\u2_Display/n1995 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1991 ,\u2_Display/n1988 }),
    .f({\u2_Display/n2026 ,\u2_Display/n2023 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2575|_al_u2576  (
    .b({\u2_Display/n1997 [4],\u2_Display/n1997 [5]}),
    .c({\u2_Display/n1995 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1990 ,\u2_Display/n1989 }),
    .f({\u2_Display/n2025 ,\u2_Display/n2024 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2578|_al_u2583  (
    .b({\u2_Display/n1997 [7],\u2_Display/n1997 [12]}),
    .c({\u2_Display/n1995 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1987 ,\u2_Display/n1982 }),
    .f({\u2_Display/n2022 ,\u2_Display/n2017 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2579|_al_u2581  (
    .b({\u2_Display/n1997 [8],\u2_Display/n1997 [10]}),
    .c({\u2_Display/n1995 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1986 ,\u2_Display/n1984 }),
    .f({\u2_Display/n2021 ,\u2_Display/n2019 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2582|_al_u2585  (
    .b({\u2_Display/n1997 [11],\u2_Display/n1997 [14]}),
    .c({\u2_Display/n1995 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1983 ,\u2_Display/n1980 }),
    .f({\u2_Display/n2018 ,\u2_Display/n2015 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2584|_al_u2588  (
    .b({\u2_Display/n1997 [13],\u2_Display/n1997 [17]}),
    .c({\u2_Display/n1995 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1981 ,\u2_Display/n1977 }),
    .f({\u2_Display/n2016 ,\u2_Display/n2012 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2586|_al_u2591  (
    .b({\u2_Display/n1997 [15],\u2_Display/n1997 [20]}),
    .c({\u2_Display/n1995 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1979 ,\u2_Display/n1974 }),
    .f({\u2_Display/n2014 ,\u2_Display/n2009 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2587|_al_u2589  (
    .b({\u2_Display/n1997 [16],\u2_Display/n1997 [18]}),
    .c({\u2_Display/n1995 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1978 ,\u2_Display/n1976 }),
    .f({\u2_Display/n2013 ,\u2_Display/n2011 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2590|_al_u2593  (
    .b({\u2_Display/n1997 [19],\u2_Display/n1997 [22]}),
    .c({\u2_Display/n1995 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1975 ,\u2_Display/n1972 }),
    .f({\u2_Display/n2010 ,\u2_Display/n2007 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2592|_al_u2596  (
    .b({\u2_Display/n1997 [21],\u2_Display/n1997 [25]}),
    .c({\u2_Display/n1995 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1973 ,\u2_Display/n1969 }),
    .f({\u2_Display/n2008 ,\u2_Display/n2004 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2594|_al_u2601  (
    .b({\u2_Display/n1997 [23],\u2_Display/n1997 [30]}),
    .c({\u2_Display/n1995 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1971 ,\u2_Display/n1964 }),
    .f({\u2_Display/n2006 ,\u2_Display/n1999 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2595|_al_u2597  (
    .b({\u2_Display/n1997 [24],\u2_Display/n1997 [26]}),
    .c({\u2_Display/n1995 ,\u2_Display/n1995 }),
    .d({\u2_Display/n1970 ,\u2_Display/n1968 }),
    .f({\u2_Display/n2005 ,\u2_Display/n2003 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2598|_al_u2733  (
    .b({\u2_Display/n1997 [27],\u2_Display/n2032 [2]}),
    .c({\u2_Display/n1995 ,\u2_Display/n2030 }),
    .d({\u2_Display/n1967 ,\u2_Display/n2027 }),
    .f({\u2_Display/n2002 ,\u2_Display/n2062 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2599|_al_u2732  (
    .b({\u2_Display/n1997 [28],\u2_Display/n2032 [1]}),
    .c({\u2_Display/n1995 ,\u2_Display/n2030 }),
    .d({\u2_Display/n1966 ,\u2_Display/n2028 }),
    .f({\u2_Display/n2001 ,\u2_Display/n2063 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2600|_al_u2731  (
    .b({\u2_Display/n1997 [29],\u2_Display/n2032 [0]}),
    .c({\u2_Display/n1995 ,\u2_Display/n2030 }),
    .d({\u2_Display/n1965 ,\u2_Display/n2029 }),
    .f({\u2_Display/n2000 ,\u2_Display/n2064 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2602|_al_u2740  (
    .b({\u2_Display/n1997 [31],\u2_Display/n2032 [9]}),
    .c({\u2_Display/n1995 ,\u2_Display/n2030 }),
    .d({\u2_Display/n1963 ,\u2_Display/n2020 }),
    .f({\u2_Display/n1998 ,\u2_Display/n2055 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2603|_al_u2605  (
    .b({\u2_Display/n3120 [0],\u2_Display/n3120 [2]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3117 ,\u2_Display/n3115 }),
    .f({\u2_Display/n3152 ,\u2_Display/n3150 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2604|_al_u2607  (
    .b({\u2_Display/n3120 [1],\u2_Display/n3120 [4]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3116 ,\u2_Display/n3113 }),
    .f({\u2_Display/n3151 ,\u2_Display/n3148 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2606|_al_u2609  (
    .b({\u2_Display/n3120 [3],\u2_Display/n3120 [6]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3114 ,\u2_Display/n3111 }),
    .f({\u2_Display/n3149 ,\u2_Display/n3146 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2608|_al_u2611  (
    .b({\u2_Display/n3120 [5],\u2_Display/n3120 [8]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3112 ,\u2_Display/n3109 }),
    .f({\u2_Display/n3147 ,\u2_Display/n3144 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2610|_al_u2613  (
    .b({\u2_Display/n3120 [7],\u2_Display/n3120 [10]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3110 ,\u2_Display/n3107 }),
    .f({\u2_Display/n3145 ,\u2_Display/n3142 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2612|_al_u2615  (
    .b({\u2_Display/n3120 [9],\u2_Display/n3120 [12]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3108 ,\u2_Display/n3105 }),
    .f({\u2_Display/n3143 ,\u2_Display/n3140 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2614|_al_u2617  (
    .b({\u2_Display/n3120 [11],\u2_Display/n3120 [14]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3106 ,\u2_Display/n3103 }),
    .f({\u2_Display/n3141 ,\u2_Display/n3138 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2616|_al_u2619  (
    .b({\u2_Display/n3120 [13],\u2_Display/n3120 [16]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3104 ,\u2_Display/n3101 }),
    .f({\u2_Display/n3139 ,\u2_Display/n3136 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2618|_al_u2621  (
    .b({\u2_Display/n3120 [15],\u2_Display/n3120 [18]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3102 ,\u2_Display/n3099 }),
    .f({\u2_Display/n3137 ,\u2_Display/n3134 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2620|_al_u2623  (
    .b({\u2_Display/n3120 [17],\u2_Display/n3120 [20]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3100 ,\u2_Display/n3097 }),
    .f({\u2_Display/n3135 ,\u2_Display/n3132 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2622|_al_u2625  (
    .b({\u2_Display/n3120 [19],\u2_Display/n3120 [22]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3098 ,\u2_Display/n3095 }),
    .f({\u2_Display/n3133 ,\u2_Display/n3130 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2624|_al_u2627  (
    .b({\u2_Display/n3120 [21],\u2_Display/n3120 [24]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3096 ,\u2_Display/n3093 }),
    .f({\u2_Display/n3131 ,\u2_Display/n3128 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2626|_al_u2629  (
    .b({\u2_Display/n3120 [23],\u2_Display/n3120 [26]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3094 ,\u2_Display/n3091 }),
    .f({\u2_Display/n3129 ,\u2_Display/n3126 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2628|_al_u2763  (
    .b({\u2_Display/n3118 ,\u2_Display/n3155 [0]}),
    .c({\u2_Display/n3120 [25],\u2_Display/n3153 }),
    .d({\u2_Display/n3092 ,\u2_Display/n3152 }),
    .f({\u2_Display/n3127 ,\u2_Display/n3187 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2630|_al_u2633  (
    .b({\u2_Display/n3120 [27],\u2_Display/n3120 [30]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3090 ,\u2_Display/n3087 }),
    .f({\u2_Display/n3125 ,\u2_Display/n3122 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2631|_al_u2632  (
    .b({\u2_Display/n3120 [28],\u2_Display/n3120 [29]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3118 }),
    .d({\u2_Display/n3089 ,\u2_Display/n3088 }),
    .f({\u2_Display/n3124 ,\u2_Display/n3123 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2634|_al_u2772  (
    .b({\u2_Display/n3120 [31],\u2_Display/n3155 [9]}),
    .c({\u2_Display/n3118 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3086 ,\u2_Display/n3143 }),
    .f({\u2_Display/n3121 ,\u2_Display/n3178 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2635|_al_u2637  (
    .b({\u2_Display/n4278 [0],\u2_Display/n4278 [2]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4275 ,\u2_Display/n4273 }),
    .f({\u2_Display/n4310 ,\u2_Display/n4308 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2636|_al_u2640  (
    .b({\u2_Display/n4278 [1],\u2_Display/n4278 [5]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4274 ,\u2_Display/n4270 }),
    .f({\u2_Display/n4309 ,\u2_Display/n4305 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2638|_al_u2644  (
    .b({\u2_Display/n4278 [3],\u2_Display/n4278 [9]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4272 ,\u2_Display/n4266 }),
    .f({\u2_Display/n4307 ,\u2_Display/n4301 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2639|_al_u2641  (
    .b({\u2_Display/n4278 [4],\u2_Display/n4278 [6]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4271 ,\u2_Display/n4269 }),
    .f({\u2_Display/n4306 ,\u2_Display/n4304 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2642|_al_u2647  (
    .b({\u2_Display/n4278 [7],\u2_Display/n4278 [12]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4268 ,\u2_Display/n4263 }),
    .f({\u2_Display/n4303 ,\u2_Display/n4298 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2643|_al_u2645  (
    .b({\u2_Display/n4278 [8],\u2_Display/n4278 [10]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4267 ,\u2_Display/n4265 }),
    .f({\u2_Display/n4302 ,\u2_Display/n4300 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2646|_al_u2649  (
    .b({\u2_Display/n4278 [11],\u2_Display/n4278 [14]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4264 ,\u2_Display/n4261 }),
    .f({\u2_Display/n4299 ,\u2_Display/n4296 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2648|_al_u2651  (
    .b({\u2_Display/n4278 [13],\u2_Display/n4278 [16]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4262 ,\u2_Display/n4259 }),
    .f({\u2_Display/n4297 ,\u2_Display/n4294 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2650|_al_u2653  (
    .b({\u2_Display/n4278 [15],\u2_Display/n4278 [18]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4260 ,\u2_Display/n4257 }),
    .f({\u2_Display/n4295 ,\u2_Display/n4292 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2652|_al_u2655  (
    .b({\u2_Display/n4278 [17],\u2_Display/n4278 [20]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4258 ,\u2_Display/n4255 }),
    .f({\u2_Display/n4293 ,\u2_Display/n4290 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2654|_al_u2657  (
    .b({\u2_Display/n4278 [19],\u2_Display/n4278 [22]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4256 ,\u2_Display/n4253 }),
    .f({\u2_Display/n4291 ,\u2_Display/n4288 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2656|_al_u2659  (
    .b({\u2_Display/n4278 [21],\u2_Display/n4278 [24]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4254 ,\u2_Display/n4251 }),
    .f({\u2_Display/n4289 ,\u2_Display/n4286 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2658|_al_u2661  (
    .b({\u2_Display/n4278 [23],\u2_Display/n4278 [26]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4252 ,\u2_Display/n4249 }),
    .f({\u2_Display/n4287 ,\u2_Display/n4284 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2660|_al_u2664  (
    .b({\u2_Display/n4278 [25],\u2_Display/n4278 [29]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4250 ,\u2_Display/n4246 }),
    .f({\u2_Display/n4285 ,\u2_Display/n4281 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2662|_al_u2666  (
    .b({\u2_Display/n4278 [27],\u2_Display/n4278 [31]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4248 ,\u2_Display/n4244 }),
    .f({\u2_Display/n4283 ,\u2_Display/n4279 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2663|_al_u2665  (
    .b({\u2_Display/n4278 [28],\u2_Display/n4278 [30]}),
    .c({\u2_Display/n4276 ,\u2_Display/n4276 }),
    .d({\u2_Display/n4247 ,\u2_Display/n4245 }),
    .f({\u2_Display/n4282 ,\u2_Display/n4280 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2667|_al_u2672  (
    .b({\u2_Display/n5401 [0],\u2_Display/n5401 [5]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5398 ,\u2_Display/n5393 }),
    .f({\u2_Display/n5433 ,\u2_Display/n5428 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2668|_al_u2669  (
    .b({\u2_Display/n5401 [1],\u2_Display/n5401 [2]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5397 ,\u2_Display/n5396 }),
    .f({\u2_Display/n5432 ,\u2_Display/n5431 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2670|_al_u2676  (
    .b({\u2_Display/n5401 [3],\u2_Display/n5401 [9]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5395 ,\u2_Display/n5389 }),
    .f({\u2_Display/n5430 ,\u2_Display/n5424 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2671|_al_u2673  (
    .b({\u2_Display/n5401 [4],\u2_Display/n5401 [6]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5394 ,\u2_Display/n5392 }),
    .f({\u2_Display/n5429 ,\u2_Display/n5427 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2674|_al_u2679  (
    .b({\u2_Display/n5401 [7],\u2_Display/n5401 [12]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5391 ,\u2_Display/n5386 }),
    .f({\u2_Display/n5426 ,\u2_Display/n5421 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2675|_al_u2677  (
    .b({\u2_Display/n5401 [8],\u2_Display/n5401 [10]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5390 ,\u2_Display/n5388 }),
    .f({\u2_Display/n5425 ,\u2_Display/n5423 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2678|_al_u2681  (
    .b({\u2_Display/n5401 [11],\u2_Display/n5401 [14]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5387 ,\u2_Display/n5384 }),
    .f({\u2_Display/n5422 ,\u2_Display/n5419 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2680|_al_u2684  (
    .b({\u2_Display/n5401 [13],\u2_Display/n5401 [17]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5385 ,\u2_Display/n5381 }),
    .f({\u2_Display/n5420 ,\u2_Display/n5416 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2682|_al_u2688  (
    .b({\u2_Display/n5401 [15],\u2_Display/n5401 [21]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5383 ,\u2_Display/n5377 }),
    .f({\u2_Display/n5418 ,\u2_Display/n5412 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2683|_al_u2685  (
    .b({\u2_Display/n5401 [16],\u2_Display/n5401 [18]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5382 ,\u2_Display/n5380 }),
    .f({\u2_Display/n5417 ,\u2_Display/n5415 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2686|_al_u2691  (
    .b({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .c({\u2_Display/n5401 [19],\u2_Display/n5401 [24]}),
    .d({\u2_Display/n5379 ,\u2_Display/n5374 }),
    .f({\u2_Display/n5414 ,\u2_Display/n5409 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2687|_al_u2689  (
    .b({\u2_Display/n5401 [20],\u2_Display/n5401 [22]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5378 ,\u2_Display/n5376 }),
    .f({\u2_Display/n5413 ,\u2_Display/n5411 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTF1("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTG0("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTG1("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    .INIT_LUTF0(16'b1111101001010000),
    .INIT_LUTF1(16'b1111101001010000),
    .INIT_LUTG0(16'b1111101001010000),
    .INIT_LUTG1(16'b1111101001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2690|_al_u2693  (
    .a({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .c({\u2_Display/n5401 [23],\u2_Display/n5401 [26]}),
    .d({\u2_Display/n5375 ,\u2_Display/n5372 }),
    .f({\u2_Display/n5410 ,\u2_Display/n5407 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2692|_al_u2695  (
    .b({\u2_Display/n5401 [25],\u2_Display/n5401 [28]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5373 ,\u2_Display/n5370 }),
    .f({\u2_Display/n5408 ,\u2_Display/n5405 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2694|_al_u2697  (
    .b({\u2_Display/n5401 [27],\u2_Display/n5401 [30]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5371 ,\u2_Display/n5368 }),
    .f({\u2_Display/n5406 ,\u2_Display/n5403 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2696|_al_u2698  (
    .b({\u2_Display/n5401 [29],\u2_Display/n5401 [31]}),
    .c({\u2_Display/n5399 ,\u2_Display/n5399 }),
    .d({\u2_Display/n5369 ,\u2_Display/n5367 }),
    .f({\u2_Display/n5404 ,\u2_Display/n5402 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2699|_al_u2701  (
    .b({\u2_Display/n909 [0],\u2_Display/n909 [2]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n906 ,\u2_Display/n904 }),
    .f({\u2_Display/n941 ,\u2_Display/n939 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2700|_al_u2704  (
    .b({\u2_Display/n909 [1],\u2_Display/n909 [5]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n905 ,\u2_Display/n901 }),
    .f({\u2_Display/n940 ,\u2_Display/n936 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2702|_al_u2707  (
    .b({\u2_Display/n909 [3],\u2_Display/n909 [8]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n903 ,\u2_Display/n898 }),
    .f({\u2_Display/n938 ,\u2_Display/n933 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2703|_al_u2705  (
    .b({\u2_Display/n909 [4],\u2_Display/n909 [6]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n902 ,\u2_Display/n900 }),
    .f({\u2_Display/n937 ,\u2_Display/n935 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2706|_al_u2709  (
    .b({\u2_Display/n909 [7],\u2_Display/n909 [10]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n899 ,\u2_Display/n896 }),
    .f({\u2_Display/n934 ,\u2_Display/n931 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2708|_al_u2711  (
    .b({\u2_Display/n909 [9],\u2_Display/n909 [12]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n897 ,\u2_Display/n894 }),
    .f({\u2_Display/n932 ,\u2_Display/n929 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2710|_al_u2713  (
    .b({\u2_Display/n909 [11],\u2_Display/n909 [14]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n895 ,\u2_Display/n892 }),
    .f({\u2_Display/n930 ,\u2_Display/n927 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2712|_al_u2715  (
    .b({\u2_Display/n909 [13],\u2_Display/n909 [16]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n893 ,\u2_Display/n890 }),
    .f({\u2_Display/n928 ,\u2_Display/n925 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2714|_al_u2717  (
    .b({\u2_Display/n909 [15],\u2_Display/n909 [18]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n891 ,\u2_Display/n888 }),
    .f({\u2_Display/n926 ,\u2_Display/n923 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2716|_al_u2720  (
    .b({\u2_Display/n909 [17],\u2_Display/n909 [21]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n889 ,\u2_Display/n885 }),
    .f({\u2_Display/n924 ,\u2_Display/n920 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2718|_al_u2724  (
    .b({\u2_Display/n909 [19],\u2_Display/n909 [25]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n887 ,\u2_Display/n881 }),
    .f({\u2_Display/n922 ,\u2_Display/n916 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2719|_al_u2721  (
    .b({\u2_Display/n909 [20],\u2_Display/n909 [22]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n886 ,\u2_Display/n884 }),
    .f({\u2_Display/n921 ,\u2_Display/n919 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2722|_al_u2727  (
    .b({\u2_Display/n909 [23],\u2_Display/n909 [28]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n883 ,\u2_Display/n878 }),
    .f({\u2_Display/n918 ,\u2_Display/n913 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2723|_al_u2725  (
    .b({\u2_Display/n909 [24],\u2_Display/n909 [26]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n882 ,\u2_Display/n880 }),
    .f({\u2_Display/n917 ,\u2_Display/n915 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2726|_al_u2729  (
    .b({\u2_Display/n909 [27],\u2_Display/n909 [30]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n879 ,\u2_Display/n876 }),
    .f({\u2_Display/n914 ,\u2_Display/n911 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2728|_al_u2730  (
    .b({\u2_Display/n909 [29],\u2_Display/n909 [31]}),
    .c({\u2_Display/n907 ,\u2_Display/n907 }),
    .d({\u2_Display/n877 ,\u2_Display/n875 }),
    .f({\u2_Display/n912 ,\u2_Display/n910 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2734|_al_u2737  (
    .b({\u2_Display/n2032 [3],\u2_Display/n2032 [6]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2030 }),
    .d({\u2_Display/n2026 ,\u2_Display/n2023 }),
    .f({\u2_Display/n2061 ,\u2_Display/n2058 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2735|_al_u2736  (
    .b({\u2_Display/n2032 [4],\u2_Display/n2032 [5]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2030 }),
    .d({\u2_Display/n2025 ,\u2_Display/n2024 }),
    .f({\u2_Display/n2060 ,\u2_Display/n2059 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2738|_al_u2744  (
    .b({\u2_Display/n2032 [7],\u2_Display/n2032 [13]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2030 }),
    .d({\u2_Display/n2022 ,\u2_Display/n2016 }),
    .f({\u2_Display/n2057 ,\u2_Display/n2051 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2739|_al_u2741  (
    .b({\u2_Display/n2032 [8],\u2_Display/n2032 [10]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2030 }),
    .d({\u2_Display/n2021 ,\u2_Display/n2019 }),
    .f({\u2_Display/n2056 ,\u2_Display/n2054 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2742|_al_u2748  (
    .b({\u2_Display/n2032 [11],\u2_Display/n2032 [17]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2030 }),
    .d({\u2_Display/n2018 ,\u2_Display/n2012 }),
    .f({\u2_Display/n2053 ,\u2_Display/n2047 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2743|_al_u2745  (
    .b({\u2_Display/n2032 [12],\u2_Display/n2032 [14]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2030 }),
    .d({\u2_Display/n2017 ,\u2_Display/n2015 }),
    .f({\u2_Display/n2052 ,\u2_Display/n2050 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2746|_al_u2751  (
    .b({\u2_Display/n2032 [15],\u2_Display/n2032 [20]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2030 }),
    .d({\u2_Display/n2014 ,\u2_Display/n2009 }),
    .f({\u2_Display/n2049 ,\u2_Display/n2044 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2747|_al_u2749  (
    .b({\u2_Display/n2032 [16],\u2_Display/n2032 [18]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2030 }),
    .d({\u2_Display/n2013 ,\u2_Display/n2011 }),
    .f({\u2_Display/n2048 ,\u2_Display/n2046 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2750|_al_u2753  (
    .b({\u2_Display/n2032 [19],\u2_Display/n2032 [22]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2030 }),
    .d({\u2_Display/n2010 ,\u2_Display/n2007 }),
    .f({\u2_Display/n2045 ,\u2_Display/n2042 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2752|_al_u2755  (
    .b({\u2_Display/n2032 [21],\u2_Display/n2032 [24]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2030 }),
    .d({\u2_Display/n2008 ,\u2_Display/n2005 }),
    .f({\u2_Display/n2043 ,\u2_Display/n2040 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2754|_al_u2757  (
    .b({\u2_Display/n2032 [23],\u2_Display/n2032 [26]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2030 }),
    .d({\u2_Display/n2006 ,\u2_Display/n2003 }),
    .f({\u2_Display/n2041 ,\u2_Display/n2038 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2756|_al_u2761  (
    .b({\u2_Display/n2032 [25],\u2_Display/n2032 [30]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2030 }),
    .d({\u2_Display/n2004 ,\u2_Display/n1999 }),
    .f({\u2_Display/n2039 ,\u2_Display/n2034 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2758|_al_u2893  (
    .b({\u2_Display/n2032 [27],\u2_Display/n2067 [2]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2002 ,\u2_Display/n2062 }),
    .f({\u2_Display/n2037 ,\u2_Display/n2097 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2759|_al_u2892  (
    .b({\u2_Display/n2032 [28],\u2_Display/n2067 [1]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2001 ,\u2_Display/n2063 }),
    .f({\u2_Display/n2036 ,\u2_Display/n2098 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2760|_al_u2891  (
    .b({\u2_Display/n2032 [29],\u2_Display/n2067 [0]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2000 ,\u2_Display/n2064 }),
    .f({\u2_Display/n2035 ,\u2_Display/n2099 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2762|_al_u2899  (
    .b({\u2_Display/n2032 [31],\u2_Display/n2067 [8]}),
    .c({\u2_Display/n2030 ,\u2_Display/n2065 }),
    .d({\u2_Display/n1998 ,\u2_Display/n2056 }),
    .f({\u2_Display/n2033 ,\u2_Display/n2091 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2764|_al_u2765  (
    .b({\u2_Display/n3155 [1],\u2_Display/n3155 [2]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3151 ,\u2_Display/n3150 }),
    .f({\u2_Display/n3186 ,\u2_Display/n3185 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2766|_al_u2769  (
    .b({\u2_Display/n3155 [3],\u2_Display/n3155 [6]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3149 ,\u2_Display/n3146 }),
    .f({\u2_Display/n3184 ,\u2_Display/n3181 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2767|_al_u2768  (
    .b({\u2_Display/n3155 [4],\u2_Display/n3155 [5]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3148 ,\u2_Display/n3147 }),
    .f({\u2_Display/n3183 ,\u2_Display/n3182 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2770|_al_u2775  (
    .b({\u2_Display/n3155 [7],\u2_Display/n3155 [12]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3145 ,\u2_Display/n3140 }),
    .f({\u2_Display/n3180 ,\u2_Display/n3175 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2771|_al_u2773  (
    .b({\u2_Display/n3155 [8],\u2_Display/n3155 [10]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3144 ,\u2_Display/n3142 }),
    .f({\u2_Display/n3179 ,\u2_Display/n3177 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2774|_al_u2777  (
    .b({\u2_Display/n3155 [11],\u2_Display/n3155 [14]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3141 ,\u2_Display/n3138 }),
    .f({\u2_Display/n3176 ,\u2_Display/n3173 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2776|_al_u2779  (
    .b({\u2_Display/n3155 [13],\u2_Display/n3155 [16]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3139 ,\u2_Display/n3136 }),
    .f({\u2_Display/n3174 ,\u2_Display/n3171 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2778|_al_u2781  (
    .b({\u2_Display/n3155 [15],\u2_Display/n3155 [18]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3137 ,\u2_Display/n3134 }),
    .f({\u2_Display/n3172 ,\u2_Display/n3169 }));
  EG_PHY_PAD #(
    //.LOCATION("K14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u278 (
    .ipad(clk_24m),
    .di(clk_24m_pad));  // source/rtl/VGA_Demo.v(4)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2780|_al_u2783  (
    .b({\u2_Display/n3155 [17],\u2_Display/n3155 [20]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3135 ,\u2_Display/n3132 }),
    .f({\u2_Display/n3170 ,\u2_Display/n3167 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2782|_al_u2785  (
    .b({\u2_Display/n3155 [19],\u2_Display/n3155 [22]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3133 ,\u2_Display/n3130 }),
    .f({\u2_Display/n3168 ,\u2_Display/n3165 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2784|_al_u2788  (
    .b({\u2_Display/n3155 [21],\u2_Display/n3155 [25]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3131 ,\u2_Display/n3127 }),
    .f({\u2_Display/n3166 ,\u2_Display/n3162 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2786|_al_u2792  (
    .b({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .c({\u2_Display/n3155 [23],\u2_Display/n3155 [29]}),
    .d({\u2_Display/n3129 ,\u2_Display/n3123 }),
    .f({\u2_Display/n3164 ,\u2_Display/n3158 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2787|_al_u2789  (
    .b({\u2_Display/n3155 [24],\u2_Display/n3155 [26]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3128 ,\u2_Display/n3126 }),
    .f({\u2_Display/n3163 ,\u2_Display/n3161 }));
  EG_PHY_PAD #(
    //.LOCATION("P8"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u279 (
    .ipad(on_off[7]));  // source/rtl/VGA_Demo.v(6)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2790|_al_u2794  (
    .b({\u2_Display/n3155 [27],\u2_Display/n3155 [31]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3125 ,\u2_Display/n3121 }),
    .f({\u2_Display/n3160 ,\u2_Display/n3156 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2791|_al_u2793  (
    .b({\u2_Display/n3155 [28],\u2_Display/n3155 [30]}),
    .c({\u2_Display/n3153 ,\u2_Display/n3153 }),
    .d({\u2_Display/n3124 ,\u2_Display/n3122 }),
    .f({\u2_Display/n3159 ,\u2_Display/n3157 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2795|_al_u2797  (
    .b({\u2_Display/n4313 [0],\u2_Display/n4313 [2]}),
    .c({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .d({\u2_Display/n4310 ,\u2_Display/n4308 }),
    .f({\u2_Display/n4345 ,\u2_Display/n4343 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u2796 (
    .b({open_n22155,\u2_Display/n4313 [1]}),
    .c({open_n22156,\u2_Display/n4311 }),
    .d({open_n22159,\u2_Display/n4309 }),
    .f({open_n22177,\u2_Display/n4344 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2798|_al_u2799  (
    .b({\u2_Display/n4313 [3],\u2_Display/n4313 [4]}),
    .c({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .d({\u2_Display/n4307 ,\u2_Display/n4306 }),
    .f({\u2_Display/n4342 ,\u2_Display/n4341 }));
  EG_PHY_PAD #(
    //.LOCATION("N6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u280 (
    .ipad(on_off[6]));  // source/rtl/VGA_Demo.v(6)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2800|_al_u2801  (
    .b({\u2_Display/n4313 [5],\u2_Display/n4313 [6]}),
    .c({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .d({\u2_Display/n4305 ,\u2_Display/n4304 }),
    .f({\u2_Display/n4340 ,\u2_Display/n4339 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2802|_al_u2805  (
    .b({\u2_Display/n4313 [7],\u2_Display/n4313 [10]}),
    .c({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .d({\u2_Display/n4303 ,\u2_Display/n4300 }),
    .f({\u2_Display/n4338 ,\u2_Display/n4335 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2803|_al_u2804  (
    .b({\u2_Display/n4313 [8],\u2_Display/n4313 [9]}),
    .c({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .d({\u2_Display/n4302 ,\u2_Display/n4301 }),
    .f({\u2_Display/n4337 ,\u2_Display/n4336 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2806|_al_u2807  (
    .b({\u2_Display/n4313 [11],\u2_Display/n4313 [12]}),
    .c({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .d({\u2_Display/n4299 ,\u2_Display/n4298 }),
    .f({\u2_Display/n4334 ,\u2_Display/n4333 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2808|_al_u2809  (
    .b({\u2_Display/n4313 [13],\u2_Display/n4313 [14]}),
    .c({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .d({\u2_Display/n4297 ,\u2_Display/n4296 }),
    .f({\u2_Display/n4332 ,\u2_Display/n4331 }));
  EG_PHY_PAD #(
    //.LOCATION("P6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u281 (
    .ipad(on_off[5]));  // source/rtl/VGA_Demo.v(6)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2810|_al_u2811  (
    .b({\u2_Display/n4313 [15],\u2_Display/n4313 [16]}),
    .c({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .d({\u2_Display/n4295 ,\u2_Display/n4294 }),
    .f({\u2_Display/n4330 ,\u2_Display/n4329 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2812|_al_u2813  (
    .b({\u2_Display/n4313 [17],\u2_Display/n4313 [18]}),
    .c({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .d({\u2_Display/n4293 ,\u2_Display/n4292 }),
    .f({\u2_Display/n4328 ,\u2_Display/n4327 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2814|_al_u2817  (
    .b({\u2_Display/n4313 [19],\u2_Display/n4313 [22]}),
    .c({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .d({\u2_Display/n4291 ,\u2_Display/n4288 }),
    .f({\u2_Display/n4326 ,\u2_Display/n4323 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2815|_al_u2816  (
    .b({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .c({\u2_Display/n4313 [20],\u2_Display/n4313 [21]}),
    .d({\u2_Display/n4290 ,\u2_Display/n4289 }),
    .f({\u2_Display/n4325 ,\u2_Display/n4324 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    //.LUTF1("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUTG0("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    //.LUTG1("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT_LUTF0(16'b1101100011011000),
    .INIT_LUTF1(16'b1110010011100100),
    .INIT_LUTG0(16'b1101100011011000),
    .INIT_LUTG1(16'b1110010011100100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2818|_al_u2821  (
    .a({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .b({\u2_Display/n4313 [23],\u2_Display/n4284 }),
    .c({\u2_Display/n4287 ,\u2_Display/n4313 [26]}),
    .f({\u2_Display/n4322 ,\u2_Display/n4319 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2819|_al_u2820  (
    .b({\u2_Display/n4313 [24],\u2_Display/n4313 [25]}),
    .c({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .d({\u2_Display/n4286 ,\u2_Display/n4285 }),
    .f({\u2_Display/n4321 ,\u2_Display/n4320 }));
  EG_PHY_PAD #(
    //.LOCATION("M6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u282 (
    .ipad(on_off[4]),
    .di(on_off_pad[4]));  // source/rtl/VGA_Demo.v(6)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2822|_al_u2823  (
    .b({\u2_Display/n4313 [27],\u2_Display/n4313 [28]}),
    .c({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .d({\u2_Display/n4283 ,\u2_Display/n4282 }),
    .f({\u2_Display/n4318 ,\u2_Display/n4317 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2824|_al_u2825  (
    .b({\u2_Display/n4313 [29],\u2_Display/n4313 [30]}),
    .c({\u2_Display/n4311 ,\u2_Display/n4311 }),
    .d({\u2_Display/n4281 ,\u2_Display/n4280 }),
    .f({\u2_Display/n4316 ,\u2_Display/n4315 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2826|_al_u1169  (
    .b({\u2_Display/n4313 [31],open_n22602}),
    .c({\u2_Display/n4311 ,rst_n_pad}),
    .d({\u2_Display/n4279 ,_al_u1168_o}),
    .f({\u2_Display/n4314 ,\u2_Display/mux21_b0_sel_is_0_o }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2827|_al_u2832  (
    .b({\u2_Display/n5436 [0],\u2_Display/n5436 [5]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5433 ,\u2_Display/n5428 }),
    .f({\u2_Display/n5468 ,\u2_Display/n5463 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2828|_al_u2829  (
    .b({\u2_Display/n5436 [1],\u2_Display/n5436 [2]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5432 ,\u2_Display/n5431 }),
    .f({\u2_Display/n5467 ,\u2_Display/n5466 }));
  EG_PHY_PAD #(
    //.LOCATION("T6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u283 (
    .ipad(on_off[3]),
    .di(on_off_pad[3]));  // source/rtl/VGA_Demo.v(6)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2830|_al_u2835  (
    .b({\u2_Display/n5436 [3],\u2_Display/n5436 [8]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5430 ,\u2_Display/n5425 }),
    .f({\u2_Display/n5465 ,\u2_Display/n5460 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2831|_al_u2833  (
    .b({\u2_Display/n5436 [4],\u2_Display/n5436 [6]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5429 ,\u2_Display/n5427 }),
    .f({\u2_Display/n5464 ,\u2_Display/n5462 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2834|_al_u2837  (
    .b({\u2_Display/n5436 [7],\u2_Display/n5436 [10]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5426 ,\u2_Display/n5423 }),
    .f({\u2_Display/n5461 ,\u2_Display/n5458 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2836|_al_u2839  (
    .b({\u2_Display/n5436 [9],\u2_Display/n5436 [12]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5424 ,\u2_Display/n5421 }),
    .f({\u2_Display/n5459 ,\u2_Display/n5456 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2838|_al_u2841  (
    .b({\u2_Display/n5436 [11],\u2_Display/n5436 [14]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5422 ,\u2_Display/n5419 }),
    .f({\u2_Display/n5457 ,\u2_Display/n5454 }));
  EG_PHY_PAD #(
    //.LOCATION("T5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u284 (
    .ipad(on_off[2]),
    .di(on_off_pad[2]));  // source/rtl/VGA_Demo.v(6)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2840|_al_u2844  (
    .b({\u2_Display/n5436 [13],\u2_Display/n5436 [17]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5420 ,\u2_Display/n5416 }),
    .f({\u2_Display/n5455 ,\u2_Display/n5451 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2842|_al_u2847  (
    .b({\u2_Display/n5436 [15],\u2_Display/n5436 [20]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5418 ,\u2_Display/n5413 }),
    .f({\u2_Display/n5453 ,\u2_Display/n5448 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2843|_al_u2845  (
    .b({\u2_Display/n5436 [16],\u2_Display/n5436 [18]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5417 ,\u2_Display/n5415 }),
    .f({\u2_Display/n5452 ,\u2_Display/n5450 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2846|_al_u2849  (
    .b({\u2_Display/n5436 [19],\u2_Display/n5436 [22]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5414 ,\u2_Display/n5411 }),
    .f({\u2_Display/n5449 ,\u2_Display/n5446 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2848|_al_u2852  (
    .b({\u2_Display/n5436 [21],\u2_Display/n5436 [25]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5412 ,\u2_Display/n5408 }),
    .f({\u2_Display/n5447 ,\u2_Display/n5443 }));
  EG_PHY_PAD #(
    //.LOCATION("R5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u285 (
    .ipad(on_off[1]),
    .di(on_off_pad[1]));  // source/rtl/VGA_Demo.v(6)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2850|_al_u2856  (
    .b({\u2_Display/n5436 [23],\u2_Display/n5436 [29]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5410 ,\u2_Display/n5404 }),
    .f({\u2_Display/n5445 ,\u2_Display/n5439 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2851|_al_u2853  (
    .b({\u2_Display/n5436 [24],\u2_Display/n5436 [26]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5409 ,\u2_Display/n5407 }),
    .f({\u2_Display/n5444 ,\u2_Display/n5442 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2854|_al_u2858  (
    .b({\u2_Display/n5436 [27],\u2_Display/n5436 [31]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5406 ,\u2_Display/n5402 }),
    .f({\u2_Display/n5441 ,\u2_Display/n5437 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2855|_al_u2857  (
    .b({\u2_Display/n5436 [28],\u2_Display/n5436 [30]}),
    .c({\u2_Display/n5434 ,\u2_Display/n5434 }),
    .d({\u2_Display/n5405 ,\u2_Display/n5403 }),
    .f({\u2_Display/n5440 ,\u2_Display/n5438 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2859|_al_u2864  (
    .b({\u2_Display/n944 [0],\u2_Display/n944 [5]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n941 ,\u2_Display/n936 }),
    .f({\u2_Display/n976 ,\u2_Display/n971 }));
  EG_PHY_PAD #(
    //.LOCATION("T4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u286 (
    .ipad(on_off[0]),
    .di(on_off_pad[0]));  // source/rtl/VGA_Demo.v(6)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2860|_al_u2861  (
    .b({\u2_Display/n944 [1],\u2_Display/n944 [2]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n940 ,\u2_Display/n939 }),
    .f({\u2_Display/n975 ,\u2_Display/n974 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2862|_al_u2867  (
    .b({\u2_Display/n944 [3],\u2_Display/n944 [8]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n938 ,\u2_Display/n933 }),
    .f({\u2_Display/n973 ,\u2_Display/n968 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2863|_al_u2865  (
    .b({\u2_Display/n944 [4],\u2_Display/n944 [6]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n937 ,\u2_Display/n935 }),
    .f({\u2_Display/n972 ,\u2_Display/n970 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2866|_al_u2869  (
    .b({\u2_Display/n944 [7],\u2_Display/n944 [10]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n934 ,\u2_Display/n931 }),
    .f({\u2_Display/n969 ,\u2_Display/n966 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2868|_al_u2871  (
    .b({\u2_Display/n944 [9],\u2_Display/n944 [12]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n932 ,\u2_Display/n929 }),
    .f({\u2_Display/n967 ,\u2_Display/n964 }));
  EG_PHY_PAD #(
    //.LOCATION("G11"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u287 (
    .ipad(rst_n),
    .di(rst_n_pad));  // source/rtl/VGA_Demo.v(5)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2870|_al_u2873  (
    .b({\u2_Display/n944 [11],\u2_Display/n944 [14]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n930 ,\u2_Display/n927 }),
    .f({\u2_Display/n965 ,\u2_Display/n962 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2872|_al_u2875  (
    .b({\u2_Display/n944 [13],\u2_Display/n944 [16]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n928 ,\u2_Display/n925 }),
    .f({\u2_Display/n963 ,\u2_Display/n960 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2874|_al_u2877  (
    .b({\u2_Display/n944 [15],\u2_Display/n944 [18]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n926 ,\u2_Display/n923 }),
    .f({\u2_Display/n961 ,\u2_Display/n958 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2876|_al_u2880  (
    .b({\u2_Display/n944 [17],\u2_Display/n944 [21]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n924 ,\u2_Display/n920 }),
    .f({\u2_Display/n959 ,\u2_Display/n955 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2878|_al_u2884  (
    .b({\u2_Display/n944 [19],\u2_Display/n944 [25]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n922 ,\u2_Display/n916 }),
    .f({\u2_Display/n957 ,\u2_Display/n951 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2879|_al_u2881  (
    .b({\u2_Display/n944 [20],\u2_Display/n944 [22]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n921 ,\u2_Display/n919 }),
    .f({\u2_Display/n956 ,\u2_Display/n954 }));
  EG_PHY_PAD #(
    //.LOCATION("C1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u288 (
    .do({open_n23441,open_n23442,open_n23443,vga_b_pad[0]}),
    .opad(vga_b[7]));  // source/rtl/VGA_Demo.v(17)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2882|_al_u2887  (
    .b({\u2_Display/n944 [23],\u2_Display/n944 [28]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n918 ,\u2_Display/n913 }),
    .f({\u2_Display/n953 ,\u2_Display/n948 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2883|_al_u2885  (
    .b({\u2_Display/n944 [24],\u2_Display/n944 [26]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n917 ,\u2_Display/n915 }),
    .f({\u2_Display/n952 ,\u2_Display/n950 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2886|_al_u2889  (
    .b({\u2_Display/n944 [27],\u2_Display/n944 [30]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n914 ,\u2_Display/n911 }),
    .f({\u2_Display/n949 ,\u2_Display/n946 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2888|_al_u2890  (
    .b({\u2_Display/n944 [29],\u2_Display/n944 [31]}),
    .c({\u2_Display/n942 ,\u2_Display/n942 }),
    .d({\u2_Display/n912 ,\u2_Display/n910 }),
    .f({\u2_Display/n947 ,\u2_Display/n945 }));
  EG_PHY_PAD #(
    //.LOCATION("D1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u289 (
    .do({open_n23562,open_n23563,open_n23564,vga_b_pad[0]}),
    .opad(vga_b[6]));  // source/rtl/VGA_Demo.v(17)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2894|_al_u2895  (
    .b({\u2_Display/n2067 [3],\u2_Display/n2067 [4]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2061 ,\u2_Display/n2060 }),
    .f({\u2_Display/n2096 ,\u2_Display/n2095 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2896|_al_u2897  (
    .b({\u2_Display/n2067 [5],\u2_Display/n2067 [6]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2059 ,\u2_Display/n2058 }),
    .f({\u2_Display/n2094 ,\u2_Display/n2093 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2898|_al_u2901  (
    .b({\u2_Display/n2067 [7],\u2_Display/n2067 [10]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2057 ,\u2_Display/n2054 }),
    .f({\u2_Display/n2092 ,\u2_Display/n2089 }));
  EG_PHY_PAD #(
    //.LOCATION("E2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u290 (
    .do({open_n23657,open_n23658,open_n23659,vga_b_pad[0]}),
    .opad(vga_b[5]));  // source/rtl/VGA_Demo.v(17)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2900|_al_u2903  (
    .b({\u2_Display/n2067 [9],\u2_Display/n2067 [12]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2055 ,\u2_Display/n2052 }),
    .f({\u2_Display/n2090 ,\u2_Display/n2087 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2902|_al_u2905  (
    .b({\u2_Display/n2067 [11],\u2_Display/n2067 [14]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2053 ,\u2_Display/n2050 }),
    .f({\u2_Display/n2088 ,\u2_Display/n2085 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2904|_al_u2908  (
    .b({\u2_Display/n2067 [13],\u2_Display/n2067 [17]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2051 ,\u2_Display/n2047 }),
    .f({\u2_Display/n2086 ,\u2_Display/n2082 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2906|_al_u2912  (
    .b({\u2_Display/n2067 [15],\u2_Display/n2067 [21]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2049 ,\u2_Display/n2043 }),
    .f({\u2_Display/n2084 ,\u2_Display/n2078 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2907|_al_u2909  (
    .b({\u2_Display/n2067 [16],\u2_Display/n2067 [18]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2048 ,\u2_Display/n2046 }),
    .f({\u2_Display/n2083 ,\u2_Display/n2081 }));
  EG_PHY_PAD #(
    //.LOCATION("G3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u291 (
    .do({open_n23804,open_n23805,open_n23806,vga_b_pad[0]}),
    .opad(vga_b[4]));  // source/rtl/VGA_Demo.v(17)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2910|_al_u2915  (
    .b({\u2_Display/n2067 [19],\u2_Display/n2067 [24]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2045 ,\u2_Display/n2040 }),
    .f({\u2_Display/n2080 ,\u2_Display/n2075 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2911|_al_u2913  (
    .b({\u2_Display/n2067 [20],\u2_Display/n2067 [22]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2044 ,\u2_Display/n2042 }),
    .f({\u2_Display/n2079 ,\u2_Display/n2077 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2914|_al_u2917  (
    .b({\u2_Display/n2067 [23],\u2_Display/n2067 [26]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2041 ,\u2_Display/n2038 }),
    .f({\u2_Display/n2076 ,\u2_Display/n2073 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2916|_al_u2920  (
    .b({\u2_Display/n2067 [25],\u2_Display/n2067 [29]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2039 ,\u2_Display/n2035 }),
    .f({\u2_Display/n2074 ,\u2_Display/n2070 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2918|_al_u2922  (
    .b({\u2_Display/n2067 [27],\u2_Display/n2067 [31]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2037 ,\u2_Display/n2033 }),
    .f({\u2_Display/n2072 ,\u2_Display/n2068 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2919|_al_u2921  (
    .b({\u2_Display/n2067 [28],\u2_Display/n2067 [30]}),
    .c({\u2_Display/n2065 ,\u2_Display/n2065 }),
    .d({\u2_Display/n2036 ,\u2_Display/n2034 }),
    .f({\u2_Display/n2071 ,\u2_Display/n2069 }));
  EG_PHY_PAD #(
    //.LOCATION("E1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u292 (
    .do({open_n23977,open_n23978,open_n23979,vga_b_pad[0]}),
    .opad(vga_b[3]));  // source/rtl/VGA_Demo.v(17)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2923|_al_u2925  (
    .b({\u2_Display/n3190 [0],\u2_Display/n3190 [2]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3187 ,\u2_Display/n3185 }),
    .f({\u2_Display/n3222 ,\u2_Display/n3220 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2924|_al_u2927  (
    .b({\u2_Display/n3190 [1],\u2_Display/n3190 [4]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3186 ,\u2_Display/n3183 }),
    .f({\u2_Display/n3221 ,\u2_Display/n3218 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2926|_al_u2929  (
    .b({\u2_Display/n3190 [3],\u2_Display/n3190 [6]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3184 ,\u2_Display/n3181 }),
    .f({\u2_Display/n3219 ,\u2_Display/n3216 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2928|_al_u2931  (
    .b({\u2_Display/n3190 [5],\u2_Display/n3190 [8]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3182 ,\u2_Display/n3179 }),
    .f({\u2_Display/n3217 ,\u2_Display/n3214 }));
  EG_PHY_PAD #(
    //.LOCATION("F2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u293 (
    .do({open_n24098,open_n24099,open_n24100,vga_b_pad[0]}),
    .opad(vga_b[2]));  // source/rtl/VGA_Demo.v(17)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2930|_al_u2933  (
    .b({\u2_Display/n3190 [7],\u2_Display/n3190 [10]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3180 ,\u2_Display/n3177 }),
    .f({\u2_Display/n3215 ,\u2_Display/n3212 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2932|_al_u2935  (
    .b({\u2_Display/n3190 [9],\u2_Display/n3190 [12]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3178 ,\u2_Display/n3175 }),
    .f({\u2_Display/n3213 ,\u2_Display/n3210 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2934|_al_u2937  (
    .b({\u2_Display/n3190 [11],\u2_Display/n3190 [14]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3176 ,\u2_Display/n3173 }),
    .f({\u2_Display/n3211 ,\u2_Display/n3208 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2936|_al_u2939  (
    .b({\u2_Display/n3190 [13],\u2_Display/n3190 [16]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3174 ,\u2_Display/n3171 }),
    .f({\u2_Display/n3209 ,\u2_Display/n3206 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2938|_al_u2941  (
    .b({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .c({\u2_Display/n3190 [15],\u2_Display/n3190 [18]}),
    .d({\u2_Display/n3172 ,\u2_Display/n3169 }),
    .f({\u2_Display/n3207 ,\u2_Display/n3204 }));
  EG_PHY_PAD #(
    //.LOCATION("F1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u294 (
    .do({open_n24245,open_n24246,open_n24247,vga_b_pad[0]}),
    .opad(vga_b[1]));  // source/rtl/VGA_Demo.v(17)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2940|_al_u2944  (
    .b({\u2_Display/n3190 [17],\u2_Display/n3190 [21]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3170 ,\u2_Display/n3166 }),
    .f({\u2_Display/n3205 ,\u2_Display/n3201 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2942|_al_u2948  (
    .b({\u2_Display/n3190 [19],\u2_Display/n3190 [25]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3168 ,\u2_Display/n3162 }),
    .f({\u2_Display/n3203 ,\u2_Display/n3197 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2943|_al_u2945  (
    .b({\u2_Display/n3190 [20],\u2_Display/n3190 [22]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3167 ,\u2_Display/n3165 }),
    .f({\u2_Display/n3202 ,\u2_Display/n3200 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2946|_al_u3084  (
    .b({\u2_Display/n3190 [23],\u2_Display/n3225 [1]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3164 ,\u2_Display/n3221 }),
    .f({\u2_Display/n3199 ,\u2_Display/n3256 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2947|_al_u2949  (
    .b({\u2_Display/n3190 [24],\u2_Display/n3190 [26]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3163 ,\u2_Display/n3161 }),
    .f({\u2_Display/n3198 ,\u2_Display/n3196 }));
  EG_PHY_PAD #(
    //.LOCATION("G1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u295 (
    .do({open_n24392,open_n24393,open_n24394,vga_b_pad[0]}),
    .opad(vga_b[0]));  // source/rtl/VGA_Demo.v(17)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2950|_al_u2953  (
    .b({\u2_Display/n3190 [27],\u2_Display/n3190 [30]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3160 ,\u2_Display/n3157 }),
    .f({\u2_Display/n3195 ,\u2_Display/n3192 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2951|_al_u2952  (
    .b({\u2_Display/n3190 [28],\u2_Display/n3190 [29]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3188 }),
    .d({\u2_Display/n3159 ,\u2_Display/n3158 }),
    .f({\u2_Display/n3194 ,\u2_Display/n3193 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2954|_al_u3091  (
    .b({\u2_Display/n3190 [31],\u2_Display/n3225 [8]}),
    .c({\u2_Display/n3188 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3156 ,\u2_Display/n3214 }),
    .f({\u2_Display/n3191 ,\u2_Display/n3249 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2955|_al_u2960  (
    .b({\u2_Display/n4348 [0],\u2_Display/n4348 [5]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4345 ,\u2_Display/n4340 }),
    .f({\u2_Display/n4380 ,\u2_Display/n4375 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2956|_al_u2957  (
    .b({\u2_Display/n4348 [1],\u2_Display/n4348 [2]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4344 ,\u2_Display/n4343 }),
    .f({\u2_Display/n4379 ,\u2_Display/n4378 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2958|_al_u2964  (
    .b({\u2_Display/n4348 [3],\u2_Display/n4348 [9]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4342 ,\u2_Display/n4336 }),
    .f({\u2_Display/n4377 ,\u2_Display/n4371 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2959|_al_u2961  (
    .b({\u2_Display/n4348 [4],\u2_Display/n4348 [6]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4341 ,\u2_Display/n4339 }),
    .f({\u2_Display/n4376 ,\u2_Display/n4374 }));
  EG_PHY_PAD #(
    //.LOCATION("H2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u296 (
    .do({open_n24591,open_n24592,open_n24593,vga_clk_pad}),
    .opad(vga_clk));  // source/rtl/VGA_Demo.v(9)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2962|_al_u2968  (
    .b({\u2_Display/n4348 [7],\u2_Display/n4348 [13]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4338 ,\u2_Display/n4332 }),
    .f({\u2_Display/n4373 ,\u2_Display/n4367 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2963|_al_u2965  (
    .b({\u2_Display/n4348 [8],\u2_Display/n4348 [10]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4337 ,\u2_Display/n4335 }),
    .f({\u2_Display/n4372 ,\u2_Display/n4370 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2966|_al_u2972  (
    .b({\u2_Display/n4348 [11],\u2_Display/n4348 [17]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4334 ,\u2_Display/n4328 }),
    .f({\u2_Display/n4369 ,\u2_Display/n4363 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2967|_al_u2969  (
    .b({\u2_Display/n4348 [12],\u2_Display/n4348 [14]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4333 ,\u2_Display/n4331 }),
    .f({\u2_Display/n4368 ,\u2_Display/n4366 }));
  EG_PHY_PAD #(
    //.LOCATION("H16"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u297 (
    .do({open_n24712,open_n24713,open_n24714,vga_de_pad}),
    .opad(vga_de));  // source/rtl/VGA_Demo.v(13)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2970|_al_u2975  (
    .b({\u2_Display/n4348 [15],\u2_Display/n4348 [20]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4330 ,\u2_Display/n4325 }),
    .f({\u2_Display/n4365 ,\u2_Display/n4360 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2971|_al_u2973  (
    .b({\u2_Display/n4348 [16],\u2_Display/n4348 [18]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4329 ,\u2_Display/n4327 }),
    .f({\u2_Display/n4364 ,\u2_Display/n4362 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2974|_al_u2977  (
    .b({\u2_Display/n4348 [19],\u2_Display/n4348 [22]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4326 ,\u2_Display/n4323 }),
    .f({\u2_Display/n4361 ,\u2_Display/n4358 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2976|_al_u2979  (
    .b({\u2_Display/n4348 [21],\u2_Display/n4348 [24]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4324 ,\u2_Display/n4321 }),
    .f({\u2_Display/n4359 ,\u2_Display/n4356 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2978|_al_u2981  (
    .b({\u2_Display/n4348 [23],\u2_Display/n4348 [26]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4322 ,\u2_Display/n4319 }),
    .f({\u2_Display/n4357 ,\u2_Display/n4354 }));
  EG_PHY_PAD #(
    //.LOCATION("H5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u298 (
    .do({open_n24859,open_n24860,open_n24861,vga_b_pad[0]}),
    .opad(vga_g[7]));  // source/rtl/VGA_Demo.v(16)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2980|_al_u2984  (
    .b({\u2_Display/n4348 [25],\u2_Display/n4348 [29]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4320 ,\u2_Display/n4316 }),
    .f({\u2_Display/n4355 ,\u2_Display/n4351 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2982|_al_u2986  (
    .b({\u2_Display/n4348 [27],\u2_Display/n4348 [31]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4318 ,\u2_Display/n4314 }),
    .f({\u2_Display/n4353 ,\u2_Display/n4349 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2983|_al_u2985  (
    .b({\u2_Display/n4348 [28],\u2_Display/n4348 [30]}),
    .c({\u2_Display/n4346 ,\u2_Display/n4346 }),
    .d({\u2_Display/n4317 ,\u2_Display/n4315 }),
    .f({\u2_Display/n4352 ,\u2_Display/n4350 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2987|_al_u2989  (
    .b({\u2_Display/n5471 [0],\u2_Display/n5471 [2]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5468 ,\u2_Display/n5466 }),
    .f({\u2_Display/n5503 ,\u2_Display/n5501 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2988|_al_u2991  (
    .b({\u2_Display/n5471 [1],\u2_Display/n5471 [4]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5467 ,\u2_Display/n5464 }),
    .f({\u2_Display/n5502 ,\u2_Display/n5499 }));
  EG_PHY_PAD #(
    //.LOCATION("H1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u299 (
    .do({open_n25006,open_n25007,open_n25008,vga_b_pad[0]}),
    .opad(vga_g[6]));  // source/rtl/VGA_Demo.v(16)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2990|_al_u2993  (
    .b({\u2_Display/n5471 [3],\u2_Display/n5471 [6]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5465 ,\u2_Display/n5462 }),
    .f({\u2_Display/n5500 ,\u2_Display/n5497 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2992|_al_u2995  (
    .b({\u2_Display/n5471 [5],\u2_Display/n5471 [8]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5463 ,\u2_Display/n5460 }),
    .f({\u2_Display/n5498 ,\u2_Display/n5495 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2994|_al_u2997  (
    .b({\u2_Display/n5471 [7],\u2_Display/n5471 [10]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5461 ,\u2_Display/n5458 }),
    .f({\u2_Display/n5496 ,\u2_Display/n5493 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2996|_al_u3000  (
    .b({\u2_Display/n5471 [9],\u2_Display/n5471 [13]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5459 ,\u2_Display/n5455 }),
    .f({\u2_Display/n5494 ,\u2_Display/n5490 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2998|_al_u3003  (
    .b({\u2_Display/n5471 [11],\u2_Display/n5471 [16]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5457 ,\u2_Display/n5452 }),
    .f({\u2_Display/n5492 ,\u2_Display/n5487 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2999|_al_u3001  (
    .b({\u2_Display/n5471 [12],\u2_Display/n5471 [14]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5456 ,\u2_Display/n5454 }),
    .f({\u2_Display/n5491 ,\u2_Display/n5489 }));
  EG_PHY_PAD #(
    //.LOCATION("J6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u300 (
    .do({open_n25179,open_n25180,open_n25181,vga_b_pad[0]}),
    .opad(vga_g[5]));  // source/rtl/VGA_Demo.v(16)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3002|_al_u3005  (
    .b({\u2_Display/n5471 [15],\u2_Display/n5471 [18]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5453 ,\u2_Display/n5450 }),
    .f({\u2_Display/n5488 ,\u2_Display/n5485 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3004|_al_u3008  (
    .b({\u2_Display/n5471 [17],\u2_Display/n5471 [21]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5451 ,\u2_Display/n5447 }),
    .f({\u2_Display/n5486 ,\u2_Display/n5482 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3006|_al_u3011  (
    .b({\u2_Display/n5471 [19],\u2_Display/n5471 [24]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5449 ,\u2_Display/n5444 }),
    .f({\u2_Display/n5484 ,\u2_Display/n5479 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3007|_al_u3009  (
    .b({\u2_Display/n5471 [20],\u2_Display/n5471 [22]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5448 ,\u2_Display/n5446 }),
    .f({\u2_Display/n5483 ,\u2_Display/n5481 }));
  EG_PHY_PAD #(
    //.LOCATION("H3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u301 (
    .do({open_n25300,open_n25301,open_n25302,vga_b_pad[0]}),
    .opad(vga_g[4]));  // source/rtl/VGA_Demo.v(16)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3010|_al_u3013  (
    .b({\u2_Display/n5471 [23],\u2_Display/n5471 [26]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5445 ,\u2_Display/n5442 }),
    .f({\u2_Display/n5480 ,\u2_Display/n5477 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3012|_al_u3015  (
    .b({\u2_Display/n5471 [25],\u2_Display/n5471 [28]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5443 ,\u2_Display/n5440 }),
    .f({\u2_Display/n5478 ,\u2_Display/n5475 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3014|_al_u3017  (
    .b({\u2_Display/n5471 [27],\u2_Display/n5471 [30]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5441 ,\u2_Display/n5438 }),
    .f({\u2_Display/n5476 ,\u2_Display/n5473 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3016|_al_u3018  (
    .b({\u2_Display/n5471 [29],\u2_Display/n5471 [31]}),
    .c({\u2_Display/n5469 ,\u2_Display/n5469 }),
    .d({\u2_Display/n5439 ,\u2_Display/n5437 }),
    .f({\u2_Display/n5474 ,\u2_Display/n5472 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3019|_al_u3023  (
    .b({\u2_Display/n979 [0],\u2_Display/n979 [4]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n976 ,\u2_Display/n972 }),
    .f({\u2_Display/n1011 ,\u2_Display/n1007 }));
  EG_PHY_PAD #(
    //.LOCATION("J1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u302 (
    .do({open_n25447,open_n25448,open_n25449,vga_b_pad[0]}),
    .opad(vga_g[3]));  // source/rtl/VGA_Demo.v(16)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3020|_al_u3021  (
    .b({\u2_Display/n979 [1],\u2_Display/n979 [2]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n975 ,\u2_Display/n974 }),
    .f({\u2_Display/n1010 ,\u2_Display/n1009 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3022|_al_u3025  (
    .b({\u2_Display/n979 [3],\u2_Display/n979 [6]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n973 ,\u2_Display/n970 }),
    .f({\u2_Display/n1008 ,\u2_Display/n1005 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3024|_al_u3028  (
    .b({\u2_Display/n979 [5],\u2_Display/n979 [9]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n971 ,\u2_Display/n967 }),
    .f({\u2_Display/n1006 ,\u2_Display/n1002 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3026|_al_u3031  (
    .b({\u2_Display/n979 [7],\u2_Display/n979 [12]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n969 ,\u2_Display/n964 }),
    .f({\u2_Display/n1004 ,\u2_Display/n999 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3027|_al_u3029  (
    .b({\u2_Display/n979 [8],\u2_Display/n979 [10]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n968 ,\u2_Display/n966 }),
    .f({\u2_Display/n1003 ,\u2_Display/n1001 }));
  EG_PHY_PAD #(
    //.LOCATION("K1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u303 (
    .do({open_n25594,open_n25595,open_n25596,vga_b_pad[0]}),
    .opad(vga_g[2]));  // source/rtl/VGA_Demo.v(16)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3030|_al_u3033  (
    .b({\u2_Display/n979 [11],\u2_Display/n979 [14]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n965 ,\u2_Display/n962 }),
    .f({\u2_Display/n1000 ,\u2_Display/n997 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3032|_al_u3036  (
    .b({\u2_Display/n979 [13],\u2_Display/n979 [17]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n963 ,\u2_Display/n959 }),
    .f({\u2_Display/n998 ,\u2_Display/n994 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3034|_al_u3039  (
    .b({\u2_Display/n979 [15],\u2_Display/n979 [20]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n961 ,\u2_Display/n956 }),
    .f({\u2_Display/n996 ,\u2_Display/n991 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3035|_al_u3037  (
    .b({\u2_Display/n979 [16],\u2_Display/n979 [18]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n960 ,\u2_Display/n958 }),
    .f({\u2_Display/n995 ,\u2_Display/n993 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3038|_al_u3041  (
    .b({\u2_Display/n979 [19],\u2_Display/n979 [22]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n957 ,\u2_Display/n954 }),
    .f({\u2_Display/n992 ,\u2_Display/n989 }));
  EG_PHY_PAD #(
    //.LOCATION("K2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u304 (
    .do({open_n25741,open_n25742,open_n25743,vga_b_pad[0]}),
    .opad(vga_g[1]));  // source/rtl/VGA_Demo.v(16)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3040|_al_u3043  (
    .b({\u2_Display/n979 [21],\u2_Display/n979 [24]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n955 ,\u2_Display/n952 }),
    .f({\u2_Display/n990 ,\u2_Display/n987 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3042|_al_u3045  (
    .b({\u2_Display/n979 [23],\u2_Display/n979 [26]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n953 ,\u2_Display/n950 }),
    .f({\u2_Display/n988 ,\u2_Display/n985 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3044|_al_u3047  (
    .b({\u2_Display/n979 [25],\u2_Display/n979 [28]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n951 ,\u2_Display/n948 }),
    .f({\u2_Display/n986 ,\u2_Display/n983 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3046|_al_u3049  (
    .b({\u2_Display/n979 [27],\u2_Display/n979 [30]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n949 ,\u2_Display/n946 }),
    .f({\u2_Display/n984 ,\u2_Display/n981 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3048|_al_u3050  (
    .b({\u2_Display/n979 [29],\u2_Display/n979 [31]}),
    .c({\u2_Display/n977 ,\u2_Display/n977 }),
    .d({\u2_Display/n947 ,\u2_Display/n945 }),
    .f({\u2_Display/n982 ,\u2_Display/n980 }));
  EG_PHY_PAD #(
    //.LOCATION("L1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u305 (
    .do({open_n25888,open_n25889,open_n25890,vga_b_pad[0]}),
    .opad(vga_g[0]));  // source/rtl/VGA_Demo.v(16)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3051|_al_u3053  (
    .b({\u2_Display/n2102 [0],\u2_Display/n2102 [2]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .d({\u2_Display/n2099 ,\u2_Display/n2097 }),
    .f({\u2_Display/n2134 ,\u2_Display/n2132 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3052|_al_u3055  (
    .b({\u2_Display/n2102 [1],\u2_Display/n2102 [4]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .d({\u2_Display/n2098 ,\u2_Display/n2095 }),
    .f({\u2_Display/n2133 ,\u2_Display/n2130 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3054|_al_u3057  (
    .b({\u2_Display/n2102 [3],\u2_Display/n2102 [6]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .d({\u2_Display/n2096 ,\u2_Display/n2093 }),
    .f({\u2_Display/n2131 ,\u2_Display/n2128 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3056|_al_u3060  (
    .b({\u2_Display/n2102 [5],\u2_Display/n2102 [9]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .d({\u2_Display/n2094 ,\u2_Display/n2090 }),
    .f({\u2_Display/n2129 ,\u2_Display/n2125 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3058|_al_u3063  (
    .b({\u2_Display/n2102 [7],\u2_Display/n2102 [12]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .d({\u2_Display/n2092 ,\u2_Display/n2087 }),
    .f({\u2_Display/n2127 ,\u2_Display/n2122 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3059|_al_u3061  (
    .b({\u2_Display/n2102 [8],\u2_Display/n2102 [10]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .d({\u2_Display/n2091 ,\u2_Display/n2089 }),
    .f({\u2_Display/n2126 ,\u2_Display/n2124 }));
  EG_PHY_PAD #(
    //.LOCATION("J3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u306 (
    .do({open_n26061,open_n26062,open_n26063,vga_hs_pad}),
    .opad(vga_hs));  // source/rtl/VGA_Demo.v(10)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3062|_al_u3065  (
    .b({\u2_Display/n2102 [11],\u2_Display/n2102 [14]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .d({\u2_Display/n2088 ,\u2_Display/n2085 }),
    .f({\u2_Display/n2123 ,\u2_Display/n2120 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3064|_al_u3068  (
    .b({\u2_Display/n2102 [13],\u2_Display/n2102 [17]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .d({\u2_Display/n2086 ,\u2_Display/n2082 }),
    .f({\u2_Display/n2121 ,\u2_Display/n2117 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3066|_al_u3071  (
    .b({\u2_Display/n2102 [15],\u2_Display/n2102 [20]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .d({\u2_Display/n2084 ,\u2_Display/n2079 }),
    .f({\u2_Display/n2119 ,\u2_Display/n2114 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3067|_al_u3069  (
    .b({\u2_Display/n2102 [16],\u2_Display/n2102 [18]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .d({\u2_Display/n2083 ,\u2_Display/n2081 }),
    .f({\u2_Display/n2118 ,\u2_Display/n2116 }));
  EG_PHY_PAD #(
    //.LOCATION("K6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u307 (
    .do({open_n26182,open_n26183,open_n26184,vga_b_pad[0]}),
    .opad(vga_r[7]));  // source/rtl/VGA_Demo.v(15)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3070|_al_u3073  (
    .b({\u2_Display/n2102 [19],\u2_Display/n2102 [22]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .d({\u2_Display/n2080 ,\u2_Display/n2077 }),
    .f({\u2_Display/n2115 ,\u2_Display/n2112 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3072|_al_u3076  (
    .b({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .c({\u2_Display/n2102 [21],\u2_Display/n2102 [25]}),
    .d({\u2_Display/n2078 ,\u2_Display/n2074 }),
    .f({\u2_Display/n2113 ,\u2_Display/n2109 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3074|_al_u3212  (
    .b({\u2_Display/n2102 [23],\u2_Display/n2137 [1]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2076 ,\u2_Display/n2133 }),
    .f({\u2_Display/n2111 ,\u2_Display/n2168 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3075|_al_u3077  (
    .b({\u2_Display/n2102 [24],\u2_Display/n2102 [26]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .d({\u2_Display/n2075 ,\u2_Display/n2073 }),
    .f({\u2_Display/n2110 ,\u2_Display/n2108 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    //.LUTF1("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUTG0("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    //.LUTG1("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT_LUTF0(16'b1101100011011000),
    .INIT_LUTF1(16'b1110010011100100),
    .INIT_LUTG0(16'b1101100011011000),
    .INIT_LUTG1(16'b1110010011100100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3078|_al_u3079  (
    .a({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .b({\u2_Display/n2102 [27],\u2_Display/n2071 }),
    .c({\u2_Display/n2072 ,\u2_Display/n2102 [28]}),
    .f({\u2_Display/n2107 ,\u2_Display/n2106 }));
  EG_PHY_PAD #(
    //.LOCATION("K3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u308 (
    .do({open_n26329,open_n26330,open_n26331,vga_b_pad[0]}),
    .opad(vga_r[6]));  // source/rtl/VGA_Demo.v(15)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3080|_al_u3081  (
    .b({\u2_Display/n2102 [29],\u2_Display/n2102 [30]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2100 }),
    .d({\u2_Display/n2070 ,\u2_Display/n2069 }),
    .f({\u2_Display/n2105 ,\u2_Display/n2104 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3082|_al_u3219  (
    .b({\u2_Display/n2102 [31],\u2_Display/n2137 [8]}),
    .c({\u2_Display/n2100 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2068 ,\u2_Display/n2126 }),
    .f({\u2_Display/n2103 ,\u2_Display/n2161 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3083|_al_u3085  (
    .b({\u2_Display/n3225 [0],\u2_Display/n3225 [2]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3222 ,\u2_Display/n3220 }),
    .f({\u2_Display/n3257 ,\u2_Display/n3255 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3086|_al_u3089  (
    .b({\u2_Display/n3225 [3],\u2_Display/n3225 [6]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3219 ,\u2_Display/n3216 }),
    .f({\u2_Display/n3254 ,\u2_Display/n3251 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3087|_al_u3088  (
    .b({\u2_Display/n3225 [4],\u2_Display/n3225 [5]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3218 ,\u2_Display/n3217 }),
    .f({\u2_Display/n3253 ,\u2_Display/n3252 }));
  EG_PHY_PAD #(
    //.LOCATION("K5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u309 (
    .do({open_n26476,open_n26477,open_n26478,vga_b_pad[0]}),
    .opad(vga_r[5]));  // source/rtl/VGA_Demo.v(15)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3090|_al_u3093  (
    .b({\u2_Display/n3225 [7],\u2_Display/n3225 [10]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3215 ,\u2_Display/n3212 }),
    .f({\u2_Display/n3250 ,\u2_Display/n3247 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3092|_al_u3095  (
    .b({\u2_Display/n3225 [9],\u2_Display/n3225 [12]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3213 ,\u2_Display/n3210 }),
    .f({\u2_Display/n3248 ,\u2_Display/n3245 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3094|_al_u3097  (
    .b({\u2_Display/n3225 [11],\u2_Display/n3225 [14]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3211 ,\u2_Display/n3208 }),
    .f({\u2_Display/n3246 ,\u2_Display/n3243 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3096|_al_u3100  (
    .b({\u2_Display/n3225 [13],\u2_Display/n3225 [17]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3209 ,\u2_Display/n3205 }),
    .f({\u2_Display/n3244 ,\u2_Display/n3240 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3098|_al_u3103  (
    .b({\u2_Display/n3225 [15],\u2_Display/n3225 [20]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3207 ,\u2_Display/n3202 }),
    .f({\u2_Display/n3242 ,\u2_Display/n3237 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3099|_al_u3101  (
    .b({\u2_Display/n3225 [16],\u2_Display/n3225 [18]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3206 ,\u2_Display/n3204 }),
    .f({\u2_Display/n3241 ,\u2_Display/n3239 }));
  EG_PHY_PAD #(
    //.LOCATION("L4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u310 (
    .do({open_n26649,open_n26650,open_n26651,vga_b_pad[0]}),
    .opad(vga_r[4]));  // source/rtl/VGA_Demo.v(15)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3102|_al_u3105  (
    .b({\u2_Display/n3225 [19],\u2_Display/n3225 [22]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3203 ,\u2_Display/n3200 }),
    .f({\u2_Display/n3238 ,\u2_Display/n3235 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3104|_al_u3107  (
    .b({\u2_Display/n3225 [21],\u2_Display/n3225 [24]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3201 ,\u2_Display/n3198 }),
    .f({\u2_Display/n3236 ,\u2_Display/n3233 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3106|_al_u3244  (
    .b({\u2_Display/n3225 [23],\u2_Display/n3260 [1]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3199 ,\u2_Display/n3256 }),
    .f({\u2_Display/n3234 ,\u2_Display/n3291 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUTF1("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    //.LUTG0("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUTG1("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    .INIT_LUTF0(16'b1110010011100100),
    .INIT_LUTF1(16'b1110111001000100),
    .INIT_LUTG0(16'b1110010011100100),
    .INIT_LUTG1(16'b1110111001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3108|_al_u3109  (
    .a({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .b({\u2_Display/n3225 [25],\u2_Display/n3225 [26]}),
    .c({open_n26743,\u2_Display/n3196 }),
    .d({\u2_Display/n3197 ,open_n26746}),
    .f({\u2_Display/n3232 ,\u2_Display/n3231 }));
  EG_PHY_PAD #(
    //.LOCATION("M1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u311 (
    .do({open_n26770,open_n26771,open_n26772,vga_b_pad[0]}),
    .opad(vga_r[3]));  // source/rtl/VGA_Demo.v(15)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3110|_al_u3111  (
    .b({\u2_Display/n3225 [27],\u2_Display/n3225 [28]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3195 ,\u2_Display/n3194 }),
    .f({\u2_Display/n3230 ,\u2_Display/n3229 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3112|_al_u3113  (
    .b({\u2_Display/n3225 [29],\u2_Display/n3225 [30]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3223 }),
    .d({\u2_Display/n3193 ,\u2_Display/n3192 }),
    .f({\u2_Display/n3228 ,\u2_Display/n3227 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3114|_al_u3252  (
    .b({\u2_Display/n3225 [31],\u2_Display/n3260 [9]}),
    .c({\u2_Display/n3223 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3191 ,\u2_Display/n3248 }),
    .f({\u2_Display/n3226 ,\u2_Display/n3283 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3115|_al_u3117  (
    .b({\u2_Display/n4383 [0],\u2_Display/n4383 [2]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4380 ,\u2_Display/n4378 }),
    .f({\u2_Display/n4415 ,\u2_Display/n4413 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3116|_al_u3119  (
    .b({\u2_Display/n4383 [1],\u2_Display/n4383 [4]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4379 ,\u2_Display/n4376 }),
    .f({\u2_Display/n4414 ,\u2_Display/n4411 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3118|_al_u3121  (
    .b({\u2_Display/n4383 [3],\u2_Display/n4383 [6]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4377 ,\u2_Display/n4374 }),
    .f({\u2_Display/n4412 ,\u2_Display/n4409 }));
  EG_PHY_PAD #(
    //.LOCATION("M2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u312 (
    .do({open_n26943,open_n26944,open_n26945,vga_b_pad[0]}),
    .opad(vga_r[2]));  // source/rtl/VGA_Demo.v(15)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3120|_al_u3124  (
    .b({\u2_Display/n4383 [5],\u2_Display/n4383 [9]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4375 ,\u2_Display/n4371 }),
    .f({\u2_Display/n4410 ,\u2_Display/n4406 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3122|_al_u3128  (
    .b({\u2_Display/n4383 [7],\u2_Display/n4383 [13]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4373 ,\u2_Display/n4367 }),
    .f({\u2_Display/n4408 ,\u2_Display/n4402 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3123|_al_u3125  (
    .b({\u2_Display/n4383 [8],\u2_Display/n4383 [10]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4372 ,\u2_Display/n4370 }),
    .f({\u2_Display/n4407 ,\u2_Display/n4405 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3126|_al_u3131  (
    .b({\u2_Display/n4383 [11],\u2_Display/n4383 [16]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4369 ,\u2_Display/n4364 }),
    .f({\u2_Display/n4404 ,\u2_Display/n4399 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3127|_al_u3129  (
    .b({\u2_Display/n4383 [12],\u2_Display/n4383 [14]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4368 ,\u2_Display/n4366 }),
    .f({\u2_Display/n4403 ,\u2_Display/n4401 }));
  EG_PHY_PAD #(
    //.LOCATION("L3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u313 (
    .do({open_n27090,open_n27091,open_n27092,vga_b_pad[0]}),
    .opad(vga_r[1]));  // source/rtl/VGA_Demo.v(15)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3130|_al_u3133  (
    .b({\u2_Display/n4383 [15],\u2_Display/n4383 [18]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4365 ,\u2_Display/n4362 }),
    .f({\u2_Display/n4400 ,\u2_Display/n4397 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3132|_al_u3136  (
    .b({\u2_Display/n4383 [17],\u2_Display/n4383 [21]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4363 ,\u2_Display/n4359 }),
    .f({\u2_Display/n4398 ,\u2_Display/n4394 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3134|_al_u3139  (
    .b({\u2_Display/n4383 [19],\u2_Display/n4383 [24]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4361 ,\u2_Display/n4356 }),
    .f({\u2_Display/n4396 ,\u2_Display/n4391 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3135|_al_u3137  (
    .b({\u2_Display/n4383 [20],\u2_Display/n4383 [22]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4360 ,\u2_Display/n4358 }),
    .f({\u2_Display/n4395 ,\u2_Display/n4393 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3138|_al_u3141  (
    .b({\u2_Display/n4383 [23],\u2_Display/n4383 [26]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4357 ,\u2_Display/n4354 }),
    .f({\u2_Display/n4392 ,\u2_Display/n4389 }));
  EG_PHY_PAD #(
    //.LOCATION("L5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u314 (
    .do({open_n27237,open_n27238,open_n27239,vga_b_pad[0]}),
    .opad(vga_r[0]));  // source/rtl/VGA_Demo.v(15)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3140|_al_u3144  (
    .b({\u2_Display/n4383 [25],\u2_Display/n4383 [29]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4355 ,\u2_Display/n4351 }),
    .f({\u2_Display/n4390 ,\u2_Display/n4386 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3142|_al_u3146  (
    .b({\u2_Display/n4383 [27],\u2_Display/n4383 [31]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4353 ,\u2_Display/n4349 }),
    .f({\u2_Display/n4388 ,\u2_Display/n4384 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3143|_al_u3145  (
    .b({\u2_Display/n4383 [28],\u2_Display/n4383 [30]}),
    .c({\u2_Display/n4381 ,\u2_Display/n4381 }),
    .d({\u2_Display/n4352 ,\u2_Display/n4350 }),
    .f({\u2_Display/n4387 ,\u2_Display/n4385 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3147|_al_u3152  (
    .b({\u2_Display/n5506 [0],\u2_Display/n5506 [5]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5503 ,\u2_Display/n5498 }),
    .f({\u2_Display/n5538 ,\u2_Display/n5533 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3148|_al_u3149  (
    .b({\u2_Display/n5506 [1],\u2_Display/n5506 [2]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5502 ,\u2_Display/n5501 }),
    .f({\u2_Display/n5537 ,\u2_Display/n5536 }));
  EG_PHY_PAD #(
    //.LOCATION("J4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u315 (
    .do({open_n27384,open_n27385,open_n27386,vga_vs_pad}),
    .opad(vga_vs));  // source/rtl/VGA_Demo.v(11)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3150|_al_u3156  (
    .b({\u2_Display/n5506 [3],\u2_Display/n5506 [9]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5500 ,\u2_Display/n5494 }),
    .f({\u2_Display/n5535 ,\u2_Display/n5529 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3151|_al_u3153  (
    .b({\u2_Display/n5506 [4],\u2_Display/n5506 [6]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5499 ,\u2_Display/n5497 }),
    .f({\u2_Display/n5534 ,\u2_Display/n5532 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3154|_al_u3160  (
    .b({\u2_Display/n5506 [7],\u2_Display/n5506 [13]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5496 ,\u2_Display/n5490 }),
    .f({\u2_Display/n5531 ,\u2_Display/n5525 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3155|_al_u3157  (
    .b({\u2_Display/n5506 [8],\u2_Display/n5506 [10]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5495 ,\u2_Display/n5493 }),
    .f({\u2_Display/n5530 ,\u2_Display/n5528 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3158|_al_u3164  (
    .b({\u2_Display/n5506 [11],\u2_Display/n5506 [17]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5492 ,\u2_Display/n5486 }),
    .f({\u2_Display/n5527 ,\u2_Display/n5521 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3159|_al_u3161  (
    .b({\u2_Display/n5506 [12],\u2_Display/n5506 [14]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5491 ,\u2_Display/n5489 }),
    .f({\u2_Display/n5526 ,\u2_Display/n5524 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3162|_al_u3167  (
    .b({\u2_Display/n5506 [15],\u2_Display/n5506 [20]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5488 ,\u2_Display/n5483 }),
    .f({\u2_Display/n5523 ,\u2_Display/n5518 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3163|_al_u3165  (
    .b({\u2_Display/n5506 [16],\u2_Display/n5506 [18]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5487 ,\u2_Display/n5485 }),
    .f({\u2_Display/n5522 ,\u2_Display/n5520 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3166|_al_u3169  (
    .b({\u2_Display/n5506 [19],\u2_Display/n5506 [22]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5484 ,\u2_Display/n5481 }),
    .f({\u2_Display/n5519 ,\u2_Display/n5516 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3168|_al_u3171  (
    .b({\u2_Display/n5506 [21],\u2_Display/n5506 [24]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5482 ,\u2_Display/n5479 }),
    .f({\u2_Display/n5517 ,\u2_Display/n5514 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3170|_al_u3173  (
    .b({\u2_Display/n5506 [23],\u2_Display/n5506 [26]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5480 ,\u2_Display/n5477 }),
    .f({\u2_Display/n5515 ,\u2_Display/n5512 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3172|_al_u3175  (
    .b({\u2_Display/n5506 [25],\u2_Display/n5506 [28]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5478 ,\u2_Display/n5475 }),
    .f({\u2_Display/n5513 ,\u2_Display/n5510 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3174|_al_u3177  (
    .b({\u2_Display/n5506 [27],\u2_Display/n5506 [30]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5476 ,\u2_Display/n5473 }),
    .f({\u2_Display/n5511 ,\u2_Display/n5508 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3176|_al_u3178  (
    .b({\u2_Display/n5506 [29],\u2_Display/n5506 [31]}),
    .c({\u2_Display/n5504 ,\u2_Display/n5504 }),
    .d({\u2_Display/n5474 ,\u2_Display/n5472 }),
    .f({\u2_Display/n5509 ,\u2_Display/n5507 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3179|_al_u3181  (
    .b({\u2_Display/n1014 [0],\u2_Display/n1014 [2]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n1011 ,\u2_Display/n1009 }),
    .f({\u2_Display/n1046 ,\u2_Display/n1044 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3180|_al_u3183  (
    .b({\u2_Display/n1014 [1],\u2_Display/n1014 [4]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n1010 ,\u2_Display/n1007 }),
    .f({\u2_Display/n1045 ,\u2_Display/n1042 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3182|_al_u3185  (
    .b({\u2_Display/n1014 [3],\u2_Display/n1014 [6]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n1008 ,\u2_Display/n1005 }),
    .f({\u2_Display/n1043 ,\u2_Display/n1040 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3184|_al_u3188  (
    .b({\u2_Display/n1014 [5],\u2_Display/n1014 [9]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n1006 ,\u2_Display/n1002 }),
    .f({\u2_Display/n1041 ,\u2_Display/n1037 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3186|_al_u3191  (
    .b({\u2_Display/n1014 [7],\u2_Display/n1014 [12]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n1004 ,\u2_Display/n999 }),
    .f({\u2_Display/n1039 ,\u2_Display/n1034 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3187|_al_u3189  (
    .b({\u2_Display/n1014 [8],\u2_Display/n1014 [10]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n1003 ,\u2_Display/n1001 }),
    .f({\u2_Display/n1038 ,\u2_Display/n1036 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3190|_al_u3193  (
    .b({\u2_Display/n1014 [11],\u2_Display/n1014 [14]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n1000 ,\u2_Display/n997 }),
    .f({\u2_Display/n1035 ,\u2_Display/n1032 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3192|_al_u3196  (
    .b({\u2_Display/n1014 [13],\u2_Display/n1014 [17]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n998 ,\u2_Display/n994 }),
    .f({\u2_Display/n1033 ,\u2_Display/n1029 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3194|_al_u3199  (
    .b({\u2_Display/n1014 [15],\u2_Display/n1014 [20]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n996 ,\u2_Display/n991 }),
    .f({\u2_Display/n1031 ,\u2_Display/n1026 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3195|_al_u3197  (
    .b({\u2_Display/n1014 [16],\u2_Display/n1014 [18]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n995 ,\u2_Display/n993 }),
    .f({\u2_Display/n1030 ,\u2_Display/n1028 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3198|_al_u3201  (
    .b({\u2_Display/n1014 [19],\u2_Display/n1014 [22]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n992 ,\u2_Display/n989 }),
    .f({\u2_Display/n1027 ,\u2_Display/n1024 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3200|_al_u3203  (
    .b({\u2_Display/n1014 [21],\u2_Display/n1014 [24]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n990 ,\u2_Display/n987 }),
    .f({\u2_Display/n1025 ,\u2_Display/n1022 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3202|_al_u3205  (
    .b({\u2_Display/n1014 [23],\u2_Display/n1014 [26]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n988 ,\u2_Display/n985 }),
    .f({\u2_Display/n1023 ,\u2_Display/n1020 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3204|_al_u3207  (
    .b({\u2_Display/n1014 [25],\u2_Display/n1014 [28]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n986 ,\u2_Display/n983 }),
    .f({\u2_Display/n1021 ,\u2_Display/n1018 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3206|_al_u3209  (
    .b({\u2_Display/n1014 [27],\u2_Display/n1014 [30]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n984 ,\u2_Display/n981 }),
    .f({\u2_Display/n1019 ,\u2_Display/n1016 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3208|_al_u3210  (
    .b({\u2_Display/n1014 [29],\u2_Display/n1014 [31]}),
    .c({\u2_Display/n1012 ,\u2_Display/n1012 }),
    .d({\u2_Display/n982 ,\u2_Display/n980 }),
    .f({\u2_Display/n1017 ,\u2_Display/n1015 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3211|_al_u3213  (
    .b({\u2_Display/n2137 [0],\u2_Display/n2137 [2]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2134 ,\u2_Display/n2132 }),
    .f({\u2_Display/n2169 ,\u2_Display/n2167 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3214|_al_u3217  (
    .b({\u2_Display/n2137 [3],\u2_Display/n2137 [6]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2131 ,\u2_Display/n2128 }),
    .f({\u2_Display/n2166 ,\u2_Display/n2163 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3215|_al_u3216  (
    .b({\u2_Display/n2137 [4],\u2_Display/n2137 [5]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2130 ,\u2_Display/n2129 }),
    .f({\u2_Display/n2165 ,\u2_Display/n2164 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3218|_al_u3221  (
    .b({\u2_Display/n2137 [7],\u2_Display/n2137 [10]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2127 ,\u2_Display/n2124 }),
    .f({\u2_Display/n2162 ,\u2_Display/n2159 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3220|_al_u3223  (
    .b({\u2_Display/n2137 [9],\u2_Display/n2137 [12]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2125 ,\u2_Display/n2122 }),
    .f({\u2_Display/n2160 ,\u2_Display/n2157 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3222|_al_u3225  (
    .b({\u2_Display/n2137 [11],\u2_Display/n2137 [14]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2123 ,\u2_Display/n2120 }),
    .f({\u2_Display/n2158 ,\u2_Display/n2155 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3224|_al_u3228  (
    .b({\u2_Display/n2137 [13],\u2_Display/n2137 [17]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2121 ,\u2_Display/n2117 }),
    .f({\u2_Display/n2156 ,\u2_Display/n2152 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3226|_al_u3232  (
    .b({\u2_Display/n2137 [15],\u2_Display/n2137 [21]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2119 ,\u2_Display/n2113 }),
    .f({\u2_Display/n2154 ,\u2_Display/n2148 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3227|_al_u3229  (
    .b({\u2_Display/n2137 [16],\u2_Display/n2137 [18]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2118 ,\u2_Display/n2116 }),
    .f({\u2_Display/n2153 ,\u2_Display/n2151 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3230|_al_u3235  (
    .b({\u2_Display/n2137 [19],\u2_Display/n2137 [24]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2115 ,\u2_Display/n2110 }),
    .f({\u2_Display/n2150 ,\u2_Display/n2145 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3231|_al_u3233  (
    .b({\u2_Display/n2137 [20],\u2_Display/n2137 [22]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2114 ,\u2_Display/n2112 }),
    .f({\u2_Display/n2149 ,\u2_Display/n2147 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3234|_al_u3371  (
    .b({\u2_Display/n2135 ,\u2_Display/n2172 [0]}),
    .c({\u2_Display/n2137 [23],\u2_Display/n2170 }),
    .d({\u2_Display/n2111 ,\u2_Display/n2169 }),
    .f({\u2_Display/n2146 ,\u2_Display/n2204 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTF1("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    //.LUTG0("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTG1("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    .INIT_LUTF0(16'b1111101001010000),
    .INIT_LUTF1(16'b1110111001000100),
    .INIT_LUTG0(16'b1111101001010000),
    .INIT_LUTG1(16'b1110111001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3236|_al_u3237  (
    .a({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .b({\u2_Display/n2137 [25],open_n28492}),
    .c({open_n28493,\u2_Display/n2137 [26]}),
    .d({\u2_Display/n2109 ,\u2_Display/n2108 }),
    .f({\u2_Display/n2144 ,\u2_Display/n2143 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3238|_al_u3241  (
    .b({\u2_Display/n2137 [27],\u2_Display/n2137 [30]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2107 ,\u2_Display/n2104 }),
    .f({\u2_Display/n2142 ,\u2_Display/n2139 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3239|_al_u3240  (
    .b({\u2_Display/n2137 [28],\u2_Display/n2137 [29]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2135 }),
    .d({\u2_Display/n2106 ,\u2_Display/n2105 }),
    .f({\u2_Display/n2141 ,\u2_Display/n2140 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3242|_al_u3379  (
    .b({\u2_Display/n2137 [31],\u2_Display/n2172 [8]}),
    .c({\u2_Display/n2135 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2103 ,\u2_Display/n2161 }),
    .f({\u2_Display/n2138 ,\u2_Display/n2196 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3243|_al_u3245  (
    .b({\u2_Display/n3260 [0],\u2_Display/n3260 [2]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3257 ,\u2_Display/n3255 }),
    .f({\u2_Display/n3292 ,\u2_Display/n3290 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3246|_al_u3249  (
    .b({\u2_Display/n3260 [3],\u2_Display/n3260 [6]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3254 ,\u2_Display/n3251 }),
    .f({\u2_Display/n3289 ,\u2_Display/n3286 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3247|_al_u3248  (
    .b({\u2_Display/n3260 [4],\u2_Display/n3260 [5]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3253 ,\u2_Display/n3252 }),
    .f({\u2_Display/n3288 ,\u2_Display/n3287 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3250|_al_u3255  (
    .b({\u2_Display/n3260 [7],\u2_Display/n3260 [12]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3250 ,\u2_Display/n3245 }),
    .f({\u2_Display/n3285 ,\u2_Display/n3280 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3251|_al_u3253  (
    .b({\u2_Display/n3260 [8],\u2_Display/n3260 [10]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3249 ,\u2_Display/n3247 }),
    .f({\u2_Display/n3284 ,\u2_Display/n3282 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3254|_al_u3257  (
    .b({\u2_Display/n3260 [11],\u2_Display/n3260 [14]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3246 ,\u2_Display/n3243 }),
    .f({\u2_Display/n3281 ,\u2_Display/n3278 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3256|_al_u3260  (
    .b({\u2_Display/n3260 [13],\u2_Display/n3260 [17]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3244 ,\u2_Display/n3240 }),
    .f({\u2_Display/n3279 ,\u2_Display/n3275 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3258|_al_u3264  (
    .b({\u2_Display/n3260 [15],\u2_Display/n3260 [21]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3242 ,\u2_Display/n3236 }),
    .f({\u2_Display/n3277 ,\u2_Display/n3271 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3259|_al_u3261  (
    .b({\u2_Display/n3260 [16],\u2_Display/n3260 [18]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3241 ,\u2_Display/n3239 }),
    .f({\u2_Display/n3276 ,\u2_Display/n3274 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3262|_al_u3267  (
    .b({\u2_Display/n3260 [19],\u2_Display/n3260 [24]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3238 ,\u2_Display/n3233 }),
    .f({\u2_Display/n3273 ,\u2_Display/n3268 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3263|_al_u3265  (
    .b({\u2_Display/n3260 [20],\u2_Display/n3260 [22]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3237 ,\u2_Display/n3235 }),
    .f({\u2_Display/n3272 ,\u2_Display/n3270 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3266|_al_u3404  (
    .b({\u2_Display/n3260 [23],\u2_Display/n3295 [1]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3234 ,\u2_Display/n3291 }),
    .f({\u2_Display/n3269 ,\u2_Display/n3326 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3268|_al_u3269  (
    .b({\u2_Display/n3260 [25],\u2_Display/n3260 [26]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3232 ,\u2_Display/n3231 }),
    .f({\u2_Display/n3267 ,\u2_Display/n3266 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3270|_al_u3273  (
    .b({\u2_Display/n3260 [27],\u2_Display/n3260 [30]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3230 ,\u2_Display/n3227 }),
    .f({\u2_Display/n3265 ,\u2_Display/n3262 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3271|_al_u3272  (
    .b({\u2_Display/n3260 [28],\u2_Display/n3260 [29]}),
    .c({\u2_Display/n3258 ,\u2_Display/n3258 }),
    .d({\u2_Display/n3229 ,\u2_Display/n3228 }),
    .f({\u2_Display/n3264 ,\u2_Display/n3263 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111101001010000),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111101001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3274|_al_u3416  (
    .a({\u2_Display/n3258 ,open_n28986}),
    .b({open_n28987,\u2_Display/n3295 [13]}),
    .c({\u2_Display/n3260 [31],\u2_Display/n3293 }),
    .d({\u2_Display/n3226 ,\u2_Display/n3279 }),
    .f({\u2_Display/n3261 ,\u2_Display/n3314 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3275|_al_u3279  (
    .b({\u2_Display/n4418 [0],\u2_Display/n4418 [4]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4415 ,\u2_Display/n4411 }),
    .f({\u2_Display/n4450 ,\u2_Display/n4446 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3276|_al_u3277  (
    .b({\u2_Display/n4418 [1],\u2_Display/n4418 [2]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4414 ,\u2_Display/n4413 }),
    .f({\u2_Display/n4449 ,\u2_Display/n4448 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3278|_al_u3281  (
    .b({\u2_Display/n4418 [3],\u2_Display/n4418 [6]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4412 ,\u2_Display/n4409 }),
    .f({\u2_Display/n4447 ,\u2_Display/n4444 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3280|_al_u3283  (
    .b({\u2_Display/n4418 [5],\u2_Display/n4418 [8]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4410 ,\u2_Display/n4407 }),
    .f({\u2_Display/n4445 ,\u2_Display/n4442 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3282|_al_u3285  (
    .b({\u2_Display/n4418 [7],\u2_Display/n4418 [10]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4408 ,\u2_Display/n4405 }),
    .f({\u2_Display/n4443 ,\u2_Display/n4440 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3284|_al_u3287  (
    .b({\u2_Display/n4418 [9],\u2_Display/n4418 [12]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4406 ,\u2_Display/n4403 }),
    .f({\u2_Display/n4441 ,\u2_Display/n4438 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3286|_al_u3289  (
    .b({\u2_Display/n4418 [11],\u2_Display/n4418 [14]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4404 ,\u2_Display/n4401 }),
    .f({\u2_Display/n4439 ,\u2_Display/n4436 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3288|_al_u3292  (
    .b({\u2_Display/n4418 [13],\u2_Display/n4418 [17]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4402 ,\u2_Display/n4398 }),
    .f({\u2_Display/n4437 ,\u2_Display/n4433 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C@D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111111110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u328|_al_u329  (
    .c({\u2_Display/i [9],\u2_Display/i [9]}),
    .d({\u2_Display/i [10],\u2_Display/i [10]}),
    .f({\u2_Display/add7_2_co ,\u2_Display/n140 [1]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3290|_al_u3295  (
    .b({\u2_Display/n4418 [15],\u2_Display/n4418 [20]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4400 ,\u2_Display/n4395 }),
    .f({\u2_Display/n4435 ,\u2_Display/n4430 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3291|_al_u3293  (
    .b({\u2_Display/n4418 [16],\u2_Display/n4418 [18]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4399 ,\u2_Display/n4397 }),
    .f({\u2_Display/n4434 ,\u2_Display/n4432 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3294|_al_u3297  (
    .b({\u2_Display/n4418 [19],\u2_Display/n4418 [22]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4396 ,\u2_Display/n4393 }),
    .f({\u2_Display/n4431 ,\u2_Display/n4428 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3296|_al_u3300  (
    .b({\u2_Display/n4418 [21],\u2_Display/n4418 [25]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4394 ,\u2_Display/n4390 }),
    .f({\u2_Display/n4429 ,\u2_Display/n4425 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3298|_al_u3304  (
    .b({\u2_Display/n4418 [23],\u2_Display/n4418 [29]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4392 ,\u2_Display/n4386 }),
    .f({\u2_Display/n4427 ,\u2_Display/n4421 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3299|_al_u3301  (
    .b({\u2_Display/n4418 [24],\u2_Display/n4418 [26]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4391 ,\u2_Display/n4389 }),
    .f({\u2_Display/n4426 ,\u2_Display/n4424 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTG0("(D*C*B*A)"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u330 (
    .a({open_n29400,\u1_Driver/n11 }),
    .b({open_n29401,\u1_Driver/n12 }),
    .c({open_n29402,\u1_Driver/n14 }),
    .d({open_n29405,\u1_Driver/n15 }),
    .f({open_n29423,vga_de_pad}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3302|_al_u3306  (
    .b({\u2_Display/n4418 [27],\u2_Display/n4418 [31]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4388 ,\u2_Display/n4384 }),
    .f({\u2_Display/n4423 ,\u2_Display/n4419 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3303|_al_u3305  (
    .b({\u2_Display/n4418 [28],\u2_Display/n4418 [30]}),
    .c({\u2_Display/n4416 ,\u2_Display/n4416 }),
    .d({\u2_Display/n4387 ,\u2_Display/n4385 }),
    .f({\u2_Display/n4422 ,\u2_Display/n4420 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3307|_al_u3311  (
    .b({\u2_Display/n5541 [0],\u2_Display/n5541 [4]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5538 ,\u2_Display/n5534 }),
    .f({\u2_Display/n5573 ,\u2_Display/n5569 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3308|_al_u3309  (
    .b({\u2_Display/n5541 [1],\u2_Display/n5541 [2]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5537 ,\u2_Display/n5536 }),
    .f({\u2_Display/n5572 ,\u2_Display/n5571 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3310|_al_u3313  (
    .b({\u2_Display/n5541 [3],\u2_Display/n5541 [6]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5535 ,\u2_Display/n5532 }),
    .f({\u2_Display/n5570 ,\u2_Display/n5567 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3312|_al_u3315  (
    .b({\u2_Display/n5541 [5],\u2_Display/n5541 [8]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5533 ,\u2_Display/n5530 }),
    .f({\u2_Display/n5568 ,\u2_Display/n5565 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3314|_al_u3317  (
    .b({\u2_Display/n5541 [7],\u2_Display/n5541 [10]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5531 ,\u2_Display/n5528 }),
    .f({\u2_Display/n5566 ,\u2_Display/n5563 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3316|_al_u3319  (
    .b({\u2_Display/n5541 [9],\u2_Display/n5541 [12]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5529 ,\u2_Display/n5526 }),
    .f({\u2_Display/n5564 ,\u2_Display/n5561 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3318|_al_u3321  (
    .b({\u2_Display/n5541 [11],\u2_Display/n5541 [14]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5527 ,\u2_Display/n5524 }),
    .f({\u2_Display/n5562 ,\u2_Display/n5559 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u331|_al_u333  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [0],\u2_Display/counta [2]}),
    .d({\u2_Display/n3788 [0],\u2_Display/n3788 [2]}),
    .f({\u2_Display/n3820 ,\u2_Display/n3818 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u332 (
    .b({open_n29691,\u2_Display/n3786 }),
    .c({open_n29692,\u2_Display/counta [1]}),
    .d({open_n29695,\u2_Display/n3788 [1]}),
    .f({open_n29713,\u2_Display/n3819 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3320|_al_u3324  (
    .b({\u2_Display/n5541 [13],\u2_Display/n5541 [17]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5525 ,\u2_Display/n5521 }),
    .f({\u2_Display/n5560 ,\u2_Display/n5556 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3322|_al_u3328  (
    .b({\u2_Display/n5541 [15],\u2_Display/n5541 [21]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5523 ,\u2_Display/n5517 }),
    .f({\u2_Display/n5558 ,\u2_Display/n5552 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3323|_al_u3325  (
    .b({\u2_Display/n5541 [16],\u2_Display/n5541 [18]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5522 ,\u2_Display/n5520 }),
    .f({\u2_Display/n5557 ,\u2_Display/n5555 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3326|_al_u3331  (
    .b({\u2_Display/n5541 [19],\u2_Display/n5541 [24]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5519 ,\u2_Display/n5514 }),
    .f({\u2_Display/n5554 ,\u2_Display/n5549 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3327|_al_u3329  (
    .b({\u2_Display/n5541 [20],\u2_Display/n5541 [22]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5518 ,\u2_Display/n5516 }),
    .f({\u2_Display/n5553 ,\u2_Display/n5551 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3330|_al_u3333  (
    .b({\u2_Display/n5541 [23],\u2_Display/n5541 [26]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5515 ,\u2_Display/n5512 }),
    .f({\u2_Display/n5550 ,\u2_Display/n5547 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3332|_al_u3335  (
    .b({\u2_Display/n5541 [25],\u2_Display/n5541 [28]}),
    .c({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .d({\u2_Display/n5513 ,\u2_Display/n5510 }),
    .f({\u2_Display/n5548 ,\u2_Display/n5545 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    //.LUTF1("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    //.LUTG0("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    //.LUTG1("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    .INIT_LUTF0(16'b1101100011011000),
    .INIT_LUTF1(16'b1110111001000100),
    .INIT_LUTG0(16'b1101100011011000),
    .INIT_LUTG1(16'b1110111001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3334|_al_u3337  (
    .a({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .b({\u2_Display/n5541 [27],\u2_Display/n5508 }),
    .c({open_n29901,\u2_Display/n5541 [30]}),
    .d({\u2_Display/n5511 ,open_n29904}),
    .f({\u2_Display/n5546 ,\u2_Display/n5543 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3336|_al_u3338  (
    .b({\u2_Display/n5539 ,\u2_Display/n5539 }),
    .c({\u2_Display/n5541 [29],\u2_Display/n5541 [31]}),
    .d({\u2_Display/n5509 ,\u2_Display/n5507 }),
    .f({\u2_Display/n5544 ,\u2_Display/n5542 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3339|_al_u3343  (
    .b({\u2_Display/n1049 [0],\u2_Display/n1049 [4]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1046 ,\u2_Display/n1042 }),
    .f({\u2_Display/n1081 ,\u2_Display/n1077 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3340|_al_u3341  (
    .b({\u2_Display/n1049 [1],\u2_Display/n1049 [2]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1045 ,\u2_Display/n1044 }),
    .f({\u2_Display/n1080 ,\u2_Display/n1079 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3342|_al_u3345  (
    .b({\u2_Display/n1049 [3],\u2_Display/n1049 [6]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1043 ,\u2_Display/n1040 }),
    .f({\u2_Display/n1078 ,\u2_Display/n1075 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3344|_al_u3347  (
    .b({\u2_Display/n1049 [5],\u2_Display/n1049 [8]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1041 ,\u2_Display/n1038 }),
    .f({\u2_Display/n1076 ,\u2_Display/n1073 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3346|_al_u3349  (
    .b({\u2_Display/n1049 [7],\u2_Display/n1049 [10]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1039 ,\u2_Display/n1036 }),
    .f({\u2_Display/n1074 ,\u2_Display/n1071 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3348|_al_u3351  (
    .b({\u2_Display/n1049 [9],\u2_Display/n1049 [12]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1037 ,\u2_Display/n1034 }),
    .f({\u2_Display/n1072 ,\u2_Display/n1069 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u334|_al_u337  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [3],\u2_Display/counta [6]}),
    .d({\u2_Display/n3788 [3],\u2_Display/n3788 [6]}),
    .f({\u2_Display/n3817 ,\u2_Display/n3814 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3350|_al_u3353  (
    .b({\u2_Display/n1049 [11],\u2_Display/n1049 [14]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1035 ,\u2_Display/n1032 }),
    .f({\u2_Display/n1070 ,\u2_Display/n1067 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3352|_al_u3355  (
    .b({\u2_Display/n1049 [13],\u2_Display/n1049 [16]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1033 ,\u2_Display/n1030 }),
    .f({\u2_Display/n1068 ,\u2_Display/n1065 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3354|_al_u3357  (
    .b({\u2_Display/n1049 [15],\u2_Display/n1049 [18]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1031 ,\u2_Display/n1028 }),
    .f({\u2_Display/n1066 ,\u2_Display/n1063 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3356|_al_u3359  (
    .b({\u2_Display/n1049 [17],\u2_Display/n1049 [20]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1029 ,\u2_Display/n1026 }),
    .f({\u2_Display/n1064 ,\u2_Display/n1061 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3358|_al_u3361  (
    .b({\u2_Display/n1049 [19],\u2_Display/n1049 [22]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1027 ,\u2_Display/n1024 }),
    .f({\u2_Display/n1062 ,\u2_Display/n1059 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u335|_al_u336  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [4],\u2_Display/counta [5]}),
    .d({\u2_Display/n3788 [4],\u2_Display/n3788 [5]}),
    .f({\u2_Display/n3816 ,\u2_Display/n3815 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3360|_al_u3363  (
    .b({\u2_Display/n1049 [21],\u2_Display/n1049 [24]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1025 ,\u2_Display/n1022 }),
    .f({\u2_Display/n1060 ,\u2_Display/n1057 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3362|_al_u3365  (
    .b({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .c({\u2_Display/n1049 [23],\u2_Display/n1049 [26]}),
    .d({\u2_Display/n1023 ,\u2_Display/n1020 }),
    .f({\u2_Display/n1058 ,\u2_Display/n1055 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3364|_al_u3368  (
    .b({\u2_Display/n1049 [25],\u2_Display/n1049 [29]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1021 ,\u2_Display/n1017 }),
    .f({\u2_Display/n1056 ,\u2_Display/n1052 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3366|_al_u3370  (
    .b({\u2_Display/n1049 [27],\u2_Display/n1049 [31]}),
    .c({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .d({\u2_Display/n1019 ,\u2_Display/n1015 }),
    .f({\u2_Display/n1054 ,\u2_Display/n1050 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    //.LUTF1("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUTG0("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    //.LUTG1("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT_LUTF0(16'b1110111001000100),
    .INIT_LUTF1(16'b1110010011100100),
    .INIT_LUTG0(16'b1110111001000100),
    .INIT_LUTG1(16'b1110010011100100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3367|_al_u3369  (
    .a({\u2_Display/n1047 ,\u2_Display/n1047 }),
    .b({\u2_Display/n1049 [28],\u2_Display/n1049 [30]}),
    .c({\u2_Display/n1018 ,open_n30395}),
    .d({open_n30398,\u2_Display/n1016 }),
    .f({\u2_Display/n1053 ,\u2_Display/n1051 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3372|_al_u3373  (
    .b({\u2_Display/n2172 [1],\u2_Display/n2172 [2]}),
    .c({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2168 ,\u2_Display/n2167 }),
    .f({\u2_Display/n2203 ,\u2_Display/n2202 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3374|_al_u3375  (
    .b({\u2_Display/n2172 [3],\u2_Display/n2172 [4]}),
    .c({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2166 ,\u2_Display/n2165 }),
    .f({\u2_Display/n2201 ,\u2_Display/n2200 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3376|_al_u3377  (
    .b({\u2_Display/n2172 [5],\u2_Display/n2172 [6]}),
    .c({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2164 ,\u2_Display/n2163 }),
    .f({\u2_Display/n2199 ,\u2_Display/n2198 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3378|_al_u3381  (
    .b({\u2_Display/n2172 [7],\u2_Display/n2172 [10]}),
    .c({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2162 ,\u2_Display/n2159 }),
    .f({\u2_Display/n2197 ,\u2_Display/n2194 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3380|_al_u3383  (
    .b({\u2_Display/n2172 [9],\u2_Display/n2172 [12]}),
    .c({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2160 ,\u2_Display/n2157 }),
    .f({\u2_Display/n2195 ,\u2_Display/n2192 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3382|_al_u3385  (
    .b({\u2_Display/n2172 [11],\u2_Display/n2172 [14]}),
    .c({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2158 ,\u2_Display/n2155 }),
    .f({\u2_Display/n2193 ,\u2_Display/n2190 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3384|_al_u3388  (
    .b({\u2_Display/n2172 [13],\u2_Display/n2172 [17]}),
    .c({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2156 ,\u2_Display/n2152 }),
    .f({\u2_Display/n2191 ,\u2_Display/n2187 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3386|_al_u3391  (
    .b({\u2_Display/n2172 [15],\u2_Display/n2172 [20]}),
    .c({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2154 ,\u2_Display/n2149 }),
    .f({\u2_Display/n2189 ,\u2_Display/n2184 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3387|_al_u3389  (
    .b({\u2_Display/n2172 [16],\u2_Display/n2172 [18]}),
    .c({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2153 ,\u2_Display/n2151 }),
    .f({\u2_Display/n2188 ,\u2_Display/n2186 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u338|_al_u340  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [7],\u2_Display/counta [9]}),
    .d({\u2_Display/n3788 [7],\u2_Display/n3788 [9]}),
    .f({\u2_Display/n3813 ,\u2_Display/n3811 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3390|_al_u3393  (
    .b({\u2_Display/n2172 [19],\u2_Display/n2172 [22]}),
    .c({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2150 ,\u2_Display/n2147 }),
    .f({\u2_Display/n2185 ,\u2_Display/n2182 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3392|_al_u3395  (
    .b({\u2_Display/n2172 [21],\u2_Display/n2172 [24]}),
    .c({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2148 ,\u2_Display/n2145 }),
    .f({\u2_Display/n2183 ,\u2_Display/n2180 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3394|_al_u3397  (
    .b({\u2_Display/n2172 [23],\u2_Display/n2172 [26]}),
    .c({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2146 ,\u2_Display/n2143 }),
    .f({\u2_Display/n2181 ,\u2_Display/n2178 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3396|_al_u3399  (
    .b({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .c({\u2_Display/n2172 [25],\u2_Display/n2172 [28]}),
    .d({\u2_Display/n2144 ,\u2_Display/n2141 }),
    .f({\u2_Display/n2179 ,\u2_Display/n2176 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    //.LUTF1("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    //.LUTG0("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    //.LUTG1("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    .INIT_LUTF0(16'b1101100011011000),
    .INIT_LUTF1(16'b1110111001000100),
    .INIT_LUTG0(16'b1101100011011000),
    .INIT_LUTG1(16'b1110111001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3398|_al_u3401  (
    .a({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .b({\u2_Display/n2172 [27],\u2_Display/n2139 }),
    .c({open_n30785,\u2_Display/n2172 [30]}),
    .d({\u2_Display/n2142 ,open_n30788}),
    .f({\u2_Display/n2177 ,\u2_Display/n2174 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3400|_al_u3402  (
    .b({\u2_Display/n2172 [29],\u2_Display/n2172 [31]}),
    .c({\u2_Display/n2170 ,\u2_Display/n2170 }),
    .d({\u2_Display/n2140 ,\u2_Display/n2138 }),
    .f({\u2_Display/n2175 ,\u2_Display/n2173 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3403|_al_u3405  (
    .b({\u2_Display/n3295 [0],\u2_Display/n3295 [2]}),
    .c({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3292 ,\u2_Display/n3290 }),
    .f({\u2_Display/n3327 ,\u2_Display/n3325 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3406|_al_u3407  (
    .b({\u2_Display/n3295 [3],\u2_Display/n3295 [4]}),
    .c({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3289 ,\u2_Display/n3288 }),
    .f({\u2_Display/n3324 ,\u2_Display/n3323 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3408|_al_u3409  (
    .b({\u2_Display/n3295 [5],\u2_Display/n3295 [6]}),
    .c({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3287 ,\u2_Display/n3286 }),
    .f({\u2_Display/n3322 ,\u2_Display/n3321 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3410|_al_u3413  (
    .b({\u2_Display/n3295 [7],\u2_Display/n3295 [10]}),
    .c({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3285 ,\u2_Display/n3282 }),
    .f({\u2_Display/n3320 ,\u2_Display/n3317 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3411|_al_u3412  (
    .b({\u2_Display/n3295 [8],\u2_Display/n3295 [9]}),
    .c({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3284 ,\u2_Display/n3283 }),
    .f({\u2_Display/n3319 ,\u2_Display/n3318 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3414|_al_u3419  (
    .b({\u2_Display/n3295 [11],\u2_Display/n3295 [16]}),
    .c({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3281 ,\u2_Display/n3276 }),
    .f({\u2_Display/n3316 ,\u2_Display/n3311 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3415|_al_u3417  (
    .b({\u2_Display/n3295 [12],\u2_Display/n3295 [14]}),
    .c({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3280 ,\u2_Display/n3278 }),
    .f({\u2_Display/n3315 ,\u2_Display/n3313 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3418|_al_u3421  (
    .b({\u2_Display/n3295 [15],\u2_Display/n3295 [18]}),
    .c({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3277 ,\u2_Display/n3274 }),
    .f({\u2_Display/n3312 ,\u2_Display/n3309 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u341|_al_u339  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .d({\u2_Display/n3788 [10],\u2_Display/n3788 [8]}),
    .f({\u2_Display/n3810 ,\u2_Display/n3812 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3420|_al_u3424  (
    .b({\u2_Display/n3295 [17],\u2_Display/n3295 [21]}),
    .c({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3275 ,\u2_Display/n3271 }),
    .f({\u2_Display/n3310 ,\u2_Display/n3306 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3422|_al_u3427  (
    .b({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .c({\u2_Display/n3295 [19],\u2_Display/n3295 [24]}),
    .d({\u2_Display/n3273 ,\u2_Display/n3268 }),
    .f({\u2_Display/n3308 ,\u2_Display/n3303 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3423|_al_u3425  (
    .b({\u2_Display/n3295 [20],\u2_Display/n3295 [22]}),
    .c({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3272 ,\u2_Display/n3270 }),
    .f({\u2_Display/n3307 ,\u2_Display/n3305 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTF1("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    //.LUTG0("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTG1("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT_LUTF0(16'b1111101001010000),
    .INIT_LUTF1(16'b1101100011011000),
    .INIT_LUTG0(16'b1111101001010000),
    .INIT_LUTG1(16'b1101100011011000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3426|_al_u3429  (
    .a({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .b({\u2_Display/n3269 ,open_n31149}),
    .c({\u2_Display/n3295 [23],\u2_Display/n3295 [26]}),
    .d({open_n31152,\u2_Display/n3266 }),
    .f({\u2_Display/n3304 ,\u2_Display/n3301 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3428|_al_u3431  (
    .b({\u2_Display/n3295 [25],\u2_Display/n3295 [28]}),
    .c({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3267 ,\u2_Display/n3264 }),
    .f({\u2_Display/n3302 ,\u2_Display/n3299 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u342|_al_u347  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [11],\u2_Display/counta [16]}),
    .d({\u2_Display/n3788 [11],\u2_Display/n3788 [16]}),
    .f({\u2_Display/n3809 ,\u2_Display/n3804 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3430|_al_u3433  (
    .b({\u2_Display/n3295 [27],\u2_Display/n3295 [30]}),
    .c({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3265 ,\u2_Display/n3262 }),
    .f({\u2_Display/n3300 ,\u2_Display/n3297 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3432|_al_u3434  (
    .b({\u2_Display/n3295 [29],\u2_Display/n3295 [31]}),
    .c({\u2_Display/n3293 ,\u2_Display/n3293 }),
    .d({\u2_Display/n3263 ,\u2_Display/n3261 }),
    .f({\u2_Display/n3298 ,\u2_Display/n3296 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3435|_al_u3437  (
    .b({\u2_Display/n4453 [0],\u2_Display/n4453 [2]}),
    .c({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .d({\u2_Display/n4450 ,\u2_Display/n4448 }),
    .f({\u2_Display/n4485 ,\u2_Display/n4483 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u3436 (
    .b({open_n31307,\u2_Display/n4453 [1]}),
    .c({open_n31308,\u2_Display/n4451 }),
    .d({open_n31311,\u2_Display/n4449 }),
    .f({open_n31329,\u2_Display/n4484 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3438|_al_u3439  (
    .b({\u2_Display/n4453 [3],\u2_Display/n4453 [4]}),
    .c({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .d({\u2_Display/n4447 ,\u2_Display/n4446 }),
    .f({\u2_Display/n4482 ,\u2_Display/n4481 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u343|_al_u345  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [12],\u2_Display/counta [14]}),
    .d({\u2_Display/n3788 [12],\u2_Display/n3788 [14]}),
    .f({\u2_Display/n3808 ,\u2_Display/n3806 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u344 (
    .b({open_n31389,\u2_Display/n3786 }),
    .c({open_n31390,\u2_Display/counta [13]}),
    .d({open_n31393,\u2_Display/n3788 [13]}),
    .f({open_n31411,\u2_Display/n3807 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3440|_al_u3441  (
    .b({\u2_Display/n4453 [5],\u2_Display/n4453 [6]}),
    .c({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .d({\u2_Display/n4445 ,\u2_Display/n4444 }),
    .f({\u2_Display/n4480 ,\u2_Display/n4479 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3442|_al_u3443  (
    .b({\u2_Display/n4453 [7],\u2_Display/n4453 [8]}),
    .c({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .d({\u2_Display/n4443 ,\u2_Display/n4442 }),
    .f({\u2_Display/n4478 ,\u2_Display/n4477 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3444|_al_u3445  (
    .b({\u2_Display/n4453 [9],\u2_Display/n4453 [10]}),
    .c({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .d({\u2_Display/n4441 ,\u2_Display/n4440 }),
    .f({\u2_Display/n4476 ,\u2_Display/n4475 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3446|_al_u3447  (
    .b({\u2_Display/n4453 [11],\u2_Display/n4453 [12]}),
    .c({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .d({\u2_Display/n4439 ,\u2_Display/n4438 }),
    .f({\u2_Display/n4474 ,\u2_Display/n4473 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3448|_al_u3449  (
    .b({\u2_Display/n4453 [13],\u2_Display/n4453 [14]}),
    .c({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .d({\u2_Display/n4437 ,\u2_Display/n4436 }),
    .f({\u2_Display/n4472 ,\u2_Display/n4471 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3450|_al_u3453  (
    .b({\u2_Display/n4453 [15],\u2_Display/n4453 [18]}),
    .c({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .d({\u2_Display/n4435 ,\u2_Display/n4432 }),
    .f({\u2_Display/n4470 ,\u2_Display/n4467 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u3451 (
    .b({open_n31575,\u2_Display/n4453 [16]}),
    .c({open_n31576,\u2_Display/n4451 }),
    .d({open_n31579,\u2_Display/n4434 }),
    .f({open_n31597,\u2_Display/n4469 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3452|_al_u3455  (
    .b({\u2_Display/n4453 [17],\u2_Display/n4453 [20]}),
    .c({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .d({\u2_Display/n4433 ,\u2_Display/n4430 }),
    .f({\u2_Display/n4468 ,\u2_Display/n4465 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3454|_al_u3457  (
    .b({\u2_Display/n4453 [19],\u2_Display/n4453 [22]}),
    .c({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .d({\u2_Display/n4431 ,\u2_Display/n4428 }),
    .f({\u2_Display/n4466 ,\u2_Display/n4463 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3456|_al_u3460  (
    .b({\u2_Display/n4453 [21],\u2_Display/n4453 [25]}),
    .c({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .d({\u2_Display/n4429 ,\u2_Display/n4425 }),
    .f({\u2_Display/n4464 ,\u2_Display/n4460 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3458|_al_u3464  (
    .b({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .c({\u2_Display/n4453 [23],\u2_Display/n4453 [29]}),
    .d({\u2_Display/n4427 ,\u2_Display/n4421 }),
    .f({\u2_Display/n4462 ,\u2_Display/n4456 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3459|_al_u3461  (
    .b({\u2_Display/n4453 [24],\u2_Display/n4453 [26]}),
    .c({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .d({\u2_Display/n4426 ,\u2_Display/n4424 }),
    .f({\u2_Display/n4461 ,\u2_Display/n4459 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUTF1("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTG0("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUTG1("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    .INIT_LUTF0(16'b1110010011100100),
    .INIT_LUTF1(16'b1111101001010000),
    .INIT_LUTG0(16'b1110010011100100),
    .INIT_LUTG1(16'b1111101001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3462|_al_u3466  (
    .a({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .b({open_n31733,\u2_Display/n4453 [31]}),
    .c({\u2_Display/n4453 [27],\u2_Display/n4419 }),
    .d({\u2_Display/n4423 ,open_n31736}),
    .f({\u2_Display/n4458 ,\u2_Display/n4454 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3463|_al_u3465  (
    .b({\u2_Display/n4453 [28],\u2_Display/n4453 [30]}),
    .c({\u2_Display/n4451 ,\u2_Display/n4451 }),
    .d({\u2_Display/n4422 ,\u2_Display/n4420 }),
    .f({\u2_Display/n4457 ,\u2_Display/n4455 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3467|_al_u3472  (
    .b({\u2_Display/n5576 [0],\u2_Display/n5576 [5]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5573 ,\u2_Display/n5568 }),
    .f({\u2_Display/n5608 ,\u2_Display/n5603 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3468|_al_u3469  (
    .b({\u2_Display/n5576 [1],\u2_Display/n5576 [2]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5572 ,\u2_Display/n5571 }),
    .f({\u2_Display/n5607 ,\u2_Display/n5606 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u346|_al_u349  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [15],\u2_Display/counta [18]}),
    .d({\u2_Display/n3788 [15],\u2_Display/n3788 [18]}),
    .f({\u2_Display/n3805 ,\u2_Display/n3802 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3470|_al_u3476  (
    .b({\u2_Display/n5576 [3],\u2_Display/n5576 [9]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5570 ,\u2_Display/n5564 }),
    .f({\u2_Display/n5605 ,\u2_Display/n5599 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3471|_al_u3473  (
    .b({\u2_Display/n5576 [4],\u2_Display/n5576 [6]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5569 ,\u2_Display/n5567 }),
    .f({\u2_Display/n5604 ,\u2_Display/n5602 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3474|_al_u3480  (
    .b({\u2_Display/n5576 [7],\u2_Display/n5576 [13]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5566 ,\u2_Display/n5560 }),
    .f({\u2_Display/n5601 ,\u2_Display/n5595 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3475|_al_u3477  (
    .b({\u2_Display/n5576 [8],\u2_Display/n5576 [10]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5565 ,\u2_Display/n5563 }),
    .f({\u2_Display/n5600 ,\u2_Display/n5598 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3478|_al_u3484  (
    .b({\u2_Display/n5576 [11],\u2_Display/n5576 [17]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5562 ,\u2_Display/n5556 }),
    .f({\u2_Display/n5597 ,\u2_Display/n5591 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3479|_al_u3481  (
    .b({\u2_Display/n5576 [12],\u2_Display/n5576 [14]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5561 ,\u2_Display/n5559 }),
    .f({\u2_Display/n5596 ,\u2_Display/n5594 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3482|_al_u3487  (
    .b({\u2_Display/n5576 [15],\u2_Display/n5576 [20]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5558 ,\u2_Display/n5553 }),
    .f({\u2_Display/n5593 ,\u2_Display/n5588 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3483|_al_u3485  (
    .b({\u2_Display/n5576 [16],\u2_Display/n5576 [18]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5557 ,\u2_Display/n5555 }),
    .f({\u2_Display/n5592 ,\u2_Display/n5590 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3486|_al_u3489  (
    .b({\u2_Display/n5576 [19],\u2_Display/n5576 [22]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5554 ,\u2_Display/n5551 }),
    .f({\u2_Display/n5589 ,\u2_Display/n5586 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3488|_al_u3492  (
    .b({\u2_Display/n5576 [21],\u2_Display/n5576 [25]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5552 ,\u2_Display/n5548 }),
    .f({\u2_Display/n5587 ,\u2_Display/n5583 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u348|_al_u351  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [17],\u2_Display/counta [20]}),
    .d({\u2_Display/n3788 [17],\u2_Display/n3788 [20]}),
    .f({\u2_Display/n3803 ,\u2_Display/n3800 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3490|_al_u3495  (
    .b({\u2_Display/n5576 [23],\u2_Display/n5576 [28]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5550 ,\u2_Display/n5545 }),
    .f({\u2_Display/n5585 ,\u2_Display/n5580 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3491|_al_u3493  (
    .b({\u2_Display/n5576 [24],\u2_Display/n5576 [26]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5549 ,\u2_Display/n5547 }),
    .f({\u2_Display/n5584 ,\u2_Display/n5582 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3494|_al_u3497  (
    .b({\u2_Display/n5576 [27],\u2_Display/n5576 [30]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5546 ,\u2_Display/n5543 }),
    .f({\u2_Display/n5581 ,\u2_Display/n5578 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3496|_al_u3498  (
    .b({\u2_Display/n5576 [29],\u2_Display/n5576 [31]}),
    .c({\u2_Display/n5574 ,\u2_Display/n5574 }),
    .d({\u2_Display/n5544 ,\u2_Display/n5542 }),
    .f({\u2_Display/n5579 ,\u2_Display/n5577 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3499|_al_u3503  (
    .b({\u2_Display/n1084 [0],\u2_Display/n1084 [4]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1081 ,\u2_Display/n1077 }),
    .f({\u2_Display/n1116 ,\u2_Display/n1112 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3500|_al_u3501  (
    .b({\u2_Display/n1084 [1],\u2_Display/n1084 [2]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1080 ,\u2_Display/n1079 }),
    .f({\u2_Display/n1115 ,\u2_Display/n1114 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3502|_al_u3505  (
    .b({\u2_Display/n1084 [3],\u2_Display/n1084 [6]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1078 ,\u2_Display/n1075 }),
    .f({\u2_Display/n1113 ,\u2_Display/n1110 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3504|_al_u3507  (
    .b({\u2_Display/n1084 [5],\u2_Display/n1084 [8]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1076 ,\u2_Display/n1073 }),
    .f({\u2_Display/n1111 ,\u2_Display/n1108 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3506|_al_u3509  (
    .b({\u2_Display/n1084 [7],\u2_Display/n1084 [10]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1074 ,\u2_Display/n1071 }),
    .f({\u2_Display/n1109 ,\u2_Display/n1106 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3508|_al_u3511  (
    .b({\u2_Display/n1084 [9],\u2_Display/n1084 [12]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1072 ,\u2_Display/n1069 }),
    .f({\u2_Display/n1107 ,\u2_Display/n1104 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u350|_al_u353  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [19],\u2_Display/counta [22]}),
    .d({\u2_Display/n3788 [19],\u2_Display/n3788 [22]}),
    .f({\u2_Display/n3801 ,\u2_Display/n3798 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3510|_al_u3513  (
    .b({\u2_Display/n1084 [11],\u2_Display/n1084 [14]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1070 ,\u2_Display/n1067 }),
    .f({\u2_Display/n1105 ,\u2_Display/n1102 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3512|_al_u3515  (
    .b({\u2_Display/n1084 [13],\u2_Display/n1084 [16]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1068 ,\u2_Display/n1065 }),
    .f({\u2_Display/n1103 ,\u2_Display/n1100 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3514|_al_u3517  (
    .b({\u2_Display/n1084 [15],\u2_Display/n1084 [18]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1066 ,\u2_Display/n1063 }),
    .f({\u2_Display/n1101 ,\u2_Display/n1098 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3516|_al_u3519  (
    .b({\u2_Display/n1084 [17],\u2_Display/n1084 [20]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1064 ,\u2_Display/n1061 }),
    .f({\u2_Display/n1099 ,\u2_Display/n1096 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3518|_al_u3521  (
    .b({\u2_Display/n1084 [19],\u2_Display/n1084 [22]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1062 ,\u2_Display/n1059 }),
    .f({\u2_Display/n1097 ,\u2_Display/n1094 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3520|_al_u3523  (
    .b({\u2_Display/n1084 [21],\u2_Display/n1084 [24]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1060 ,\u2_Display/n1057 }),
    .f({\u2_Display/n1095 ,\u2_Display/n1092 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3522|_al_u3525  (
    .b({\u2_Display/n1084 [23],\u2_Display/n1084 [26]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1058 ,\u2_Display/n1055 }),
    .f({\u2_Display/n1093 ,\u2_Display/n1090 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3524|_al_u3527  (
    .b({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .c({\u2_Display/n1084 [25],\u2_Display/n1084 [28]}),
    .d({\u2_Display/n1056 ,\u2_Display/n1053 }),
    .f({\u2_Display/n1091 ,\u2_Display/n1088 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3526|_al_u3529  (
    .b({\u2_Display/n1084 [27],\u2_Display/n1084 [30]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1054 ,\u2_Display/n1051 }),
    .f({\u2_Display/n1089 ,\u2_Display/n1086 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3528|_al_u3530  (
    .b({\u2_Display/n1084 [29],\u2_Display/n1084 [31]}),
    .c({\u2_Display/n1082 ,\u2_Display/n1082 }),
    .d({\u2_Display/n1052 ,\u2_Display/n1050 }),
    .f({\u2_Display/n1087 ,\u2_Display/n1085 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u352|_al_u355  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [21],\u2_Display/counta [24]}),
    .d({\u2_Display/n3788 [21],\u2_Display/n3788 [24]}),
    .f({\u2_Display/n3799 ,\u2_Display/n3796 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3531|_al_u3533  (
    .b({\u2_Display/n2207 [0],\u2_Display/n2207 [2]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2204 ,\u2_Display/n2202 }),
    .f({\u2_Display/n2239 ,\u2_Display/n2237 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3532|_al_u3536  (
    .b({\u2_Display/n2207 [1],\u2_Display/n2207 [5]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2203 ,\u2_Display/n2199 }),
    .f({\u2_Display/n2238 ,\u2_Display/n2234 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3534|_al_u3539  (
    .b({\u2_Display/n2207 [3],\u2_Display/n2207 [8]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2201 ,\u2_Display/n2196 }),
    .f({\u2_Display/n2236 ,\u2_Display/n2231 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3535|_al_u3537  (
    .b({\u2_Display/n2207 [4],\u2_Display/n2207 [6]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2200 ,\u2_Display/n2198 }),
    .f({\u2_Display/n2235 ,\u2_Display/n2233 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3538|_al_u3541  (
    .b({\u2_Display/n2207 [7],\u2_Display/n2207 [10]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2197 ,\u2_Display/n2194 }),
    .f({\u2_Display/n2232 ,\u2_Display/n2229 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3540|_al_u3543  (
    .b({\u2_Display/n2207 [9],\u2_Display/n2207 [12]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2195 ,\u2_Display/n2192 }),
    .f({\u2_Display/n2230 ,\u2_Display/n2227 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3542|_al_u3545  (
    .b({\u2_Display/n2207 [11],\u2_Display/n2207 [14]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2193 ,\u2_Display/n2190 }),
    .f({\u2_Display/n2228 ,\u2_Display/n2225 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3544|_al_u3548  (
    .b({\u2_Display/n2207 [13],\u2_Display/n2207 [17]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2191 ,\u2_Display/n2187 }),
    .f({\u2_Display/n2226 ,\u2_Display/n2222 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3546|_al_u3552  (
    .b({\u2_Display/n2207 [15],\u2_Display/n2207 [21]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2189 ,\u2_Display/n2183 }),
    .f({\u2_Display/n2224 ,\u2_Display/n2218 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3547|_al_u3549  (
    .b({\u2_Display/n2207 [16],\u2_Display/n2207 [18]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2188 ,\u2_Display/n2186 }),
    .f({\u2_Display/n2223 ,\u2_Display/n2221 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u354|_al_u357  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [23],\u2_Display/counta [26]}),
    .d({\u2_Display/n3788 [23],\u2_Display/n3788 [26]}),
    .f({\u2_Display/n3797 ,\u2_Display/n3794 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3550|_al_u3555  (
    .b({\u2_Display/n2207 [19],\u2_Display/n2207 [24]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2185 ,\u2_Display/n2180 }),
    .f({\u2_Display/n2220 ,\u2_Display/n2215 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3551|_al_u3553  (
    .b({\u2_Display/n2207 [20],\u2_Display/n2207 [22]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2184 ,\u2_Display/n2182 }),
    .f({\u2_Display/n2219 ,\u2_Display/n2217 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3554|_al_u3557  (
    .b({\u2_Display/n2207 [23],\u2_Display/n2207 [26]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2181 ,\u2_Display/n2178 }),
    .f({\u2_Display/n2216 ,\u2_Display/n2213 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3556|_al_u3559  (
    .b({\u2_Display/n2207 [25],\u2_Display/n2207 [28]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2179 ,\u2_Display/n2176 }),
    .f({\u2_Display/n2214 ,\u2_Display/n2211 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3558|_al_u3561  (
    .b({\u2_Display/n2207 [27],\u2_Display/n2207 [30]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2177 ,\u2_Display/n2174 }),
    .f({\u2_Display/n2212 ,\u2_Display/n2209 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3560|_al_u3562  (
    .b({\u2_Display/n2207 [29],\u2_Display/n2207 [31]}),
    .c({\u2_Display/n2205 ,\u2_Display/n2205 }),
    .d({\u2_Display/n2175 ,\u2_Display/n2173 }),
    .f({\u2_Display/n2210 ,\u2_Display/n2208 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3563|_al_u3565  (
    .b({\u2_Display/n3330 [0],\u2_Display/n3330 [2]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .d({\u2_Display/n3327 ,\u2_Display/n3325 }),
    .f({\u2_Display/n3362 ,\u2_Display/n3360 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3564|_al_u3567  (
    .b({\u2_Display/n3330 [1],\u2_Display/n3330 [4]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .d({\u2_Display/n3326 ,\u2_Display/n3323 }),
    .f({\u2_Display/n3361 ,\u2_Display/n3358 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3566|_al_u3569  (
    .b({\u2_Display/n3330 [3],\u2_Display/n3330 [6]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .d({\u2_Display/n3324 ,\u2_Display/n3321 }),
    .f({\u2_Display/n3359 ,\u2_Display/n3356 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3568|_al_u3572  (
    .b({\u2_Display/n3330 [5],\u2_Display/n3330 [9]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .d({\u2_Display/n3322 ,\u2_Display/n3318 }),
    .f({\u2_Display/n3357 ,\u2_Display/n3353 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u356|_al_u360  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [25],\u2_Display/counta [29]}),
    .d({\u2_Display/n3788 [25],\u2_Display/n3788 [29]}),
    .f({\u2_Display/n3795 ,\u2_Display/n3791 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3570|_al_u3575  (
    .b({\u2_Display/n3330 [7],\u2_Display/n3330 [12]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .d({\u2_Display/n3320 ,\u2_Display/n3315 }),
    .f({\u2_Display/n3355 ,\u2_Display/n3350 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3571|_al_u3573  (
    .b({\u2_Display/n3330 [8],\u2_Display/n3330 [10]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .d({\u2_Display/n3319 ,\u2_Display/n3317 }),
    .f({\u2_Display/n3354 ,\u2_Display/n3352 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3574|_al_u3577  (
    .b({\u2_Display/n3330 [11],\u2_Display/n3330 [14]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .d({\u2_Display/n3316 ,\u2_Display/n3313 }),
    .f({\u2_Display/n3351 ,\u2_Display/n3348 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3576|_al_u3579  (
    .b({\u2_Display/n3330 [13],\u2_Display/n3330 [16]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .d({\u2_Display/n3314 ,\u2_Display/n3311 }),
    .f({\u2_Display/n3349 ,\u2_Display/n3346 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3578|_al_u3581  (
    .b({\u2_Display/n3330 [15],\u2_Display/n3330 [18]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .d({\u2_Display/n3312 ,\u2_Display/n3309 }),
    .f({\u2_Display/n3347 ,\u2_Display/n3344 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3580|_al_u3583  (
    .b({\u2_Display/n3330 [17],\u2_Display/n3330 [20]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .d({\u2_Display/n3310 ,\u2_Display/n3307 }),
    .f({\u2_Display/n3345 ,\u2_Display/n3342 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3582|_al_u3585  (
    .b({\u2_Display/n3330 [19],\u2_Display/n3330 [22]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .d({\u2_Display/n3308 ,\u2_Display/n3305 }),
    .f({\u2_Display/n3343 ,\u2_Display/n3340 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3584|_al_u3588  (
    .b({\u2_Display/n3330 [21],\u2_Display/n3330 [25]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .d({\u2_Display/n3306 ,\u2_Display/n3302 }),
    .f({\u2_Display/n3341 ,\u2_Display/n3337 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3586|_al_u3723  (
    .b({\u2_Display/n3330 [23],\u2_Display/n3365 [0]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3304 ,\u2_Display/n3362 }),
    .f({\u2_Display/n3339 ,\u2_Display/n3397 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3587|_al_u3589  (
    .b({\u2_Display/n3330 [24],\u2_Display/n3330 [26]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .d({\u2_Display/n3303 ,\u2_Display/n3301 }),
    .f({\u2_Display/n3338 ,\u2_Display/n3336 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u358|_al_u362  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [27],\u2_Display/counta [31]}),
    .d({\u2_Display/n3788 [27],\u2_Display/n3788 [31]}),
    .f({\u2_Display/n3793 ,\u2_Display/n3789 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3590|_al_u3593  (
    .b({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .c({\u2_Display/n3330 [27],\u2_Display/n3330 [30]}),
    .d({\u2_Display/n3300 ,\u2_Display/n3297 }),
    .f({\u2_Display/n3335 ,\u2_Display/n3332 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUTF1("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTG0("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUTG1("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    .INIT_LUTF0(16'b1110010011100100),
    .INIT_LUTF1(16'b1111101001010000),
    .INIT_LUTG0(16'b1110010011100100),
    .INIT_LUTG1(16'b1111101001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3591|_al_u3592  (
    .a({\u2_Display/n3328 ,\u2_Display/n3328 }),
    .b({open_n33605,\u2_Display/n3330 [29]}),
    .c({\u2_Display/n3330 [28],\u2_Display/n3298 }),
    .d({\u2_Display/n3299 ,open_n33608}),
    .f({\u2_Display/n3334 ,\u2_Display/n3333 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3594|_al_u3731  (
    .b({\u2_Display/n3330 [31],\u2_Display/n3365 [8]}),
    .c({\u2_Display/n3328 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3296 ,\u2_Display/n3354 }),
    .f({\u2_Display/n3331 ,\u2_Display/n3389 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3595|_al_u3599  (
    .b({\u2_Display/n4488 [0],\u2_Display/n4488 [4]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4485 ,\u2_Display/n4481 }),
    .f({\u2_Display/n4520 ,\u2_Display/n4516 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3596|_al_u3597  (
    .b({\u2_Display/n4488 [1],\u2_Display/n4488 [2]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4484 ,\u2_Display/n4483 }),
    .f({\u2_Display/n4519 ,\u2_Display/n4518 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3598|_al_u3601  (
    .b({\u2_Display/n4488 [3],\u2_Display/n4488 [6]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4482 ,\u2_Display/n4479 }),
    .f({\u2_Display/n4517 ,\u2_Display/n4514 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u359|_al_u361  (
    .b({\u2_Display/n3786 ,\u2_Display/n3786 }),
    .c({\u2_Display/counta [28],\u2_Display/counta [30]}),
    .d({\u2_Display/n3788 [28],\u2_Display/n3788 [30]}),
    .f({\u2_Display/n3792 ,\u2_Display/n3790 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3600|_al_u3603  (
    .b({\u2_Display/n4488 [5],\u2_Display/n4488 [8]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4480 ,\u2_Display/n4477 }),
    .f({\u2_Display/n4515 ,\u2_Display/n4512 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3602|_al_u3604  (
    .b({\u2_Display/n4488 [7],\u2_Display/n4488 [9]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4478 ,\u2_Display/n4476 }),
    .f({\u2_Display/n4513 ,\u2_Display/n4511 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3605|_al_u3607  (
    .b({\u2_Display/n4488 [10],\u2_Display/n4488 [12]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4475 ,\u2_Display/n4473 }),
    .f({\u2_Display/n4510 ,\u2_Display/n4508 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3606|_al_u3609  (
    .b({\u2_Display/n4488 [11],\u2_Display/n4488 [14]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4474 ,\u2_Display/n4471 }),
    .f({\u2_Display/n4509 ,\u2_Display/n4506 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3608|_al_u3612  (
    .b({\u2_Display/n4488 [13],\u2_Display/n4488 [17]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4472 ,\u2_Display/n4468 }),
    .f({\u2_Display/n4507 ,\u2_Display/n4503 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3610|_al_u3615  (
    .b({\u2_Display/n4488 [15],\u2_Display/n4488 [20]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4470 ,\u2_Display/n4465 }),
    .f({\u2_Display/n4505 ,\u2_Display/n4500 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3611|_al_u3613  (
    .b({\u2_Display/n4488 [16],\u2_Display/n4488 [18]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4469 ,\u2_Display/n4467 }),
    .f({\u2_Display/n4504 ,\u2_Display/n4502 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3614|_al_u3617  (
    .b({\u2_Display/n4488 [19],\u2_Display/n4488 [22]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4466 ,\u2_Display/n4463 }),
    .f({\u2_Display/n4501 ,\u2_Display/n4498 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3616|_al_u3619  (
    .b({\u2_Display/n4488 [21],\u2_Display/n4488 [24]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4464 ,\u2_Display/n4461 }),
    .f({\u2_Display/n4499 ,\u2_Display/n4496 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3618|_al_u3621  (
    .b({\u2_Display/n4488 [23],\u2_Display/n4488 [26]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4462 ,\u2_Display/n4459 }),
    .f({\u2_Display/n4497 ,\u2_Display/n4494 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3620|_al_u3623  (
    .b({\u2_Display/n4488 [25],\u2_Display/n4488 [28]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4460 ,\u2_Display/n4457 }),
    .f({\u2_Display/n4495 ,\u2_Display/n4492 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3622|_al_u3625  (
    .b({\u2_Display/n4488 [27],\u2_Display/n4488 [30]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4458 ,\u2_Display/n4455 }),
    .f({\u2_Display/n4493 ,\u2_Display/n4490 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3624|_al_u3626  (
    .b({\u2_Display/n4488 [29],\u2_Display/n4488 [31]}),
    .c({\u2_Display/n4486 ,\u2_Display/n4486 }),
    .d({\u2_Display/n4456 ,\u2_Display/n4454 }),
    .f({\u2_Display/n4491 ,\u2_Display/n4489 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3627|_al_u3632  (
    .b({\u2_Display/n5611 [0],\u2_Display/n5611 [5]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5608 ,\u2_Display/n5603 }),
    .f({\u2_Display/n5643 ,\u2_Display/n5638 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3628|_al_u3629  (
    .b({\u2_Display/n5611 [1],\u2_Display/n5611 [2]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5607 ,\u2_Display/n5606 }),
    .f({\u2_Display/n5642 ,\u2_Display/n5641 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3630|_al_u3635  (
    .b({\u2_Display/n5611 [3],\u2_Display/n5611 [8]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5605 ,\u2_Display/n5600 }),
    .f({\u2_Display/n5640 ,\u2_Display/n5635 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3631|_al_u3633  (
    .b({\u2_Display/n5611 [4],\u2_Display/n5611 [6]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5604 ,\u2_Display/n5602 }),
    .f({\u2_Display/n5639 ,\u2_Display/n5637 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3634|_al_u3637  (
    .b({\u2_Display/n5611 [7],\u2_Display/n5611 [10]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5601 ,\u2_Display/n5598 }),
    .f({\u2_Display/n5636 ,\u2_Display/n5633 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3636|_al_u3639  (
    .b({\u2_Display/n5611 [9],\u2_Display/n5611 [12]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5599 ,\u2_Display/n5596 }),
    .f({\u2_Display/n5634 ,\u2_Display/n5631 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3638|_al_u3641  (
    .b({\u2_Display/n5611 [11],\u2_Display/n5611 [14]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5597 ,\u2_Display/n5594 }),
    .f({\u2_Display/n5632 ,\u2_Display/n5629 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u363|_al_u365  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [0],\u2_Display/counta [2]}),
    .d({\u2_Display/n4911 [0],\u2_Display/n4911 [2]}),
    .f({\u2_Display/n6101 ,\u2_Display/n6099 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u364 (
    .b({open_n34309,\u2_Display/n4909 }),
    .c({open_n34310,\u2_Display/counta [1]}),
    .d({open_n34313,\u2_Display/n4911 [1]}),
    .f({open_n34331,\u2_Display/n6100 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3640|_al_u3643  (
    .b({\u2_Display/n5611 [13],\u2_Display/n5611 [16]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5595 ,\u2_Display/n5592 }),
    .f({\u2_Display/n5630 ,\u2_Display/n5627 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3642|_al_u3645  (
    .b({\u2_Display/n5611 [15],\u2_Display/n5611 [18]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5593 ,\u2_Display/n5590 }),
    .f({\u2_Display/n5628 ,\u2_Display/n5625 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3644|_al_u3647  (
    .b({\u2_Display/n5611 [17],\u2_Display/n5611 [20]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5591 ,\u2_Display/n5588 }),
    .f({\u2_Display/n5626 ,\u2_Display/n5623 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3646|_al_u3649  (
    .b({\u2_Display/n5611 [19],\u2_Display/n5611 [22]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5589 ,\u2_Display/n5586 }),
    .f({\u2_Display/n5624 ,\u2_Display/n5621 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3648|_al_u3652  (
    .b({\u2_Display/n5611 [21],\u2_Display/n5611 [25]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5587 ,\u2_Display/n5583 }),
    .f({\u2_Display/n5622 ,\u2_Display/n5618 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3650|_al_u3656  (
    .b({\u2_Display/n5611 [23],\u2_Display/n5611 [29]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5585 ,\u2_Display/n5579 }),
    .f({\u2_Display/n5620 ,\u2_Display/n5614 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3651|_al_u3653  (
    .b({\u2_Display/n5611 [24],\u2_Display/n5611 [26]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5584 ,\u2_Display/n5582 }),
    .f({\u2_Display/n5619 ,\u2_Display/n5617 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3654|_al_u3658  (
    .b({\u2_Display/n5611 [27],\u2_Display/n5609 }),
    .c({\u2_Display/n5609 ,\u2_Display/n5611 [31]}),
    .d({\u2_Display/n5581 ,\u2_Display/n5577 }),
    .f({\u2_Display/n5616 ,\u2_Display/n5612 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3655|_al_u3657  (
    .b({\u2_Display/n5611 [28],\u2_Display/n5611 [30]}),
    .c({\u2_Display/n5609 ,\u2_Display/n5609 }),
    .d({\u2_Display/n5580 ,\u2_Display/n5578 }),
    .f({\u2_Display/n5615 ,\u2_Display/n5613 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3659|_al_u3663  (
    .b({\u2_Display/n1119 [0],\u2_Display/n1119 [4]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1116 ,\u2_Display/n1112 }),
    .f({\u2_Display/n1151 ,\u2_Display/n1147 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3660|_al_u3661  (
    .b({\u2_Display/n1119 [1],\u2_Display/n1119 [2]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1115 ,\u2_Display/n1114 }),
    .f({\u2_Display/n1150 ,\u2_Display/n1149 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3662|_al_u3665  (
    .b({\u2_Display/n1119 [3],\u2_Display/n1119 [6]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1113 ,\u2_Display/n1110 }),
    .f({\u2_Display/n1148 ,\u2_Display/n1145 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3664|_al_u3667  (
    .b({\u2_Display/n1119 [5],\u2_Display/n1119 [8]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1111 ,\u2_Display/n1108 }),
    .f({\u2_Display/n1146 ,\u2_Display/n1143 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3666|_al_u3669  (
    .b({\u2_Display/n1119 [7],\u2_Display/n1119 [10]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1109 ,\u2_Display/n1106 }),
    .f({\u2_Display/n1144 ,\u2_Display/n1141 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3668|_al_u3671  (
    .b({\u2_Display/n1119 [9],\u2_Display/n1119 [12]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1107 ,\u2_Display/n1104 }),
    .f({\u2_Display/n1142 ,\u2_Display/n1139 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u366|_al_u367  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [3],\u2_Display/counta [4]}),
    .d({\u2_Display/n4911 [3],\u2_Display/n4911 [4]}),
    .f({\u2_Display/n6098 ,\u2_Display/n6097 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3670|_al_u3673  (
    .b({\u2_Display/n1119 [11],\u2_Display/n1119 [14]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1105 ,\u2_Display/n1102 }),
    .f({\u2_Display/n1140 ,\u2_Display/n1137 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3672|_al_u3676  (
    .b({\u2_Display/n1119 [13],\u2_Display/n1119 [17]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1103 ,\u2_Display/n1099 }),
    .f({\u2_Display/n1138 ,\u2_Display/n1134 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3674|_al_u3680  (
    .b({\u2_Display/n1119 [15],\u2_Display/n1119 [21]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1101 ,\u2_Display/n1095 }),
    .f({\u2_Display/n1136 ,\u2_Display/n1130 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3675|_al_u3677  (
    .b({\u2_Display/n1119 [16],\u2_Display/n1119 [18]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1100 ,\u2_Display/n1098 }),
    .f({\u2_Display/n1135 ,\u2_Display/n1133 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUTF1("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTG0("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUTG1("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    .INIT_LUTF0(16'b1110010011100100),
    .INIT_LUTF1(16'b1111101001010000),
    .INIT_LUTG0(16'b1110010011100100),
    .INIT_LUTG1(16'b1111101001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3678|_al_u3683  (
    .a({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .b({open_n34857,\u2_Display/n1119 [24]}),
    .c({\u2_Display/n1119 [19],\u2_Display/n1092 }),
    .d({\u2_Display/n1097 ,open_n34860}),
    .f({\u2_Display/n1132 ,\u2_Display/n1127 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3679|_al_u3681  (
    .b({\u2_Display/n1119 [20],\u2_Display/n1119 [22]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1096 ,\u2_Display/n1094 }),
    .f({\u2_Display/n1131 ,\u2_Display/n1129 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3682|_al_u3685  (
    .b({\u2_Display/n1119 [23],\u2_Display/n1119 [26]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1093 ,\u2_Display/n1090 }),
    .f({\u2_Display/n1128 ,\u2_Display/n1125 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3684|_al_u3687  (
    .b({\u2_Display/n1119 [25],\u2_Display/n1119 [28]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1091 ,\u2_Display/n1088 }),
    .f({\u2_Display/n1126 ,\u2_Display/n1123 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3686|_al_u3689  (
    .b({\u2_Display/n1119 [27],\u2_Display/n1119 [30]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1089 ,\u2_Display/n1086 }),
    .f({\u2_Display/n1124 ,\u2_Display/n1121 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3688|_al_u3690  (
    .b({\u2_Display/n1119 [29],\u2_Display/n1119 [31]}),
    .c({\u2_Display/n1117 ,\u2_Display/n1117 }),
    .d({\u2_Display/n1087 ,\u2_Display/n1085 }),
    .f({\u2_Display/n1122 ,\u2_Display/n1120 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u368|_al_u369  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [5],\u2_Display/counta [6]}),
    .d({\u2_Display/n4911 [5],\u2_Display/n4911 [6]}),
    .f({\u2_Display/n6096 ,\u2_Display/n6095 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u3691 (
    .b({open_n35041,\u2_Display/n2242 [0]}),
    .c({open_n35042,\u2_Display/n2240 }),
    .d({open_n35045,\u2_Display/n2239 }),
    .f({open_n35063,\u2_Display/n2274 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3692|_al_u3693  (
    .b({\u2_Display/n2242 [1],\u2_Display/n2242 [2]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2238 ,\u2_Display/n2237 }),
    .f({\u2_Display/n2273 ,\u2_Display/n2272 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3694|_al_u3697  (
    .b({\u2_Display/n2242 [3],\u2_Display/n2242 [6]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2236 ,\u2_Display/n2233 }),
    .f({\u2_Display/n2271 ,\u2_Display/n2268 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3695|_al_u3696  (
    .b({\u2_Display/n2242 [4],\u2_Display/n2242 [5]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2235 ,\u2_Display/n2234 }),
    .f({\u2_Display/n2270 ,\u2_Display/n2269 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3698|_al_u3699  (
    .b({\u2_Display/n2242 [7],\u2_Display/n2242 [8]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2232 ,\u2_Display/n2231 }),
    .f({\u2_Display/n2267 ,\u2_Display/n2266 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3700|_al_u3701  (
    .b({\u2_Display/n2242 [9],\u2_Display/n2242 [10]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2230 ,\u2_Display/n2229 }),
    .f({\u2_Display/n2265 ,\u2_Display/n2264 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3702|_al_u3703  (
    .b({\u2_Display/n2242 [11],\u2_Display/n2242 [12]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2228 ,\u2_Display/n2227 }),
    .f({\u2_Display/n2263 ,\u2_Display/n2262 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3704|_al_u3705  (
    .b({\u2_Display/n2242 [13],\u2_Display/n2242 [14]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2226 ,\u2_Display/n2225 }),
    .f({\u2_Display/n2261 ,\u2_Display/n2260 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3706|_al_u3709  (
    .b({\u2_Display/n2242 [15],\u2_Display/n2242 [18]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2224 ,\u2_Display/n2221 }),
    .f({\u2_Display/n2259 ,\u2_Display/n2256 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u3707 (
    .b({open_n35279,\u2_Display/n2242 [16]}),
    .c({open_n35280,\u2_Display/n2240 }),
    .d({open_n35283,\u2_Display/n2223 }),
    .f({open_n35301,\u2_Display/n2258 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3708|_al_u3712  (
    .b({\u2_Display/n2242 [17],\u2_Display/n2242 [21]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2222 ,\u2_Display/n2218 }),
    .f({\u2_Display/n2257 ,\u2_Display/n2253 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u370|_al_u371  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [7],\u2_Display/counta [8]}),
    .d({\u2_Display/n4911 [7],\u2_Display/n4911 [8]}),
    .f({\u2_Display/n6094 ,\u2_Display/n6093 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3710|_al_u3715  (
    .b({\u2_Display/n2242 [19],\u2_Display/n2242 [24]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2220 ,\u2_Display/n2215 }),
    .f({\u2_Display/n2255 ,\u2_Display/n2250 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3711|_al_u3713  (
    .b({\u2_Display/n2242 [20],\u2_Display/n2242 [22]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2219 ,\u2_Display/n2217 }),
    .f({\u2_Display/n2254 ,\u2_Display/n2252 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3714|_al_u3717  (
    .b({\u2_Display/n2242 [23],\u2_Display/n2242 [26]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2216 ,\u2_Display/n2213 }),
    .f({\u2_Display/n2251 ,\u2_Display/n2248 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3716|_al_u3720  (
    .b({\u2_Display/n2242 [25],\u2_Display/n2242 [29]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2214 ,\u2_Display/n2210 }),
    .f({\u2_Display/n2249 ,\u2_Display/n2245 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3718|_al_u3722  (
    .b({\u2_Display/n2242 [27],\u2_Display/n2240 }),
    .c({\u2_Display/n2240 ,\u2_Display/n2242 [31]}),
    .d({\u2_Display/n2212 ,\u2_Display/n2208 }),
    .f({\u2_Display/n2247 ,\u2_Display/n2243 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3719|_al_u3721  (
    .b({\u2_Display/n2242 [28],\u2_Display/n2242 [30]}),
    .c({\u2_Display/n2240 ,\u2_Display/n2240 }),
    .d({\u2_Display/n2211 ,\u2_Display/n2209 }),
    .f({\u2_Display/n2246 ,\u2_Display/n2244 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3724|_al_u3725  (
    .b({\u2_Display/n3365 [1],\u2_Display/n3365 [2]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3361 ,\u2_Display/n3360 }),
    .f({\u2_Display/n3396 ,\u2_Display/n3395 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3726|_al_u3727  (
    .b({\u2_Display/n3365 [3],\u2_Display/n3365 [4]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3359 ,\u2_Display/n3358 }),
    .f({\u2_Display/n3394 ,\u2_Display/n3393 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3728|_al_u3729  (
    .b({\u2_Display/n3365 [5],\u2_Display/n3365 [6]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3357 ,\u2_Display/n3356 }),
    .f({\u2_Display/n3392 ,\u2_Display/n3391 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3730|_al_u3733  (
    .b({\u2_Display/n3365 [7],\u2_Display/n3365 [10]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3355 ,\u2_Display/n3352 }),
    .f({\u2_Display/n3390 ,\u2_Display/n3387 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3732|_al_u3736  (
    .b({\u2_Display/n3365 [9],\u2_Display/n3365 [13]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3353 ,\u2_Display/n3349 }),
    .f({\u2_Display/n3388 ,\u2_Display/n3384 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3734|_al_u3740  (
    .b({\u2_Display/n3365 [11],\u2_Display/n3365 [17]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3351 ,\u2_Display/n3345 }),
    .f({\u2_Display/n3386 ,\u2_Display/n3380 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3735|_al_u3737  (
    .b({\u2_Display/n3365 [12],\u2_Display/n3365 [14]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3350 ,\u2_Display/n3348 }),
    .f({\u2_Display/n3385 ,\u2_Display/n3383 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3738|_al_u3743  (
    .b({\u2_Display/n3365 [15],\u2_Display/n3365 [20]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3347 ,\u2_Display/n3342 }),
    .f({\u2_Display/n3382 ,\u2_Display/n3377 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3739|_al_u3741  (
    .b({\u2_Display/n3365 [16],\u2_Display/n3365 [18]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3346 ,\u2_Display/n3344 }),
    .f({\u2_Display/n3381 ,\u2_Display/n3379 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u373|_al_u372  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c(\u2_Display/counta [10:9]),
    .d(\u2_Display/n4911 [10:9]),
    .f({\u2_Display/n6091 ,\u2_Display/n6092 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3742|_al_u3745  (
    .b({\u2_Display/n3365 [19],\u2_Display/n3365 [22]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3343 ,\u2_Display/n3340 }),
    .f({\u2_Display/n3378 ,\u2_Display/n3375 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3744|_al_u3748  (
    .b({\u2_Display/n3365 [21],\u2_Display/n3365 [25]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3341 ,\u2_Display/n3337 }),
    .f({\u2_Display/n3376 ,\u2_Display/n3372 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3746|_al_u3884  (
    .b({\u2_Display/n3365 [23],\u2_Display/n3400 [1]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3398 }),
    .d({\u2_Display/n3339 ,\u2_Display/n3396 }),
    .f({\u2_Display/n3374 ,\u2_Display/n3431 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3747|_al_u3749  (
    .b({\u2_Display/n3365 [24],\u2_Display/n3365 [26]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3338 ,\u2_Display/n3336 }),
    .f({\u2_Display/n3373 ,\u2_Display/n3371 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u374|_al_u377  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [11],\u2_Display/counta [14]}),
    .d({\u2_Display/n4911 [11],\u2_Display/n4911 [14]}),
    .f({\u2_Display/n6090 ,\u2_Display/n6087 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u375 (
    .b({open_n35907,\u2_Display/n4909 }),
    .c({open_n35908,\u2_Display/counta [12]}),
    .d({open_n35911,\u2_Display/n4911 [12]}),
    .f({open_n35929,\u2_Display/n6089 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3750|_al_u3751  (
    .b({\u2_Display/n3365 [27],\u2_Display/n3365 [28]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3335 ,\u2_Display/n3334 }),
    .f({\u2_Display/n3370 ,\u2_Display/n3369 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3752|_al_u3753  (
    .b({\u2_Display/n3365 [29],\u2_Display/n3365 [30]}),
    .c({\u2_Display/n3363 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3333 ,\u2_Display/n3332 }),
    .f({\u2_Display/n3368 ,\u2_Display/n3367 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3756|_al_u3757  (
    .b({\u2_Display/n4523 [1],\u2_Display/n4523 [2]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4519 ,\u2_Display/n4518 }),
    .f({\u2_Display/n4554 ,\u2_Display/n4553 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3758|_al_u3761  (
    .b({\u2_Display/n4523 [3],\u2_Display/n4523 [6]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4517 ,\u2_Display/n4514 }),
    .f({\u2_Display/n4552 ,\u2_Display/n4549 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3759|_al_u3760  (
    .b({\u2_Display/n4523 [4],\u2_Display/n4523 [5]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4516 ,\u2_Display/n4515 }),
    .f({\u2_Display/n4551 ,\u2_Display/n4550 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3762|_al_u3764  (
    .b({\u2_Display/n4523 [7],\u2_Display/n4523 [9]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4513 ,\u2_Display/n4511 }),
    .f({\u2_Display/n4548 ,\u2_Display/n4546 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3765|_al_u3763  (
    .b({\u2_Display/n4523 [10],\u2_Display/n4523 [8]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4510 ,\u2_Display/n4512 }),
    .f({\u2_Display/n4545 ,\u2_Display/n4547 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3766|_al_u3769  (
    .b({\u2_Display/n4523 [11],\u2_Display/n4523 [14]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4509 ,\u2_Display/n4506 }),
    .f({\u2_Display/n4544 ,\u2_Display/n4541 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u3767 (
    .b({open_n36141,\u2_Display/n4523 [12]}),
    .c({open_n36142,\u2_Display/n4521 }),
    .d({open_n36145,\u2_Display/n4508 }),
    .f({open_n36163,\u2_Display/n4543 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3768|_al_u3772  (
    .b({\u2_Display/n4523 [13],\u2_Display/n4523 [17]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4507 ,\u2_Display/n4503 }),
    .f({\u2_Display/n4542 ,\u2_Display/n4538 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u376|_al_u379  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [13],\u2_Display/counta [16]}),
    .d({\u2_Display/n4911 [13],\u2_Display/n4911 [16]}),
    .f({\u2_Display/n6088 ,\u2_Display/n6085 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3770|_al_u3775  (
    .b({\u2_Display/n4523 [15],\u2_Display/n4523 [20]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4505 ,\u2_Display/n4500 }),
    .f({\u2_Display/n4540 ,\u2_Display/n4535 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3771|_al_u3773  (
    .b({\u2_Display/n4523 [16],\u2_Display/n4523 [18]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4504 ,\u2_Display/n4502 }),
    .f({\u2_Display/n4539 ,\u2_Display/n4537 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3774|_al_u3777  (
    .b({\u2_Display/n4523 [19],\u2_Display/n4523 [22]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4501 ,\u2_Display/n4498 }),
    .f({\u2_Display/n4536 ,\u2_Display/n4533 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3776|_al_u3779  (
    .b({\u2_Display/n4523 [21],\u2_Display/n4523 [24]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4499 ,\u2_Display/n4496 }),
    .f({\u2_Display/n4534 ,\u2_Display/n4531 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3778|_al_u3781  (
    .b({\u2_Display/n4523 [23],\u2_Display/n4523 [26]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4497 ,\u2_Display/n4494 }),
    .f({\u2_Display/n4532 ,\u2_Display/n4529 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3780|_al_u3783  (
    .b({\u2_Display/n4523 [25],\u2_Display/n4523 [28]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4495 ,\u2_Display/n4492 }),
    .f({\u2_Display/n4530 ,\u2_Display/n4527 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3782|_al_u3785  (
    .b({\u2_Display/n4523 [27],\u2_Display/n4523 [30]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4493 ,\u2_Display/n4490 }),
    .f({\u2_Display/n4528 ,\u2_Display/n4525 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3784|_al_u3786  (
    .b({\u2_Display/n4523 [29],\u2_Display/n4523 [31]}),
    .c({\u2_Display/n4521 ,\u2_Display/n4521 }),
    .d({\u2_Display/n4491 ,\u2_Display/n4489 }),
    .f({\u2_Display/n4526 ,\u2_Display/n4524 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u3787 (
    .b({open_n36411,\u2_Display/n5646 [0]}),
    .c({open_n36412,\u2_Display/n5644 }),
    .d({open_n36415,\u2_Display/n5643 }),
    .f({open_n36433,\u2_Display/n5678 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3788|_al_u3789  (
    .b({\u2_Display/n5646 [1],\u2_Display/n5646 [2]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5642 ,\u2_Display/n5641 }),
    .f({\u2_Display/n5677 ,\u2_Display/n5676 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u378|_al_u381  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [15],\u2_Display/counta [18]}),
    .d({\u2_Display/n4911 [15],\u2_Display/n4911 [18]}),
    .f({\u2_Display/n6086 ,\u2_Display/n6083 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3790|_al_u3791  (
    .b({\u2_Display/n5646 [3],\u2_Display/n5646 [4]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5640 ,\u2_Display/n5639 }),
    .f({\u2_Display/n5675 ,\u2_Display/n5674 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3792|_al_u3793  (
    .b({\u2_Display/n5646 [5],\u2_Display/n5646 [6]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5638 ,\u2_Display/n5637 }),
    .f({\u2_Display/n5673 ,\u2_Display/n5672 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3794|_al_u3796  (
    .b({\u2_Display/n5646 [7],\u2_Display/n5646 [9]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5636 ,\u2_Display/n5634 }),
    .f({\u2_Display/n5671 ,\u2_Display/n5669 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3798|_al_u3795  (
    .b({\u2_Display/n5646 [11],\u2_Display/n5646 [8]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5632 ,\u2_Display/n5635 }),
    .f({\u2_Display/n5667 ,\u2_Display/n5670 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3799|_al_u3797  (
    .b({\u2_Display/n5646 [12],\u2_Display/n5646 [10]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5631 ,\u2_Display/n5633 }),
    .f({\u2_Display/n5666 ,\u2_Display/n5668 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3800|_al_u3803  (
    .b({\u2_Display/n5646 [13],\u2_Display/n5646 [16]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5630 ,\u2_Display/n5627 }),
    .f({\u2_Display/n5665 ,\u2_Display/n5662 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u3801 (
    .b({open_n36649,\u2_Display/n5646 [14]}),
    .c({open_n36650,\u2_Display/n5644 }),
    .d({open_n36653,\u2_Display/n5629 }),
    .f({open_n36671,\u2_Display/n5664 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3802|_al_u3805  (
    .b({\u2_Display/n5646 [15],\u2_Display/n5646 [18]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5628 ,\u2_Display/n5625 }),
    .f({\u2_Display/n5663 ,\u2_Display/n5660 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3804|_al_u3807  (
    .b({\u2_Display/n5646 [17],\u2_Display/n5646 [20]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5626 ,\u2_Display/n5623 }),
    .f({\u2_Display/n5661 ,\u2_Display/n5658 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3806|_al_u3809  (
    .b({\u2_Display/n5646 [19],\u2_Display/n5646 [22]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5624 ,\u2_Display/n5621 }),
    .f({\u2_Display/n5659 ,\u2_Display/n5656 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3808|_al_u3812  (
    .b({\u2_Display/n5646 [21],\u2_Display/n5646 [25]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5622 ,\u2_Display/n5618 }),
    .f({\u2_Display/n5657 ,\u2_Display/n5653 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u380|_al_u383  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [17],\u2_Display/counta [20]}),
    .d({\u2_Display/n4911 [17],\u2_Display/n4911 [20]}),
    .f({\u2_Display/n6084 ,\u2_Display/n6081 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3810|_al_u3815  (
    .b({\u2_Display/n5646 [23],\u2_Display/n5646 [28]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5620 ,\u2_Display/n5615 }),
    .f({\u2_Display/n5655 ,\u2_Display/n5650 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3811|_al_u3813  (
    .b({\u2_Display/n5646 [24],\u2_Display/n5646 [26]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5619 ,\u2_Display/n5617 }),
    .f({\u2_Display/n5654 ,\u2_Display/n5652 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3814|_al_u3817  (
    .b({\u2_Display/n5646 [27],\u2_Display/n5646 [30]}),
    .c({\u2_Display/n5644 ,\u2_Display/n5644 }),
    .d({\u2_Display/n5616 ,\u2_Display/n5613 }),
    .f({\u2_Display/n5651 ,\u2_Display/n5648 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3816|_al_u3818  (
    .b({\u2_Display/n5646 [29],\u2_Display/n5644 }),
    .c({\u2_Display/n5644 ,\u2_Display/n5646 [31]}),
    .d({\u2_Display/n5614 ,\u2_Display/n5612 }),
    .f({\u2_Display/n5649 ,\u2_Display/n5647 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3820|_al_u3821  (
    .b({\u2_Display/n1154 [1],\u2_Display/n1154 [2]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1150 ,\u2_Display/n1149 }),
    .f({\u2_Display/n1185 ,\u2_Display/n1184 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3822|_al_u3823  (
    .b({\u2_Display/n1154 [3],\u2_Display/n1154 [4]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1148 ,\u2_Display/n1147 }),
    .f({\u2_Display/n1183 ,\u2_Display/n1182 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3824|_al_u3825  (
    .b({\u2_Display/n1154 [5],\u2_Display/n1154 [6]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1146 ,\u2_Display/n1145 }),
    .f({\u2_Display/n1181 ,\u2_Display/n1180 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3826|_al_u3828  (
    .b({\u2_Display/n1154 [7],\u2_Display/n1154 [9]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1144 ,\u2_Display/n1142 }),
    .f({\u2_Display/n1179 ,\u2_Display/n1177 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3829|_al_u3819  (
    .b({\u2_Display/n1154 [10],\u2_Display/n1154 [0]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1141 ,\u2_Display/n1151 }),
    .f({\u2_Display/n1176 ,\u2_Display/n1186 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u382|_al_u385  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [19],\u2_Display/counta [22]}),
    .d({\u2_Display/n4911 [19],\u2_Display/n4911 [22]}),
    .f({\u2_Display/n6082 ,\u2_Display/n6079 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u3830|_al_u3831  (
    .b({\u2_Display/n1140 ,\u2_Display/n1154 [12]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1154 [11],\u2_Display/n1139 }),
    .f({\u2_Display/n1175 ,\u2_Display/n1174 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3832|_al_u3827  (
    .b({\u2_Display/n1154 [13],\u2_Display/n1154 [8]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1138 ,\u2_Display/n1143 }),
    .f({\u2_Display/n1173 ,\u2_Display/n1178 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3833|_al_u3835  (
    .b({\u2_Display/n1154 [14],\u2_Display/n1154 [16]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1137 ,\u2_Display/n1135 }),
    .f({\u2_Display/n1172 ,\u2_Display/n1170 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3834|_al_u3837  (
    .b({\u2_Display/n1154 [15],\u2_Display/n1154 [18]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1136 ,\u2_Display/n1133 }),
    .f({\u2_Display/n1171 ,\u2_Display/n1168 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3836|_al_u3839  (
    .b({\u2_Display/n1154 [17],\u2_Display/n1154 [20]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1134 ,\u2_Display/n1131 }),
    .f({\u2_Display/n1169 ,\u2_Display/n1166 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u3838|_al_u3841  (
    .b({\u2_Display/n1152 ,\u2_Display/n1154 [22]}),
    .c({\u2_Display/n1154 [19],\u2_Display/n1152 }),
    .d({\u2_Display/n1132 ,\u2_Display/n1129 }),
    .f({\u2_Display/n1167 ,\u2_Display/n1164 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3840|_al_u3843  (
    .b({\u2_Display/n1154 [21],\u2_Display/n1154 [24]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1130 ,\u2_Display/n1127 }),
    .f({\u2_Display/n1165 ,\u2_Display/n1162 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3842|_al_u3845  (
    .b({\u2_Display/n1154 [23],\u2_Display/n1154 [26]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1128 ,\u2_Display/n1125 }),
    .f({\u2_Display/n1163 ,\u2_Display/n1160 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3844|_al_u3847  (
    .b({\u2_Display/n1154 [25],\u2_Display/n1154 [28]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1126 ,\u2_Display/n1123 }),
    .f({\u2_Display/n1161 ,\u2_Display/n1158 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3846|_al_u3849  (
    .b({\u2_Display/n1154 [27],\u2_Display/n1154 [30]}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1124 ,\u2_Display/n1121 }),
    .f({\u2_Display/n1159 ,\u2_Display/n1156 }));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111101000001010),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3848|_al_u3850  (
    .a({open_n37291,\u2_Display/n1154 [31]}),
    .b({\u2_Display/n1154 [29],open_n37292}),
    .c({\u2_Display/n1152 ,\u2_Display/n1152 }),
    .d({\u2_Display/n1122 ,\u2_Display/n1120 }),
    .f({\u2_Display/n1157 ,\u2_Display/n1155 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u384|_al_u388  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [21],\u2_Display/counta [25]}),
    .d({\u2_Display/n4911 [21],\u2_Display/n4911 [25]}),
    .f({\u2_Display/n6080 ,\u2_Display/n6076 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3851|_al_u3853  (
    .b({\u2_Display/n2277 [0],\u2_Display/n2277 [2]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2274 ,\u2_Display/n2272 }),
    .f({\u2_Display/n2309 ,\u2_Display/n2307 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u3852 (
    .b({open_n37367,\u2_Display/n2277 [1]}),
    .c({open_n37368,\u2_Display/n2275 }),
    .d({open_n37371,\u2_Display/n2273 }),
    .f({open_n37389,\u2_Display/n2308 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3854|_al_u3855  (
    .b({\u2_Display/n2277 [3],\u2_Display/n2277 [4]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2271 ,\u2_Display/n2270 }),
    .f({\u2_Display/n2306 ,\u2_Display/n2305 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3856|_al_u3857  (
    .b({\u2_Display/n2277 [5],\u2_Display/n2277 [6]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2269 ,\u2_Display/n2268 }),
    .f({\u2_Display/n2304 ,\u2_Display/n2303 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3858|_al_u3860  (
    .b({\u2_Display/n2277 [7],\u2_Display/n2277 [9]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2267 ,\u2_Display/n2265 }),
    .f({\u2_Display/n2302 ,\u2_Display/n2300 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3861|_al_u3859  (
    .b({\u2_Display/n2277 [10],\u2_Display/n2277 [8]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2264 ,\u2_Display/n2266 }),
    .f({\u2_Display/n2299 ,\u2_Display/n2301 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3862|_al_u3863  (
    .b({\u2_Display/n2277 [11],\u2_Display/n2277 [12]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2263 ,\u2_Display/n2262 }),
    .f({\u2_Display/n2298 ,\u2_Display/n2297 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3864|_al_u3865  (
    .b({\u2_Display/n2277 [13],\u2_Display/n2277 [14]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2261 ,\u2_Display/n2260 }),
    .f({\u2_Display/n2296 ,\u2_Display/n2295 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3866|_al_u3869  (
    .b({\u2_Display/n2277 [15],\u2_Display/n2277 [18]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2259 ,\u2_Display/n2256 }),
    .f({\u2_Display/n2294 ,\u2_Display/n2291 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .MODE("LOGIC"))
    _al_u3867 (
    .b({open_n37575,\u2_Display/n2277 [16]}),
    .c({open_n37576,\u2_Display/n2275 }),
    .d({open_n37579,\u2_Display/n2258 }),
    .f({open_n37593,\u2_Display/n2293 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3868|_al_u3871  (
    .b({\u2_Display/n2277 [17],\u2_Display/n2277 [20]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2257 ,\u2_Display/n2254 }),
    .f({\u2_Display/n2292 ,\u2_Display/n2289 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u386|_al_u391  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [23],\u2_Display/counta [28]}),
    .d({\u2_Display/n4911 [23],\u2_Display/n4911 [28]}),
    .f({\u2_Display/n6078 ,\u2_Display/n6073 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3870|_al_u3873  (
    .b({\u2_Display/n2277 [19],\u2_Display/n2277 [22]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2255 ,\u2_Display/n2252 }),
    .f({\u2_Display/n2290 ,\u2_Display/n2287 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3872|_al_u3875  (
    .b({\u2_Display/n2277 [21],\u2_Display/n2277 [24]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2253 ,\u2_Display/n2250 }),
    .f({\u2_Display/n2288 ,\u2_Display/n2285 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3874|_al_u3877  (
    .b({\u2_Display/n2277 [23],\u2_Display/n2277 [26]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2251 ,\u2_Display/n2248 }),
    .f({\u2_Display/n2286 ,\u2_Display/n2283 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3876|_al_u3879  (
    .b({\u2_Display/n2277 [25],\u2_Display/n2277 [28]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2249 ,\u2_Display/n2246 }),
    .f({\u2_Display/n2284 ,\u2_Display/n2281 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3878|_al_u3881  (
    .b({\u2_Display/n2277 [27],\u2_Display/n2277 [30]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2247 ,\u2_Display/n2244 }),
    .f({\u2_Display/n2282 ,\u2_Display/n2279 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u387|_al_u389  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [24],\u2_Display/counta [26]}),
    .d({\u2_Display/n4911 [24],\u2_Display/n4911 [26]}),
    .f({\u2_Display/n6077 ,\u2_Display/n6075 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3880|_al_u3882  (
    .b({\u2_Display/n2277 [29],\u2_Display/n2277 [31]}),
    .c({\u2_Display/n2275 ,\u2_Display/n2275 }),
    .d({\u2_Display/n2245 ,\u2_Display/n2243 }),
    .f({\u2_Display/n2280 ,\u2_Display/n2278 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3883|_al_u3885  (
    .b({\u2_Display/n3400 [0],\u2_Display/n3400 [2]}),
    .c({\u2_Display/n3398 ,\u2_Display/n3398 }),
    .d({\u2_Display/n3397 ,\u2_Display/n3395 }),
    .f({\u2_Display/n3432 ,\u2_Display/n3430 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3886|_al_u3889  (
    .b({\u2_Display/n3400 [3],\u2_Display/n3400 [6]}),
    .c({\u2_Display/n3398 ,\u2_Display/n3398 }),
    .d({\u2_Display/n3394 ,\u2_Display/n3391 }),
    .f({\u2_Display/n3429 ,\u2_Display/n3426 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3887|_al_u3888  (
    .b({\u2_Display/n3400 [4],\u2_Display/n3400 [5]}),
    .c({\u2_Display/n3398 ,\u2_Display/n3398 }),
    .d({\u2_Display/n3393 ,\u2_Display/n3392 }),
    .f({\u2_Display/n3428 ,\u2_Display/n3427 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3890|_al_u3892  (
    .b({\u2_Display/n3400 [7],\u2_Display/n3400 [9]}),
    .c({\u2_Display/n3398 ,\u2_Display/n3398 }),
    .d({\u2_Display/n3390 ,\u2_Display/n3388 }),
    .f({\u2_Display/n3425 ,\u2_Display/n3423 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3893|_al_u3891  (
    .b({\u2_Display/n3400 [10],\u2_Display/n3400 [8]}),
    .c({\u2_Display/n3398 ,\u2_Display/n3398 }),
    .d({\u2_Display/n3387 ,\u2_Display/n3389 }),
    .f({\u2_Display/n3422 ,\u2_Display/n3424 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3894|_al_u3754  (
    .b({\u2_Display/n3400 [11],\u2_Display/n3365 [31]}),
    .c({\u2_Display/n3398 ,\u2_Display/n3363 }),
    .d({\u2_Display/n3386 ,\u2_Display/n3331 }),
    .f({\u2_Display/n3421 ,\u2_Display/n3366 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3895|_al_u3897  (
    .b({\u2_Display/n3400 [12],\u2_Display/n3400 [14]}),
    .c({\u2_Display/n3398 ,\u2_Display/n3398 }),
    .d({\u2_Display/n3385 ,\u2_Display/n3383 }),
    .f({\u2_Display/n3420 ,\u2_Display/n3418 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3896|_al_u3899  (
    .b({\u2_Display/n3400 [13],\u2_Display/n3400 [16]}),
    .c({\u2_Display/n3398 ,\u2_Display/n3398 }),
    .d({\u2_Display/n3384 ,\u2_Display/n3381 }),
    .f({\u2_Display/n3419 ,\u2_Display/n3416 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3898|_al_u3901  (
    .b({\u2_Display/n3400 [15],\u2_Display/n3400 [18]}),
    .c({\u2_Display/n3398 ,\u2_Display/n3398 }),
    .d({\u2_Display/n3382 ,\u2_Display/n3379 }),
    .f({\u2_Display/n3417 ,\u2_Display/n3414 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3900|_al_u3903  (
    .b({\u2_Display/n3400 [17],\u2_Display/n3400 [20]}),
    .c({\u2_Display/n3398 ,\u2_Display/n3398 }),
    .d({\u2_Display/n3380 ,\u2_Display/n3377 }),
    .f({\u2_Display/n3415 ,\u2_Display/n3412 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3902|_al_u3905  (
    .b({\u2_Display/n3400 [19],\u2_Display/n3400 [22]}),
    .c({\u2_Display/n3398 ,\u2_Display/n3398 }),
    .d({\u2_Display/n3378 ,\u2_Display/n3375 }),
    .f({\u2_Display/n3413 ,\u2_Display/n3410 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3904|_al_u3907  (
    .b({\u2_Display/n3400 [21],\u2_Display/n3400 [24]}),
    .c({\u2_Display/n3398 ,\u2_Display/n3398 }),
    .d({\u2_Display/n3376 ,\u2_Display/n3373 }),
    .f({\u2_Display/n3411 ,\u2_Display/n3408 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3906|_al_u3909  (
    .b({\u2_Display/n3400 [23],\u2_Display/n3400 [26]}),
    .c({\u2_Display/n3398 ,\u2_Display/n3398 }),
    .d({\u2_Display/n3374 ,\u2_Display/n3371 }),
    .f({\u2_Display/n3409 ,\u2_Display/n3406 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u3908|_al_u3911  (
    .b({\u2_Display/n3398 ,\u2_Display/n3400 [28]}),
    .c({\u2_Display/n3400 [25],\u2_Display/n3398 }),
    .d({\u2_Display/n3372 ,\u2_Display/n3369 }),
    .f({\u2_Display/n3407 ,\u2_Display/n3404 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u390|_al_u393  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [27],\u2_Display/counta [30]}),
    .d({\u2_Display/n4911 [27],\u2_Display/n4911 [30]}),
    .f({\u2_Display/n6074 ,\u2_Display/n6071 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"))
    \_al_u3910|_al_u3913  (
    .b({\u2_Display/n3398 ,\u2_Display/n3400 [30]}),
    .c({\u2_Display/n3400 [27],\u2_Display/n3398 }),
    .d({\u2_Display/n3370 ,\u2_Display/n3367 }),
    .f({\u2_Display/n3405 ,\u2_Display/n3402 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3912|_al_u3914  (
    .b({\u2_Display/n3400 [29],\u2_Display/n3398 }),
    .c({\u2_Display/n3398 ,\u2_Display/n3400 [31]}),
    .d({\u2_Display/n3368 ,\u2_Display/n3366 }),
    .f({\u2_Display/n3403 ,\u2_Display/n3401 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3916|_al_u3925  (
    .b({\u2_Display/n3435 [0],\u2_Display/n3435 [2]}),
    .c({\u2_Display/n3433 ,\u2_Display/n3433 }),
    .d({\u2_Display/n3432 ,\u2_Display/n3430 }),
    .f({_al_u3916_o,_al_u3925_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3917|_al_u3937  (
    .b({\u2_Display/n1189 [0],\u2_Display/n1189 [5]}),
    .c({\u2_Display/n1187 ,\u2_Display/n1187 }),
    .d({\u2_Display/n1186 ,\u2_Display/n1181 }),
    .f({_al_u3917_o,_al_u3937_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~((0*~(A)*~(D)+0*A*~(D)+~(0)*A*D+0*A*D))*~(C)+B*(0*~(A)*~(D)+0*A*~(D)+~(0)*A*D+0*A*D)*~(C)+~(B)*(0*~(A)*~(D)+0*A*~(D)+~(0)*A*D+0*A*D)*C+B*(0*~(A)*~(D)+0*A*~(D)+~(0)*A*D+0*A*D)*C)"),
    //.LUTF1("~(A*~((0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D))*~(C)+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*~(C)+~(A)*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C)"),
    //.LUTG0("(B*~((1*~(A)*~(D)+1*A*~(D)+~(1)*A*D+1*A*D))*~(C)+B*(1*~(A)*~(D)+1*A*~(D)+~(1)*A*D+1*A*D)*~(C)+~(B)*(1*~(A)*~(D)+1*A*~(D)+~(1)*A*D+1*A*D)*C+B*(1*~(A)*~(D)+1*A*~(D)+~(1)*A*D+1*A*D)*C)"),
    //.LUTG1("~(A*~((1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D))*~(C)+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*~(C)+~(A)*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C)"),
    .INIT_LUTF0(16'b1010110000001100),
    .INIT_LUTF1(16'b0011010111110101),
    .INIT_LUTG0(16'b1010110011111100),
    .INIT_LUTG1(16'b0011010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3918|_al_u3926  (
    .a({_al_u3916_o,_al_u3924_o}),
    .b({_al_u3917_o,_al_u3925_o}),
    .c({\u2_Display/mux11_b0_sel_is_0_o ,\u2_Display/mux11_b0_sel_is_0_o }),
    .d({on_off_pad[4],on_off_pad[4]}),
    .e({\u2_Display/j [0],\u2_Display/j [2]}),
    .f({_al_u3918_o,_al_u3926_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u3920 (
    .b({open_n38315,\u2_Display/n3435 [1]}),
    .c({open_n38316,\u2_Display/n3433 }),
    .d({open_n38319,\u2_Display/n3431 }),
    .f({open_n38337,_al_u3920_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3921|_al_u3924  (
    .b({\u2_Display/n1189 [1],\u2_Display/n1189 [2]}),
    .c({\u2_Display/n1187 ,\u2_Display/n1187 }),
    .d({\u2_Display/n1185 ,\u2_Display/n1184 }),
    .f({_al_u3921_o,_al_u3924_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3928|_al_u3936  (
    .b({\u2_Display/n3435 [3],\u2_Display/n3435 [5]}),
    .c({\u2_Display/n3433 ,\u2_Display/n3433 }),
    .d({\u2_Display/n3429 ,\u2_Display/n3427 }),
    .f({_al_u3928_o,_al_u3936_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3929|_al_u3948  (
    .b({\u2_Display/n1189 [3],\u2_Display/n1189 [8]}),
    .c({\u2_Display/n1187 ,\u2_Display/n1187 }),
    .d({\u2_Display/n1183 ,\u2_Display/n1178 }),
    .f({_al_u3929_o,_al_u3948_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u392|_al_u394  (
    .b({\u2_Display/n4909 ,\u2_Display/n4909 }),
    .c({\u2_Display/counta [29],\u2_Display/counta [31]}),
    .d({\u2_Display/n4911 [29],\u2_Display/n4911 [31]}),
    .f({\u2_Display/n6072 ,\u2_Display/n6070 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~((0*~(A)*~(D)+0*A*~(D)+~(0)*A*D+0*A*D))*~(C)+B*(0*~(A)*~(D)+0*A*~(D)+~(0)*A*D+0*A*D)*~(C)+~(B)*(0*~(A)*~(D)+0*A*~(D)+~(0)*A*D+0*A*D)*C+B*(0*~(A)*~(D)+0*A*~(D)+~(0)*A*D+0*A*D)*C)"),
    //.LUTF1("~(A*~((0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D))*~(C)+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*~(C)+~(A)*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C)"),
    //.LUTG0("(B*~((1*~(A)*~(D)+1*A*~(D)+~(1)*A*D+1*A*D))*~(C)+B*(1*~(A)*~(D)+1*A*~(D)+~(1)*A*D+1*A*D)*~(C)+~(B)*(1*~(A)*~(D)+1*A*~(D)+~(1)*A*D+1*A*D)*C+B*(1*~(A)*~(D)+1*A*~(D)+~(1)*A*D+1*A*D)*C)"),
    //.LUTG1("~(A*~((1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D))*~(C)+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*~(C)+~(A)*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C)"),
    .INIT_LUTF0(16'b1010110000001100),
    .INIT_LUTF1(16'b0011010111110101),
    .INIT_LUTG0(16'b1010110011111100),
    .INIT_LUTG1(16'b0011010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3930|_al_u3942  (
    .a({_al_u3928_o,_al_u3940_o}),
    .b({_al_u3929_o,_al_u3941_o}),
    .c({\u2_Display/mux11_b0_sel_is_0_o ,\u2_Display/mux11_b0_sel_is_0_o }),
    .d({on_off_pad[4],on_off_pad[4]}),
    .e({\u2_Display/j [3],\u2_Display/j [6]}),
    .f({_al_u3930_o,_al_u3942_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3932|_al_u3941  (
    .b({\u2_Display/n3435 [4],\u2_Display/n3435 [6]}),
    .c({\u2_Display/n3433 ,\u2_Display/n3433 }),
    .d({\u2_Display/n3428 ,\u2_Display/n3426 }),
    .f({_al_u3932_o,_al_u3941_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3933|_al_u3940  (
    .b({\u2_Display/n1189 [4],\u2_Display/n1189 [6]}),
    .c({\u2_Display/n1187 ,\u2_Display/n1187 }),
    .d({\u2_Display/n1182 ,\u2_Display/n1180 }),
    .f({_al_u3933_o,_al_u3940_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(A*~((0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D))*~(C)+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*~(C)+~(A)*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C)"),
    //.LUTF1("~(A*~((0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D))*~(C)+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*~(C)+~(A)*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C)"),
    //.LUTG0("~(A*~((1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D))*~(C)+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*~(C)+~(A)*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C)"),
    //.LUTG1("~(A*~((1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D))*~(C)+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*~(C)+~(A)*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C)"),
    .INIT_LUTF0(16'b0011010111110101),
    .INIT_LUTF1(16'b0011010111110101),
    .INIT_LUTG0(16'b0011010100000101),
    .INIT_LUTG1(16'b0011010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3934|_al_u3938  (
    .a({_al_u3932_o,_al_u3936_o}),
    .b({_al_u3933_o,_al_u3937_o}),
    .c({\u2_Display/mux11_b0_sel_is_0_o ,\u2_Display/mux11_b0_sel_is_0_o }),
    .d({on_off_pad[4],on_off_pad[4]}),
    .e({\u2_Display/j [4],\u2_Display/j [5]}),
    .f({_al_u3934_o,_al_u3938_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3944|_al_u3949  (
    .b({\u2_Display/n3435 [7],\u2_Display/n3435 [8]}),
    .c({\u2_Display/n3433 ,\u2_Display/n3433 }),
    .d({\u2_Display/n3425 ,\u2_Display/n3424 }),
    .f({_al_u3944_o,_al_u3949_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3945|_al_u3953  (
    .b({\u2_Display/n1189 [7],\u2_Display/n1189 [9]}),
    .c({\u2_Display/n1187 ,\u2_Display/n1187 }),
    .d({\u2_Display/n1179 ,\u2_Display/n1177 }),
    .f({_al_u3945_o,_al_u3953_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~((0*~(A)*~(D)+0*A*~(D)+~(0)*A*D+0*A*D))*~(C)+B*(0*~(A)*~(D)+0*A*~(D)+~(0)*A*D+0*A*D)*~(C)+~(B)*(0*~(A)*~(D)+0*A*~(D)+~(0)*A*D+0*A*D)*C+B*(0*~(A)*~(D)+0*A*~(D)+~(0)*A*D+0*A*D)*C)"),
    //.LUTF1("~(A*~((0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D))*~(C)+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*~(C)+~(A)*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C)"),
    //.LUTG0("(B*~((1*~(A)*~(D)+1*A*~(D)+~(1)*A*D+1*A*D))*~(C)+B*(1*~(A)*~(D)+1*A*~(D)+~(1)*A*D+1*A*D)*~(C)+~(B)*(1*~(A)*~(D)+1*A*~(D)+~(1)*A*D+1*A*D)*C+B*(1*~(A)*~(D)+1*A*~(D)+~(1)*A*D+1*A*D)*C)"),
    //.LUTG1("~(A*~((1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D))*~(C)+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*~(C)+~(A)*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C)"),
    .INIT_LUTF0(16'b1010110000001100),
    .INIT_LUTF1(16'b0011010111110101),
    .INIT_LUTG0(16'b1010110011111100),
    .INIT_LUTG1(16'b0011010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3946|_al_u3950  (
    .a({_al_u3944_o,_al_u3948_o}),
    .b({_al_u3945_o,_al_u3949_o}),
    .c({\u2_Display/mux11_b0_sel_is_0_o ,\u2_Display/mux11_b0_sel_is_0_o }),
    .d({on_off_pad[4],on_off_pad[4]}),
    .e({\u2_Display/j [7],\u2_Display/j [8]}),
    .f({_al_u3946_o,_al_u3950_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(A*~((0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D))*~(C)+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*~(C)+~(A)*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("~(A*~((1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D))*~(C)+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*~(C)+~(A)*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0011010111110101),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b0011010100000101),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3952|_al_u3922  (
    .a({open_n38601,_al_u3920_o}),
    .b({\u2_Display/n3435 [9],_al_u3921_o}),
    .c({\u2_Display/n3433 ,\u2_Display/mux11_b0_sel_is_0_o }),
    .d({\u2_Display/n3423 ,on_off_pad[4]}),
    .e({open_n38604,\u2_Display/j [1]}),
    .f({_al_u3952_o,_al_u3922_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+~(A)*B*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+~(A)*B*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .INIT_LUTF0(16'b0101001101011111),
    .INIT_LUTF1(16'b1010101010111000),
    .INIT_LUTG0(16'b0101011101010111),
    .INIT_LUTG1(16'b1010101010111000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3956|_al_u3963  (
    .a({\u2_Display/n5678 ,\u2_Display/n5677 }),
    .b({on_off_pad[0],on_off_pad[1]}),
    .c({\u2_Display/n5681 [0],on_off_pad[0]}),
    .d({\u2_Display/n5679 ,\u2_Display/n5681 [1]}),
    .e({open_n38627,\u2_Display/n5679 }),
    .f({_al_u3956_o,_al_u3963_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(0)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*0*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*B)"),
    //.LUTF1("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(0)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*0*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*B)"),
    //.LUTG0("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(1)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*1*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*B)"),
    //.LUTG1("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(1)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*1*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*B)"),
    .INIT_LUTF0(16'b1101110111001111),
    .INIT_LUTF1(16'b1101110111001111),
    .INIT_LUTG0(16'b0001000100000011),
    .INIT_LUTG1(16'b0001000100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3957|_al_u3966  (
    .a({\u2_Display/n2309 ,\u2_Display/n2307 }),
    .b({\u2_Display/mux5_b0_sel_is_0_o ,\u2_Display/mux5_b0_sel_is_0_o }),
    .c({\u2_Display/n2312 [0],\u2_Display/n2312 [2]}),
    .d({\u2_Display/n2310 ,\u2_Display/n2310 }),
    .e({\u2_Display/i [0],\u2_Display/i [2]}),
    .f({_al_u3957_o,_al_u3966_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~((D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0))*~(C)+~A*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*~(C)+~(~A)*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*C+~A*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*C)"),
    //.LUTF1("~(~A*~((D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0))*~(C)+~A*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*~(C)+~(~A)*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*C+~A*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*C)"),
    //.LUTG0("~(~A*~((D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1))*~(C)+~A*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*~(C)+~(~A)*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*C+~A*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*C)"),
    //.LUTG1("~(~A*~((D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1))*~(C)+~A*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*~(C)+~(~A)*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*C+~A*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*C)"),
    .INIT_LUTF0(16'b0000101011111010),
    .INIT_LUTF1(16'b0000101011111010),
    .INIT_LUTG0(16'b0011101000111010),
    .INIT_LUTG1(16'b0011101000111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3958|_al_u3967  (
    .a({_al_u3957_o,_al_u3966_o}),
    .b({\u2_Display/n4555 ,\u2_Display/n4553 }),
    .c({on_off_pad[2],on_off_pad[2]}),
    .d({\u2_Display/n4558 [0],\u2_Display/n4558 [2]}),
    .e({\u2_Display/n4556 ,\u2_Display/n4556 }),
    .f({_al_u3958_o,_al_u3967_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u395|_al_u397  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [0],\u2_Display/counta [2]}),
    .d({\u2_Display/n419 [0],\u2_Display/n419 [2]}),
    .f({\u2_Display/n451 ,\u2_Display/n449 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u3960|_al_u3969  (
    .b({\u2_Display/n2312 [1],\u2_Display/n2312 [3]}),
    .c({\u2_Display/n2310 ,\u2_Display/n2310 }),
    .d({\u2_Display/n2308 ,\u2_Display/n2306 }),
    .f({_al_u3960_o,_al_u3969_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1000100011000000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1000100011000000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3961|_al_u3981  (
    .a({open_n38740,\u2_Display/n4550 }),
    .b({\u2_Display/n4558 [1],on_off_pad[2]}),
    .c({\u2_Display/n4556 ,\u2_Display/n4558 [5]}),
    .d({\u2_Display/n4554 ,\u2_Display/n4556 }),
    .f({_al_u3961_o,_al_u3981_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*~(B)*~(D)+(A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*B*~(D)+~((A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C))*B*D+(A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*B*D)"),
    //.LUTF1("~((A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*~(B)*~(D)+(A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*B*~(D)+~((A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C))*B*D+(A*~(0)*~(C)+A*0*~(C)+~(A)*0*C+A*0*C)*B*D)"),
    //.LUTG0("~((A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*~(B)*~(D)+(A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*B*~(D)+~((A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C))*B*D+(A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*B*D)"),
    //.LUTG1("~((A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*~(B)*~(D)+(A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*B*~(D)+~((A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C))*B*D+(A*~(1)*~(C)+A*1*~(C)+~(A)*1*C+A*1*C)*B*D)"),
    .INIT_LUTF0(16'b0011001111110101),
    .INIT_LUTF1(16'b0011001111110101),
    .INIT_LUTG0(16'b0011001100000101),
    .INIT_LUTG1(16'b0011001100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3962|_al_u3971  (
    .a({_al_u3960_o,_al_u3969_o}),
    .b({_al_u3961_o,_al_u3970_o}),
    .c({\u2_Display/mux5_b0_sel_is_0_o ,\u2_Display/mux5_b0_sel_is_0_o }),
    .d({on_off_pad[2],on_off_pad[2]}),
    .e({\u2_Display/i [1],\u2_Display/i [3]}),
    .f({_al_u3962_o,_al_u3971_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .INIT_LUT0(16'b1010101010111000),
    .MODE("LOGIC"))
    _al_u3965 (
    .a({open_n38787,\u2_Display/n5676 }),
    .b({open_n38788,on_off_pad[0]}),
    .c({open_n38789,\u2_Display/n5681 [2]}),
    .d({open_n38792,\u2_Display/n5679 }),
    .f({open_n38806,_al_u3965_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u3970 (
    .b({open_n38814,\u2_Display/n4558 [3]}),
    .c({open_n38815,\u2_Display/n4556 }),
    .d({open_n38818,\u2_Display/n4552 }),
    .f({open_n38836,_al_u3970_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+A*~(B)*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+A*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+A*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+A*B*~(C)*D*0+A*~(B)*C*D*0+A*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+~(A)*B*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+A*~(B)*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+A*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+A*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+A*B*~(C)*D*1+A*~(B)*C*D*1+A*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+~(A)*B*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+~(A)*B*C*D*1)"),
    .INIT_LUTF0(16'b1010111110100011),
    .INIT_LUTF1(16'b0101001101011111),
    .INIT_LUTG0(16'b1010101110101011),
    .INIT_LUTG1(16'b0101011101010111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3972|_al_u3978  (
    .a({\u2_Display/n5675 ,\u2_Display/n5673 }),
    .b({on_off_pad[1],on_off_pad[1]}),
    .c({on_off_pad[0],on_off_pad[0]}),
    .d({\u2_Display/n5681 [3],\u2_Display/n5681 [5]}),
    .e({\u2_Display/n5679 ,\u2_Display/n5679 }),
    .f({_al_u3972_o,_al_u3978_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3974|_al_u3983  (
    .b({\u2_Display/n4558 [4],\u2_Display/n4558 [6]}),
    .c({\u2_Display/n4556 ,\u2_Display/n4556 }),
    .d({\u2_Display/n4551 ,\u2_Display/n4549 }),
    .f({_al_u3974_o,_al_u3983_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(0)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*0*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*B)"),
    //.LUTF1("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(0)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*0*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*B)"),
    //.LUTG0("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(1)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*1*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*B)"),
    //.LUTG1("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(1)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*1*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*B)"),
    .INIT_LUTF0(16'b1101110111001111),
    .INIT_LUTF1(16'b1101110111001111),
    .INIT_LUTG0(16'b0001000100000011),
    .INIT_LUTG1(16'b0001000100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3975|_al_u3984  (
    .a({\u2_Display/n2305 ,\u2_Display/n2303 }),
    .b({\u2_Display/mux5_b0_sel_is_0_o ,\u2_Display/mux5_b0_sel_is_0_o }),
    .c({\u2_Display/n2312 [4],\u2_Display/n2312 [6]}),
    .d({\u2_Display/n2310 ,\u2_Display/n2310 }),
    .e({\u2_Display/i [4],\u2_Display/i [6]}),
    .f({_al_u3975_o,_al_u3984_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+~(A)*B*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+~(A)*B*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+~(A)*B*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+~(A)*B*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+~(A)*B*C*D*1)"),
    .INIT_LUTF0(16'b0101001101011111),
    .INIT_LUTF1(16'b0101001101011111),
    .INIT_LUTG0(16'b0101011101010111),
    .INIT_LUTG1(16'b0101011101010111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3976|_al_u3985  (
    .a({\u2_Display/n5674 ,\u2_Display/n5672 }),
    .b({on_off_pad[1],on_off_pad[1]}),
    .c({on_off_pad[0],on_off_pad[0]}),
    .d({\u2_Display/n5681 [4],\u2_Display/n5681 [6]}),
    .e({\u2_Display/n5679 ,\u2_Display/n5679 }),
    .f({_al_u3976_o,_al_u3985_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3979|_al_u3755  (
    .b({\u2_Display/n2312 [5],\u2_Display/n4523 [0]}),
    .c({\u2_Display/n2310 ,\u2_Display/n4521 }),
    .d({\u2_Display/n2304 ,\u2_Display/n4520 }),
    .f({_al_u3979_o,\u2_Display/n4555 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    //.LUTG0("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT_LUTF0(16'b0000111000000010),
    .INIT_LUTG0(16'b0000111000000010),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u3980 (
    .a({open_n38960,_al_u3979_o}),
    .b({open_n38961,\u2_Display/mux5_b0_sel_is_0_o }),
    .c({open_n38962,on_off_pad[2]}),
    .d({open_n38965,\u2_Display/i [5]}),
    .f({open_n38983,_al_u3980_o}));
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTF1("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    //.LUTG0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG1("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110011111100),
    .INIT_LUTF1(16'b1010101010111000),
    .INIT_LUTG0(16'b0000110011111100),
    .INIT_LUTG1(16'b1010101010111000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3987|u2_Display/reg3_b2  (
    .a({\u2_Display/n5671 ,open_n38989}),
    .b({on_off_pad[0],_al_u3965_o}),
    .c({\u2_Display/n5681 [7],\u2_Display/mux19_b0_sel_is_0_o }),
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({\u2_Display/n5679 ,_al_u3967_o}),
    .f({_al_u3987_o,open_n39007}),
    .q({open_n39011,\u2_Display/i [2]}));  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(0)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*0*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*B)"),
    //.LUTF1("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(0)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*0*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*B)"),
    //.LUTG0("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(1)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*1*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*B)"),
    //.LUTG1("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(1)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*1*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*B)"),
    .INIT_LUTF0(16'b1101110111001111),
    .INIT_LUTF1(16'b1101110111001111),
    .INIT_LUTG0(16'b0001000100000011),
    .INIT_LUTG1(16'b0001000100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3988|_al_u3996  (
    .a({\u2_Display/n2302 ,\u2_Display/n2300 }),
    .b({\u2_Display/mux5_b0_sel_is_0_o ,\u2_Display/mux5_b0_sel_is_0_o }),
    .c({\u2_Display/n2312 [7],\u2_Display/n2312 [9]}),
    .d({\u2_Display/n2310 ,\u2_Display/n2310 }),
    .e({\u2_Display/i [7],\u2_Display/i [9]}),
    .f({_al_u3988_o,_al_u3996_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(0)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*0*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*0*B)"),
    //.LUTF1("~(~A*~((D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0))*~(C)+~A*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*~(C)+~(~A)*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*C+~A*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*C)"),
    //.LUTG0("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(1)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*1*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*1*B)"),
    //.LUTG1("~(~A*~((D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1))*~(C)+~A*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*~(C)+~(~A)*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*C+~A*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*C)"),
    .INIT_LUTF0(16'b1101110111001111),
    .INIT_LUTF1(16'b0000101011111010),
    .INIT_LUTG0(16'b0001000100000011),
    .INIT_LUTG1(16'b0011101000111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3989|_al_u3992  (
    .a({_al_u3988_o,\u2_Display/n2301 }),
    .b({\u2_Display/n4548 ,\u2_Display/mux5_b0_sel_is_0_o }),
    .c({on_off_pad[2],\u2_Display/n2312 [8]}),
    .d({\u2_Display/n4558 [7],\u2_Display/n2310 }),
    .e({\u2_Display/n4556 ,\u2_Display/i [8]}),
    .f({_al_u3989_o,_al_u3992_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u398|_al_u401  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [3],\u2_Display/counta [6]}),
    .d({\u2_Display/n419 [3],\u2_Display/n419 [6]}),
    .f({\u2_Display/n448 ,\u2_Display/n445 }));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~((~C*~B))+A*D*~((~C*~B))+~(A)*D*(~C*~B)+A*D*(~C*~B))"),
    //.LUT1("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .INIT_LUT0(16'b1010101110101000),
    .INIT_LUT1(16'b1010101010111000),
    .MODE("LOGIC"))
    \_al_u3991|_al_u3995  (
    .a({\u2_Display/n5670 ,\u2_Display/n5669 }),
    .b({on_off_pad[0],on_off_pad[0]}),
    .c({\u2_Display/n5681 [8],\u2_Display/n5679 }),
    .d({\u2_Display/n5679 ,\u2_Display/n5681 [9]}),
    .f({_al_u3991_o,_al_u3995_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~((D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0))*~(C)+~A*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*~(C)+~(~A)*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*C+~A*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*C)"),
    //.LUTF1("~(~A*~((D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0))*~(C)+~A*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*~(C)+~(~A)*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*C+~A*(D*~(B)*~(0)+D*B*~(0)+~(D)*B*0+D*B*0)*C)"),
    //.LUTG0("~(~A*~((D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1))*~(C)+~A*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*~(C)+~(~A)*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*C+~A*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*C)"),
    //.LUTG1("~(~A*~((D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1))*~(C)+~A*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*~(C)+~(~A)*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*C+~A*(D*~(B)*~(1)+D*B*~(1)+~(D)*B*1+D*B*1)*C)"),
    .INIT_LUTF0(16'b0000101011111010),
    .INIT_LUTF1(16'b0000101011111010),
    .INIT_LUTG0(16'b0011101000111010),
    .INIT_LUTG1(16'b0011101000111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3993|_al_u3997  (
    .a({_al_u3992_o,_al_u3996_o}),
    .b({\u2_Display/n4547 ,\u2_Display/n4546 }),
    .c({on_off_pad[2],on_off_pad[2]}),
    .d({\u2_Display/n4558 [8],\u2_Display/n4558 [9]}),
    .e({\u2_Display/n4556 ,\u2_Display/n4556 }),
    .f({_al_u3993_o,_al_u3997_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u399|_al_u400  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [4],\u2_Display/counta [5]}),
    .d({\u2_Display/n419 [4],\u2_Display/n419 [5]}),
    .f({\u2_Display/n447 ,\u2_Display/n446 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D)"),
    .INIT_LUT0(16'b0000000011111111),
    .MODE("LOGIC"))
    _al_u4001 (
    .d({open_n39158,\u1_Driver/n4 }),
    .f({open_n39172,vga_hs_pad}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D)"),
    .INIT_LUT0(16'b0000000011111111),
    .MODE("LOGIC"))
    _al_u4002 (
    .d({open_n39186,\u1_Driver/n10 }),
    .f({open_n39200,vga_vs_pad}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D)"),
    .INIT_LUT0(16'b0000000011111111),
    .MODE("LOGIC"))
    _al_u4004 (
    .d({open_n39214,\u2_Display/i [9]}),
    .f({open_n39228,\u2_Display/n140 [0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D)"),
    .INIT_LUT0(16'b0000000011111111),
    .MODE("LOGIC"))
    _al_u4005 (
    .d({open_n39242,\u2_Display/j [9]}),
    .f({open_n39256,\u2_Display/n99 [0]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u402|_al_u404  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [7],\u2_Display/counta [9]}),
    .d({\u2_Display/n419 [7],\u2_Display/n419 [9]}),
    .f({\u2_Display/n444 ,\u2_Display/n442 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u405|_al_u403  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .d({\u2_Display/n419 [10],\u2_Display/n419 [8]}),
    .f({\u2_Display/n441 ,\u2_Display/n443 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u406|_al_u396  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [11],\u2_Display/counta [1]}),
    .d({\u2_Display/n419 [11],\u2_Display/n419 [1]}),
    .f({\u2_Display/n440 ,\u2_Display/n450 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u407|_al_u409  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [12],\u2_Display/counta [14]}),
    .d({\u2_Display/n419 [12],\u2_Display/n419 [14]}),
    .f({\u2_Display/n439 ,\u2_Display/n437 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u408|_al_u412  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [13],\u2_Display/counta [17]}),
    .d({\u2_Display/n419 [13],\u2_Display/n419 [17]}),
    .f({\u2_Display/n438 ,\u2_Display/n434 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u410|_al_u415  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [15],\u2_Display/counta [20]}),
    .d({\u2_Display/n419 [15],\u2_Display/n419 [20]}),
    .f({\u2_Display/n436 ,\u2_Display/n431 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u411|_al_u413  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [16],\u2_Display/counta [18]}),
    .d({\u2_Display/n419 [16],\u2_Display/n419 [18]}),
    .f({\u2_Display/n435 ,\u2_Display/n433 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u414|_al_u417  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [19],\u2_Display/counta [22]}),
    .d({\u2_Display/n419 [19],\u2_Display/n419 [22]}),
    .f({\u2_Display/n432 ,\u2_Display/n429 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u416|_al_u419  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [21],\u2_Display/counta [24]}),
    .d({\u2_Display/n419 [21],\u2_Display/n419 [24]}),
    .f({\u2_Display/n430 ,\u2_Display/n427 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u418|_al_u421  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [23],\u2_Display/counta [26]}),
    .d({\u2_Display/n419 [23],\u2_Display/n419 [26]}),
    .f({\u2_Display/n428 ,\u2_Display/n425 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u420|_al_u424  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [25],\u2_Display/counta [29]}),
    .d({\u2_Display/n419 [25],\u2_Display/n419 [29]}),
    .f({\u2_Display/n426 ,\u2_Display/n422 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u422|_al_u426  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [27],\u2_Display/counta [31]}),
    .d({\u2_Display/n419 [27],\u2_Display/n419 [31]}),
    .f({\u2_Display/n424 ,\u2_Display/n420 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u423|_al_u425  (
    .b({\u2_Display/n417 ,\u2_Display/n417 }),
    .c({\u2_Display/counta [28],\u2_Display/counta [30]}),
    .d({\u2_Display/n419 [28],\u2_Display/n419 [30]}),
    .f({\u2_Display/n423 ,\u2_Display/n421 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u428|_al_u429  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [1],\u2_Display/counta [2]}),
    .d({\u2_Display/n1542 [1],\u2_Display/n1542 [2]}),
    .f({\u2_Display/n1573 ,\u2_Display/n1572 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u430|_al_u431  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [3],\u2_Display/counta [4]}),
    .d({\u2_Display/n1542 [3],\u2_Display/n1542 [4]}),
    .f({\u2_Display/n1571 ,\u2_Display/n1570 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u432|_al_u433  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [5],\u2_Display/counta [6]}),
    .d({\u2_Display/n1542 [5],\u2_Display/n1542 [6]}),
    .f({\u2_Display/n1569 ,\u2_Display/n1568 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u434|_al_u436  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [7],\u2_Display/counta [9]}),
    .d({\u2_Display/n1542 [7],\u2_Display/n1542 [9]}),
    .f({\u2_Display/n1567 ,\u2_Display/n1565 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u437|_al_u435  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .d({\u2_Display/n1542 [10],\u2_Display/n1542 [8]}),
    .f({\u2_Display/n1564 ,\u2_Display/n1566 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u438|_al_u441  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [11],\u2_Display/counta [14]}),
    .d({\u2_Display/n1542 [11],\u2_Display/n1542 [14]}),
    .f({\u2_Display/n1563 ,\u2_Display/n1560 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u440|_al_u444  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [13],\u2_Display/counta [17]}),
    .d({\u2_Display/n1542 [13],\u2_Display/n1542 [17]}),
    .f({\u2_Display/n1561 ,\u2_Display/n1557 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u442|_al_u448  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [15],\u2_Display/counta [21]}),
    .d({\u2_Display/n1542 [15],\u2_Display/n1542 [21]}),
    .f({\u2_Display/n1559 ,\u2_Display/n1553 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u443|_al_u445  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [16],\u2_Display/counta [18]}),
    .d({\u2_Display/n1542 [16],\u2_Display/n1542 [18]}),
    .f({\u2_Display/n1558 ,\u2_Display/n1556 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u446|_al_u452  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [19],\u2_Display/counta [25]}),
    .d({\u2_Display/n1542 [19],\u2_Display/n1542 [25]}),
    .f({\u2_Display/n1555 ,\u2_Display/n1549 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u447|_al_u449  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [20],\u2_Display/counta [22]}),
    .d({\u2_Display/n1542 [20],\u2_Display/n1542 [22]}),
    .f({\u2_Display/n1554 ,\u2_Display/n1552 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u451|_al_u453  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [24],\u2_Display/counta [26]}),
    .d({\u2_Display/n1542 [24],\u2_Display/n1542 [26]}),
    .f({\u2_Display/n1550 ,\u2_Display/n1548 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u459|_al_u461  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [0],\u2_Display/counta [2]}),
    .d({\u2_Display/n2665 [0],\u2_Display/n2665 [2]}),
    .f({\u2_Display/n2697 ,\u2_Display/n2695 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u460 (
    .b({open_n39940,\u2_Display/n2663 }),
    .c({open_n39941,\u2_Display/counta [1]}),
    .d({open_n39944,\u2_Display/n2665 [1]}),
    .f({open_n39962,\u2_Display/n2696 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u462|_al_u465  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [3],\u2_Display/counta [6]}),
    .d({\u2_Display/n2665 [3],\u2_Display/n2665 [6]}),
    .f({\u2_Display/n2694 ,\u2_Display/n2691 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u463|_al_u464  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [4],\u2_Display/counta [5]}),
    .d({\u2_Display/n2665 [4],\u2_Display/n2665 [5]}),
    .f({\u2_Display/n2693 ,\u2_Display/n2692 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u466|_al_u467  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [7],\u2_Display/counta [8]}),
    .d({\u2_Display/n2665 [7],\u2_Display/n2665 [8]}),
    .f({\u2_Display/n2690 ,\u2_Display/n2689 }));
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011111100),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b0011000011111100),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u469|u2_Display/reg4_b0  (
    .b({\u2_Display/n2663 ,\u2_Display/mux19_b0_sel_is_0_o }),
    .c({\u2_Display/counta [10],\u2_Display/counta [0]}),
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({\u2_Display/n2665 [10],_al_u3918_o}),
    .f({\u2_Display/n2687 ,open_n40065}),
    .q({open_n40069,\u2_Display/j [0]}));  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u470|_al_u468  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [11],\u2_Display/counta [9]}),
    .d({\u2_Display/n2665 [11],\u2_Display/n2665 [9]}),
    .f({\u2_Display/n2686 ,\u2_Display/n2688 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u471|_al_u475  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [12],\u2_Display/counta [16]}),
    .d({\u2_Display/n2665 [12],\u2_Display/n2665 [16]}),
    .f({\u2_Display/n2685 ,\u2_Display/n2681 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u472|_al_u473  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [13],\u2_Display/counta [14]}),
    .d({\u2_Display/n2665 [13],\u2_Display/n2665 [14]}),
    .f({\u2_Display/n2684 ,\u2_Display/n2683 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u474|_al_u477  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [15],\u2_Display/counta [18]}),
    .d({\u2_Display/n2665 [15],\u2_Display/n2665 [18]}),
    .f({\u2_Display/n2682 ,\u2_Display/n2679 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u476|_al_u479  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [17],\u2_Display/counta [20]}),
    .d({\u2_Display/n2665 [17],\u2_Display/n2665 [20]}),
    .f({\u2_Display/n2680 ,\u2_Display/n2677 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u478|_al_u481  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [19],\u2_Display/counta [22]}),
    .d({\u2_Display/n2665 [19],\u2_Display/n2665 [22]}),
    .f({\u2_Display/n2678 ,\u2_Display/n2675 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(A*~((0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D))*~(C)+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*~(C)+~(A)*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C+A*(0*~(B)*~(D)+0*B*~(D)+~(0)*B*D+0*B*D)*C)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("~(A*~((1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D))*~(C)+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*~(C)+~(A)*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C+A*(1*~(B)*~(D)+1*B*~(D)+~(1)*B*D+1*B*D)*C)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b0011010111110101),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b0011010100000101),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u480|_al_u3954  (
    .a({open_n40226,_al_u3952_o}),
    .b({\u2_Display/n2663 ,_al_u3953_o}),
    .c({\u2_Display/counta [21],\u2_Display/mux11_b0_sel_is_0_o }),
    .d({\u2_Display/n2665 [21],on_off_pad[4]}),
    .e({open_n40229,\u2_Display/j [9]}),
    .f({\u2_Display/n2676 ,_al_u3954_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u482|_al_u483  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [23],\u2_Display/counta [24]}),
    .d({\u2_Display/n2665 [23],\u2_Display/n2665 [24]}),
    .f({\u2_Display/n2674 ,\u2_Display/n2673 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u484|_al_u485  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [25],\u2_Display/counta [26]}),
    .d({\u2_Display/n2665 [25],\u2_Display/n2665 [26]}),
    .f({\u2_Display/n2672 ,\u2_Display/n2671 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u486|_al_u489  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [27],\u2_Display/counta [30]}),
    .d({\u2_Display/n2665 [27],\u2_Display/n2665 [30]}),
    .f({\u2_Display/n2670 ,\u2_Display/n2667 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u487|_al_u488  (
    .b({\u2_Display/n2663 ,\u2_Display/n2663 }),
    .c({\u2_Display/counta [28],\u2_Display/counta [29]}),
    .d({\u2_Display/n2665 [28],\u2_Display/n2665 [29]}),
    .f({\u2_Display/n2669 ,\u2_Display/n2668 }));
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000100000001),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111000100000001),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u490|u2_Display/reg4_b9  (
    .a({open_n40354,_al_u3954_o}),
    .b({\u2_Display/n2663 ,on_off_pad[1]}),
    .c({\u2_Display/counta [31],on_off_pad[0]}),
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({\u2_Display/n2665 [31],\u2_Display/counta [9]}),
    .f({\u2_Display/n2666 ,open_n40372}),
    .q({open_n40376,\u2_Display/j [9]}));  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTG0("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u491 (
    .c({open_n40381,lcd_data[23]}),
    .d({open_n40384,vga_de_pad}),
    .f({open_n40402,vga_b_pad[0]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~D*C*~B*A)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(1*~D*C*~B*A)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000000000100000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u492|_al_u999  (
    .a({\u1_Driver/n14 ,_al_u998_o}),
    .b({\u1_Driver/n15 ,\u1_Driver/hcnt [6]}),
    .c({\u1_Driver/n17 ,\u1_Driver/hcnt [7]}),
    .d({\u1_Driver/n18 ,\u1_Driver/hcnt [8]}),
    .e({open_n40410,\u1_Driver/hcnt [9]}),
    .f({\u1_Driver/lcd_request ,\u1_Driver/n5 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u493|_al_u502  (
    .c({\u1_Driver/n21 [9],\u1_Driver/n21 [10]}),
    .d({\u1_Driver/lcd_request ,\u1_Driver/lcd_request }),
    .f({lcd_ypos[9],lcd_ypos[10]}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u494|_al_u501  (
    .c({\u1_Driver/n21 [8],\u1_Driver/lcd_request }),
    .d({\u1_Driver/lcd_request ,\u1_Driver/n21 [11]}),
    .f({lcd_ypos[8],lcd_ypos[11]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u495|_al_u498  (
    .c({\u1_Driver/n21 [7],\u1_Driver/n21 [4]}),
    .d({\u1_Driver/lcd_request ,\u1_Driver/lcd_request }),
    .f({lcd_ypos[7],lcd_ypos[4]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u496|_al_u503  (
    .c({\u1_Driver/n21 [6],\u1_Driver/n21 [1]}),
    .d({\u1_Driver/lcd_request ,\u1_Driver/lcd_request }),
    .f({lcd_ypos[6],lcd_ypos[1]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u497|_al_u499  (
    .c({\u1_Driver/n21 [5],\u1_Driver/n21 [3]}),
    .d({\u1_Driver/lcd_request ,\u1_Driver/lcd_request }),
    .f({lcd_ypos[5],lcd_ypos[3]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u500|_al_u504  (
    .c({\u1_Driver/n21 [2],\u1_Driver/n21 [0]}),
    .d({\u1_Driver/lcd_request ,\u1_Driver/lcd_request }),
    .f({lcd_ypos[2],lcd_ypos[0]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u505|_al_u514  (
    .c({\u1_Driver/n20 [9],\u1_Driver/n20 [10]}),
    .d({\u1_Driver/lcd_request ,\u1_Driver/lcd_request }),
    .f({lcd_xpos[9],lcd_xpos[10]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u506|_al_u513  (
    .c({\u1_Driver/n20 [8],\u1_Driver/n20 [11]}),
    .d({\u1_Driver/lcd_request ,\u1_Driver/lcd_request }),
    .f({lcd_xpos[8],lcd_xpos[11]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u507|_al_u509  (
    .c({\u1_Driver/n20 [7],\u1_Driver/n20 [5]}),
    .d({\u1_Driver/lcd_request ,\u1_Driver/lcd_request }),
    .f({lcd_xpos[7],lcd_xpos[5]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u508|_al_u511  (
    .c({\u1_Driver/n20 [6],\u1_Driver/n20 [3]}),
    .d({\u1_Driver/lcd_request ,\u1_Driver/lcd_request }),
    .f({lcd_xpos[6],lcd_xpos[3]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u510|_al_u515  (
    .c({\u1_Driver/n20 [4],\u1_Driver/n20 [1]}),
    .d({\u1_Driver/lcd_request ,\u1_Driver/lcd_request }),
    .f({lcd_xpos[4],lcd_xpos[1]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u512|_al_u516  (
    .c({\u1_Driver/n20 [2],\u1_Driver/n20 [0]}),
    .d({\u1_Driver/lcd_request ,\u1_Driver/lcd_request }),
    .f({lcd_xpos[2],lcd_xpos[0]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u517|_al_u519  (
    .b({\u2_Display/n3823 [0],\u2_Display/n3823 [2]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3820 ,\u2_Display/n3818 }),
    .f({\u2_Display/n3855 ,\u2_Display/n3853 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u518|_al_u522  (
    .b({\u2_Display/n3823 [1],\u2_Display/n3823 [5]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3819 ,\u2_Display/n3815 }),
    .f({\u2_Display/n3854 ,\u2_Display/n3850 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u520|_al_u525  (
    .b({\u2_Display/n3823 [3],\u2_Display/n3823 [8]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3817 ,\u2_Display/n3812 }),
    .f({\u2_Display/n3852 ,\u2_Display/n3847 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u521|_al_u523  (
    .b({\u2_Display/n3823 [4],\u2_Display/n3823 [6]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3816 ,\u2_Display/n3814 }),
    .f({\u2_Display/n3851 ,\u2_Display/n3849 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u524|_al_u527  (
    .b({\u2_Display/n3823 [7],\u2_Display/n3823 [10]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3813 ,\u2_Display/n3810 }),
    .f({\u2_Display/n3848 ,\u2_Display/n3845 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u526|_al_u529  (
    .b({\u2_Display/n3823 [9],\u2_Display/n3823 [12]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3811 ,\u2_Display/n3808 }),
    .f({\u2_Display/n3846 ,\u2_Display/n3843 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u528|_al_u531  (
    .b({\u2_Display/n3823 [11],\u2_Display/n3823 [14]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3809 ,\u2_Display/n3806 }),
    .f({\u2_Display/n3844 ,\u2_Display/n3841 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u530|_al_u533  (
    .b({\u2_Display/n3823 [13],\u2_Display/n3823 [16]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3807 ,\u2_Display/n3804 }),
    .f({\u2_Display/n3842 ,\u2_Display/n3839 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u532|_al_u535  (
    .b({\u2_Display/n3823 [15],\u2_Display/n3823 [18]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3805 ,\u2_Display/n3802 }),
    .f({\u2_Display/n3840 ,\u2_Display/n3837 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u534|_al_u538  (
    .b({\u2_Display/n3823 [17],\u2_Display/n3823 [21]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3803 ,\u2_Display/n3799 }),
    .f({\u2_Display/n3838 ,\u2_Display/n3834 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u536|_al_u541  (
    .b({\u2_Display/n3823 [19],\u2_Display/n3823 [24]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3801 ,\u2_Display/n3796 }),
    .f({\u2_Display/n3836 ,\u2_Display/n3831 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u537|_al_u539  (
    .b({\u2_Display/n3823 [20],\u2_Display/n3823 [22]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3800 ,\u2_Display/n3798 }),
    .f({\u2_Display/n3835 ,\u2_Display/n3833 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u540|_al_u543  (
    .b({\u2_Display/n3823 [23],\u2_Display/n3823 [26]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3797 ,\u2_Display/n3794 }),
    .f({\u2_Display/n3832 ,\u2_Display/n3829 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u542|_al_u545  (
    .b({\u2_Display/n3823 [25],\u2_Display/n3823 [28]}),
    .c({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .d({\u2_Display/n3795 ,\u2_Display/n3792 }),
    .f({\u2_Display/n3830 ,\u2_Display/n3827 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u544|_al_u547  (
    .b({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .c({\u2_Display/n3823 [27],\u2_Display/n3823 [30]}),
    .d({\u2_Display/n3793 ,\u2_Display/n3790 }),
    .f({\u2_Display/n3828 ,\u2_Display/n3825 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTF1("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTG0("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUTG1("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    .INIT_LUTF0(16'b1111101001010000),
    .INIT_LUTF1(16'b1111101001010000),
    .INIT_LUTG0(16'b1111101001010000),
    .INIT_LUTG1(16'b1111101001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u546|_al_u548  (
    .a({\u2_Display/n3821 ,\u2_Display/n3821 }),
    .c({\u2_Display/n3823 [29],\u2_Display/n3823 [31]}),
    .d({\u2_Display/n3791 ,\u2_Display/n3789 }),
    .f({\u2_Display/n3826 ,\u2_Display/n3824 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u549|_al_u551  (
    .b({\u2_Display/n4946 [0],\u2_Display/n4946 [2]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6101 ,\u2_Display/n6099 }),
    .f({\u2_Display/n6136 ,\u2_Display/n6134 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u550|_al_u553  (
    .b({\u2_Display/n4946 [1],\u2_Display/n4946 [4]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6100 ,\u2_Display/n6097 }),
    .f({\u2_Display/n6135 ,\u2_Display/n6132 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u552|_al_u555  (
    .b({\u2_Display/n4946 [3],\u2_Display/n4946 [6]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6098 ,\u2_Display/n6095 }),
    .f({\u2_Display/n6133 ,\u2_Display/n6130 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u554|_al_u557  (
    .b({\u2_Display/n4946 [5],\u2_Display/n4946 [8]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6096 ,\u2_Display/n6093 }),
    .f({\u2_Display/n6131 ,\u2_Display/n6128 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u556|_al_u561  (
    .b({\u2_Display/n4946 [7],\u2_Display/n4946 [12]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6094 ,\u2_Display/n6089 }),
    .f({\u2_Display/n6129 ,\u2_Display/n6124 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u558|_al_u559  (
    .b({\u2_Display/n4946 [9],\u2_Display/n4946 [10]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6092 ,\u2_Display/n6091 }),
    .f({\u2_Display/n6127 ,\u2_Display/n6126 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u560|_al_u563  (
    .b({\u2_Display/n4946 [11],\u2_Display/n4946 [14]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6090 ,\u2_Display/n6087 }),
    .f({\u2_Display/n6125 ,\u2_Display/n6122 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u562|_al_u565  (
    .b({\u2_Display/n4946 [13],\u2_Display/n4946 [16]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6088 ,\u2_Display/n6085 }),
    .f({\u2_Display/n6123 ,\u2_Display/n6120 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u564|_al_u567  (
    .b({\u2_Display/n4946 [15],\u2_Display/n4946 [18]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6086 ,\u2_Display/n6083 }),
    .f({\u2_Display/n6121 ,\u2_Display/n6118 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u566|_al_u569  (
    .b({\u2_Display/n4946 [17],\u2_Display/n4946 [20]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6084 ,\u2_Display/n6081 }),
    .f({\u2_Display/n6119 ,\u2_Display/n6116 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u568|_al_u571  (
    .b({\u2_Display/n4946 [19],\u2_Display/n4946 [22]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6082 ,\u2_Display/n6079 }),
    .f({\u2_Display/n6117 ,\u2_Display/n6114 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u570|_al_u573  (
    .b({\u2_Display/n4946 [21],\u2_Display/n4946 [24]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6080 ,\u2_Display/n6077 }),
    .f({\u2_Display/n6115 ,\u2_Display/n6112 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u572|_al_u575  (
    .b({\u2_Display/n4946 [23],\u2_Display/n4946 [26]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6078 ,\u2_Display/n6075 }),
    .f({\u2_Display/n6113 ,\u2_Display/n6110 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u574|_al_u578  (
    .b({\u2_Display/n4946 [25],\u2_Display/n4946 [29]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6076 ,\u2_Display/n6072 }),
    .f({\u2_Display/n6111 ,\u2_Display/n6107 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u576|_al_u580  (
    .b({\u2_Display/n4946 [27],\u2_Display/n4946 [31]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6074 ,\u2_Display/n6070 }),
    .f({\u2_Display/n6109 ,\u2_Display/n6105 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u577|_al_u579  (
    .b({\u2_Display/n4946 [28],\u2_Display/n4946 [30]}),
    .c({\u2_Display/n4944 ,\u2_Display/n4944 }),
    .d({\u2_Display/n6073 ,\u2_Display/n6071 }),
    .f({\u2_Display/n6108 ,\u2_Display/n6106 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u581|_al_u583  (
    .b({\u2_Display/n454 [0],\u2_Display/n454 [2]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n451 ,\u2_Display/n449 }),
    .f({\u2_Display/n486 ,\u2_Display/n484 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u582|_al_u586  (
    .b({\u2_Display/n454 [1],\u2_Display/n454 [5]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n450 ,\u2_Display/n446 }),
    .f({\u2_Display/n485 ,\u2_Display/n481 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u584|_al_u589  (
    .b({\u2_Display/n454 [3],\u2_Display/n454 [8]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n448 ,\u2_Display/n443 }),
    .f({\u2_Display/n483 ,\u2_Display/n478 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u585|_al_u587  (
    .b({\u2_Display/n454 [4],\u2_Display/n454 [6]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n447 ,\u2_Display/n445 }),
    .f({\u2_Display/n482 ,\u2_Display/n480 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u588|_al_u591  (
    .b({\u2_Display/n454 [7],\u2_Display/n454 [10]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n444 ,\u2_Display/n441 }),
    .f({\u2_Display/n479 ,\u2_Display/n476 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u590|_al_u594  (
    .b({\u2_Display/n454 [9],\u2_Display/n454 [13]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n442 ,\u2_Display/n438 }),
    .f({\u2_Display/n477 ,\u2_Display/n473 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u592|_al_u597  (
    .b({\u2_Display/n454 [11],\u2_Display/n454 [16]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n440 ,\u2_Display/n435 }),
    .f({\u2_Display/n475 ,\u2_Display/n470 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u593|_al_u595  (
    .b({\u2_Display/n454 [12],\u2_Display/n454 [14]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n439 ,\u2_Display/n437 }),
    .f({\u2_Display/n474 ,\u2_Display/n472 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u596|_al_u599  (
    .b({\u2_Display/n454 [15],\u2_Display/n454 [18]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n436 ,\u2_Display/n433 }),
    .f({\u2_Display/n471 ,\u2_Display/n468 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u598|_al_u601  (
    .b({\u2_Display/n454 [17],\u2_Display/n454 [20]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n434 ,\u2_Display/n431 }),
    .f({\u2_Display/n469 ,\u2_Display/n466 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u600|_al_u603  (
    .b({\u2_Display/n454 [19],\u2_Display/n454 [22]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n432 ,\u2_Display/n429 }),
    .f({\u2_Display/n467 ,\u2_Display/n464 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u602|_al_u606  (
    .b({\u2_Display/n454 [21],\u2_Display/n454 [25]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n430 ,\u2_Display/n426 }),
    .f({\u2_Display/n465 ,\u2_Display/n461 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u604|_al_u609  (
    .b({\u2_Display/n454 [23],\u2_Display/n454 [28]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n428 ,\u2_Display/n423 }),
    .f({\u2_Display/n463 ,\u2_Display/n458 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u605|_al_u607  (
    .b({\u2_Display/n454 [24],\u2_Display/n454 [26]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n427 ,\u2_Display/n425 }),
    .f({\u2_Display/n462 ,\u2_Display/n460 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u608|_al_u611  (
    .b({\u2_Display/n454 [27],\u2_Display/n454 [30]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n424 ,\u2_Display/n421 }),
    .f({\u2_Display/n459 ,\u2_Display/n456 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u610|_al_u612  (
    .b({\u2_Display/n454 [29],\u2_Display/n454 [31]}),
    .c({\u2_Display/n452 ,\u2_Display/n452 }),
    .d({\u2_Display/n422 ,\u2_Display/n420 }),
    .f({\u2_Display/n457 ,\u2_Display/n455 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u613|_al_u618  (
    .b({\u2_Display/n1577 [0],\u2_Display/n1577 [5]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1574 ,\u2_Display/n1569 }),
    .f({\u2_Display/n1609 ,\u2_Display/n1604 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u614|_al_u615  (
    .b({\u2_Display/n1577 [1],\u2_Display/n1577 [2]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1573 ,\u2_Display/n1572 }),
    .f({\u2_Display/n1608 ,\u2_Display/n1607 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u616|_al_u621  (
    .b({\u2_Display/n1577 [3],\u2_Display/n1577 [8]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1571 ,\u2_Display/n1566 }),
    .f({\u2_Display/n1606 ,\u2_Display/n1601 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u617|_al_u619  (
    .b({\u2_Display/n1577 [4],\u2_Display/n1577 [6]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1570 ,\u2_Display/n1568 }),
    .f({\u2_Display/n1605 ,\u2_Display/n1603 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u620|_al_u622  (
    .b({\u2_Display/n1577 [7],\u2_Display/n1577 [9]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1567 ,\u2_Display/n1565 }),
    .f({\u2_Display/n1602 ,\u2_Display/n1600 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u623|_al_u625  (
    .b({\u2_Display/n1577 [10],\u2_Display/n1577 [12]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1564 ,\u2_Display/n1562 }),
    .f({\u2_Display/n1599 ,\u2_Display/n1597 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u624|_al_u627  (
    .b({\u2_Display/n1577 [11],\u2_Display/n1577 [14]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1563 ,\u2_Display/n1560 }),
    .f({\u2_Display/n1598 ,\u2_Display/n1595 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u626|_al_u629  (
    .b({\u2_Display/n1577 [13],\u2_Display/n1577 [16]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1561 ,\u2_Display/n1558 }),
    .f({\u2_Display/n1596 ,\u2_Display/n1593 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u628|_al_u631  (
    .b({\u2_Display/n1577 [15],\u2_Display/n1577 [18]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1559 ,\u2_Display/n1556 }),
    .f({\u2_Display/n1594 ,\u2_Display/n1591 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u630|_al_u634  (
    .b({\u2_Display/n1577 [17],\u2_Display/n1577 [21]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1557 ,\u2_Display/n1553 }),
    .f({\u2_Display/n1592 ,\u2_Display/n1588 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u632|_al_u637  (
    .b({\u2_Display/n1577 [19],\u2_Display/n1577 [24]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1555 ,\u2_Display/n1550 }),
    .f({\u2_Display/n1590 ,\u2_Display/n1585 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u633|_al_u635  (
    .b({\u2_Display/n1577 [20],\u2_Display/n1577 [22]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1554 ,\u2_Display/n1552 }),
    .f({\u2_Display/n1589 ,\u2_Display/n1587 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u636|_al_u427  (
    .b({\u2_Display/n1577 [23],\u2_Display/n1540 }),
    .c({\u2_Display/n1575 ,\u2_Display/counta [0]}),
    .d({\u2_Display/n1551 ,\u2_Display/n1542 [0]}),
    .f({\u2_Display/n1586 ,\u2_Display/n1574 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u638|_al_u639  (
    .b({\u2_Display/n1577 [25],\u2_Display/n1577 [26]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1549 ,\u2_Display/n1548 }),
    .f({\u2_Display/n1584 ,\u2_Display/n1583 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u640|_al_u641  (
    .b({\u2_Display/n1577 [27],\u2_Display/n1577 [28]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1547 ,\u2_Display/n1546 }),
    .f({\u2_Display/n1582 ,\u2_Display/n1581 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u642|_al_u643  (
    .b({\u2_Display/n1577 [29],\u2_Display/n1577 [30]}),
    .c({\u2_Display/n1575 ,\u2_Display/n1575 }),
    .d({\u2_Display/n1545 ,\u2_Display/n1544 }),
    .f({\u2_Display/n1580 ,\u2_Display/n1579 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u644|_al_u439  (
    .b({\u2_Display/n1577 [31],\u2_Display/n1540 }),
    .c({\u2_Display/n1575 ,\u2_Display/counta [12]}),
    .d({\u2_Display/n1543 ,\u2_Display/n1542 [12]}),
    .f({\u2_Display/n1578 ,\u2_Display/n1562 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u645|_al_u647  (
    .b({\u2_Display/n2700 [0],\u2_Display/n2700 [2]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2697 ,\u2_Display/n2695 }),
    .f({\u2_Display/n2732 ,\u2_Display/n2730 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u646|_al_u649  (
    .b({\u2_Display/n2700 [1],\u2_Display/n2700 [4]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2696 ,\u2_Display/n2693 }),
    .f({\u2_Display/n2731 ,\u2_Display/n2728 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u648|_al_u651  (
    .b({\u2_Display/n2700 [3],\u2_Display/n2700 [6]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2694 ,\u2_Display/n2691 }),
    .f({\u2_Display/n2729 ,\u2_Display/n2726 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u650|_al_u653  (
    .b({\u2_Display/n2700 [5],\u2_Display/n2700 [8]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2692 ,\u2_Display/n2689 }),
    .f({\u2_Display/n2727 ,\u2_Display/n2724 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u652|_al_u655  (
    .b({\u2_Display/n2700 [7],\u2_Display/n2700 [10]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2690 ,\u2_Display/n2687 }),
    .f({\u2_Display/n2725 ,\u2_Display/n2722 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u654|_al_u658  (
    .b({\u2_Display/n2700 [9],\u2_Display/n2700 [13]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2688 ,\u2_Display/n2684 }),
    .f({\u2_Display/n2723 ,\u2_Display/n2719 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u656|_al_u661  (
    .b({\u2_Display/n2700 [11],\u2_Display/n2700 [16]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2686 ,\u2_Display/n2681 }),
    .f({\u2_Display/n2721 ,\u2_Display/n2716 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u657|_al_u659  (
    .b({\u2_Display/n2700 [12],\u2_Display/n2700 [14]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2685 ,\u2_Display/n2683 }),
    .f({\u2_Display/n2720 ,\u2_Display/n2718 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u660|_al_u663  (
    .b({\u2_Display/n2700 [15],\u2_Display/n2700 [18]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2682 ,\u2_Display/n2679 }),
    .f({\u2_Display/n2717 ,\u2_Display/n2714 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u662|_al_u666  (
    .b({\u2_Display/n2700 [17],\u2_Display/n2700 [21]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2680 ,\u2_Display/n2676 }),
    .f({\u2_Display/n2715 ,\u2_Display/n2711 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u664|_al_u669  (
    .b({\u2_Display/n2700 [19],\u2_Display/n2700 [24]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2678 ,\u2_Display/n2673 }),
    .f({\u2_Display/n2713 ,\u2_Display/n2708 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u665|_al_u667  (
    .b({\u2_Display/n2700 [20],\u2_Display/n2700 [22]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2677 ,\u2_Display/n2675 }),
    .f({\u2_Display/n2712 ,\u2_Display/n2710 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u668|_al_u671  (
    .b({\u2_Display/n2700 [23],\u2_Display/n2700 [26]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2674 ,\u2_Display/n2671 }),
    .f({\u2_Display/n2709 ,\u2_Display/n2706 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u670|_al_u674  (
    .b({\u2_Display/n2700 [25],\u2_Display/n2700 [29]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2672 ,\u2_Display/n2668 }),
    .f({\u2_Display/n2707 ,\u2_Display/n2703 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u672|_al_u676  (
    .b({\u2_Display/n2700 [27],\u2_Display/n2700 [31]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2670 ,\u2_Display/n2666 }),
    .f({\u2_Display/n2705 ,\u2_Display/n2701 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u673|_al_u675  (
    .b({\u2_Display/n2700 [28],\u2_Display/n2700 [30]}),
    .c({\u2_Display/n2698 ,\u2_Display/n2698 }),
    .d({\u2_Display/n2669 ,\u2_Display/n2667 }),
    .f({\u2_Display/n2704 ,\u2_Display/n2702 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u677|_al_u682  (
    .b({\u2_Display/n3858 [0],\u2_Display/n3858 [5]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3855 ,\u2_Display/n3850 }),
    .f({\u2_Display/n3890 ,\u2_Display/n3885 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u678|_al_u679  (
    .b({\u2_Display/n3858 [1],\u2_Display/n3858 [2]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3854 ,\u2_Display/n3853 }),
    .f({\u2_Display/n3889 ,\u2_Display/n3888 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u680|_al_u685  (
    .b({\u2_Display/n3858 [3],\u2_Display/n3858 [8]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3852 ,\u2_Display/n3847 }),
    .f({\u2_Display/n3887 ,\u2_Display/n3882 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u681|_al_u683  (
    .b({\u2_Display/n3858 [4],\u2_Display/n3858 [6]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3851 ,\u2_Display/n3849 }),
    .f({\u2_Display/n3886 ,\u2_Display/n3884 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u684|_al_u687  (
    .b({\u2_Display/n3858 [7],\u2_Display/n3858 [10]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3848 ,\u2_Display/n3845 }),
    .f({\u2_Display/n3883 ,\u2_Display/n3880 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u686|_al_u689  (
    .b({\u2_Display/n3858 [9],\u2_Display/n3858 [12]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3846 ,\u2_Display/n3843 }),
    .f({\u2_Display/n3881 ,\u2_Display/n3878 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u688|_al_u691  (
    .b({\u2_Display/n3858 [11],\u2_Display/n3858 [14]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3844 ,\u2_Display/n3841 }),
    .f({\u2_Display/n3879 ,\u2_Display/n3876 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u690|_al_u693  (
    .b({\u2_Display/n3858 [13],\u2_Display/n3858 [16]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3842 ,\u2_Display/n3839 }),
    .f({\u2_Display/n3877 ,\u2_Display/n3874 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u692|_al_u695  (
    .b({\u2_Display/n3858 [15],\u2_Display/n3858 [18]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3840 ,\u2_Display/n3837 }),
    .f({\u2_Display/n3875 ,\u2_Display/n3872 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u694|_al_u698  (
    .b({\u2_Display/n3858 [17],\u2_Display/n3858 [21]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3838 ,\u2_Display/n3834 }),
    .f({\u2_Display/n3873 ,\u2_Display/n3869 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u696|_al_u702  (
    .b({\u2_Display/n3858 [19],\u2_Display/n3858 [25]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3836 ,\u2_Display/n3830 }),
    .f({\u2_Display/n3871 ,\u2_Display/n3865 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u697|_al_u699  (
    .b({\u2_Display/n3858 [20],\u2_Display/n3858 [22]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3835 ,\u2_Display/n3833 }),
    .f({\u2_Display/n3870 ,\u2_Display/n3868 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u700|_al_u706  (
    .b({\u2_Display/n3858 [23],\u2_Display/n3858 [29]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3832 ,\u2_Display/n3826 }),
    .f({\u2_Display/n3867 ,\u2_Display/n3861 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u701|_al_u703  (
    .b({\u2_Display/n3858 [24],\u2_Display/n3858 [26]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3831 ,\u2_Display/n3829 }),
    .f({\u2_Display/n3866 ,\u2_Display/n3864 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u704|_al_u708  (
    .b({\u2_Display/n3858 [27],\u2_Display/n3858 [31]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3828 ,\u2_Display/n3824 }),
    .f({\u2_Display/n3863 ,\u2_Display/n3859 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u705|_al_u707  (
    .b({\u2_Display/n3858 [28],\u2_Display/n3858 [30]}),
    .c({\u2_Display/n3856 ,\u2_Display/n3856 }),
    .d({\u2_Display/n3827 ,\u2_Display/n3825 }),
    .f({\u2_Display/n3862 ,\u2_Display/n3860 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u709|_al_u714  (
    .b({\u2_Display/n4981 [0],\u2_Display/n4981 [5]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6136 ,\u2_Display/n6131 }),
    .f({\u2_Display/n6171 ,\u2_Display/n6166 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u710|_al_u711  (
    .b({\u2_Display/n4981 [1],\u2_Display/n4981 [2]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6135 ,\u2_Display/n6134 }),
    .f({\u2_Display/n6170 ,\u2_Display/n6169 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u712|_al_u718  (
    .b({\u2_Display/n4981 [3],\u2_Display/n4981 [9]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6133 ,\u2_Display/n6127 }),
    .f({\u2_Display/n6168 ,\u2_Display/n6162 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u713|_al_u715  (
    .b({\u2_Display/n4981 [4],\u2_Display/n4981 [6]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6132 ,\u2_Display/n6130 }),
    .f({\u2_Display/n6167 ,\u2_Display/n6165 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u716|_al_u721  (
    .b({\u2_Display/n4981 [7],\u2_Display/n4981 [12]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6129 ,\u2_Display/n6124 }),
    .f({\u2_Display/n6164 ,\u2_Display/n6159 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u717|_al_u719  (
    .b({\u2_Display/n4981 [8],\u2_Display/n4981 [10]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6128 ,\u2_Display/n6126 }),
    .f({\u2_Display/n6163 ,\u2_Display/n6161 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u720|_al_u723  (
    .b({\u2_Display/n4981 [11],\u2_Display/n4981 [14]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6125 ,\u2_Display/n6122 }),
    .f({\u2_Display/n6160 ,\u2_Display/n6157 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u722|_al_u725  (
    .b({\u2_Display/n4981 [13],\u2_Display/n4981 [16]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6123 ,\u2_Display/n6120 }),
    .f({\u2_Display/n6158 ,\u2_Display/n6155 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u724|_al_u727  (
    .b({\u2_Display/n4981 [15],\u2_Display/n4981 [18]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6121 ,\u2_Display/n6118 }),
    .f({\u2_Display/n6156 ,\u2_Display/n6153 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u726|_al_u730  (
    .b({\u2_Display/n4981 [17],\u2_Display/n4981 [21]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6119 ,\u2_Display/n6115 }),
    .f({\u2_Display/n6154 ,\u2_Display/n6150 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u728|_al_u734  (
    .b({\u2_Display/n4981 [19],\u2_Display/n4981 [25]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6117 ,\u2_Display/n6111 }),
    .f({\u2_Display/n6152 ,\u2_Display/n6146 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u729|_al_u731  (
    .b({\u2_Display/n4981 [20],\u2_Display/n4981 [22]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6116 ,\u2_Display/n6114 }),
    .f({\u2_Display/n6151 ,\u2_Display/n6149 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u732|_al_u738  (
    .b({\u2_Display/n4981 [23],\u2_Display/n4981 [29]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6113 ,\u2_Display/n6107 }),
    .f({\u2_Display/n6148 ,\u2_Display/n6142 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u733|_al_u735  (
    .b({\u2_Display/n4981 [24],\u2_Display/n4981 [26]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6112 ,\u2_Display/n6110 }),
    .f({\u2_Display/n6147 ,\u2_Display/n6145 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u736|_al_u740  (
    .b({\u2_Display/n4981 [27],\u2_Display/n4981 [31]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6109 ,\u2_Display/n6105 }),
    .f({\u2_Display/n6144 ,\u2_Display/n6140 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u737|_al_u739  (
    .b({\u2_Display/n4981 [28],\u2_Display/n4981 [30]}),
    .c({\u2_Display/n4979 ,\u2_Display/n4979 }),
    .d({\u2_Display/n6108 ,\u2_Display/n6106 }),
    .f({\u2_Display/n6143 ,\u2_Display/n6141 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u741|_al_u745  (
    .b({\u2_Display/n489 [0],\u2_Display/n489 [4]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n486 ,\u2_Display/n482 }),
    .f({\u2_Display/n521 ,\u2_Display/n517 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u742|_al_u743  (
    .b({\u2_Display/n489 [1],\u2_Display/n489 [2]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n485 ,\u2_Display/n484 }),
    .f({\u2_Display/n520 ,\u2_Display/n519 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u744|_al_u747  (
    .b({\u2_Display/n489 [3],\u2_Display/n489 [6]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n483 ,\u2_Display/n480 }),
    .f({\u2_Display/n518 ,\u2_Display/n515 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u746|_al_u749  (
    .b({\u2_Display/n489 [5],\u2_Display/n489 [8]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n481 ,\u2_Display/n478 }),
    .f({\u2_Display/n516 ,\u2_Display/n513 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u748|_al_u751  (
    .b({\u2_Display/n489 [7],\u2_Display/n489 [10]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n479 ,\u2_Display/n476 }),
    .f({\u2_Display/n514 ,\u2_Display/n511 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u750|_al_u753  (
    .b({\u2_Display/n489 [9],\u2_Display/n489 [12]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n477 ,\u2_Display/n474 }),
    .f({\u2_Display/n512 ,\u2_Display/n509 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u752|_al_u755  (
    .b({\u2_Display/n489 [11],\u2_Display/n489 [14]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n475 ,\u2_Display/n472 }),
    .f({\u2_Display/n510 ,\u2_Display/n507 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u754|_al_u757  (
    .b({\u2_Display/n489 [13],\u2_Display/n489 [16]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n473 ,\u2_Display/n470 }),
    .f({\u2_Display/n508 ,\u2_Display/n505 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u756|_al_u759  (
    .b({\u2_Display/n489 [15],\u2_Display/n489 [18]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n471 ,\u2_Display/n468 }),
    .f({\u2_Display/n506 ,\u2_Display/n503 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u758|_al_u761  (
    .b({\u2_Display/n489 [17],\u2_Display/n489 [20]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n469 ,\u2_Display/n466 }),
    .f({\u2_Display/n504 ,\u2_Display/n501 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u760|_al_u763  (
    .b({\u2_Display/n489 [19],\u2_Display/n489 [22]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n467 ,\u2_Display/n464 }),
    .f({\u2_Display/n502 ,\u2_Display/n499 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u762|_al_u765  (
    .b({\u2_Display/n489 [21],\u2_Display/n489 [24]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n465 ,\u2_Display/n462 }),
    .f({\u2_Display/n500 ,\u2_Display/n497 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u764|_al_u767  (
    .b({\u2_Display/n489 [23],\u2_Display/n489 [26]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n463 ,\u2_Display/n460 }),
    .f({\u2_Display/n498 ,\u2_Display/n495 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u766|_al_u769  (
    .b({\u2_Display/n489 [25],\u2_Display/n489 [28]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n461 ,\u2_Display/n458 }),
    .f({\u2_Display/n496 ,\u2_Display/n493 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u768|_al_u771  (
    .b({\u2_Display/n489 [27],\u2_Display/n489 [30]}),
    .c({\u2_Display/n487 ,\u2_Display/n487 }),
    .d({\u2_Display/n459 ,\u2_Display/n456 }),
    .f({\u2_Display/n494 ,\u2_Display/n491 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u770|_al_u772  (
    .b({\u2_Display/n489 [29],\u2_Display/n487 }),
    .c({\u2_Display/n487 ,\u2_Display/n489 [31]}),
    .d({\u2_Display/n457 ,\u2_Display/n455 }),
    .f({\u2_Display/n492 ,\u2_Display/n490 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u773|_al_u958  (
    .b({\u2_Display/n1612 [0],\u2_Display/n1647 [25]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1609 ,\u2_Display/n1619 }),
    .f({\u2_Display/n1644 ,\u2_Display/n1654 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u774|_al_u778  (
    .b({\u2_Display/n1612 [1],\u2_Display/n1612 [5]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1608 ,\u2_Display/n1604 }),
    .f({\u2_Display/n1643 ,\u2_Display/n1639 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u775 (
    .b({open_n44151,\u2_Display/n1612 [2]}),
    .c({open_n44152,\u2_Display/n1610 }),
    .d({open_n44155,\u2_Display/n1607 }),
    .f({open_n44173,\u2_Display/n1642 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u776|_al_u781  (
    .b({\u2_Display/n1612 [3],\u2_Display/n1612 [8]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1606 ,\u2_Display/n1601 }),
    .f({\u2_Display/n1641 ,\u2_Display/n1636 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u777|_al_u779  (
    .b({\u2_Display/n1612 [4],\u2_Display/n1612 [6]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1605 ,\u2_Display/n1603 }),
    .f({\u2_Display/n1640 ,\u2_Display/n1638 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u780|_al_u783  (
    .b({\u2_Display/n1612 [7],\u2_Display/n1612 [10]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1602 ,\u2_Display/n1599 }),
    .f({\u2_Display/n1637 ,\u2_Display/n1634 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u782|_al_u785  (
    .b({\u2_Display/n1612 [9],\u2_Display/n1612 [12]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1600 ,\u2_Display/n1597 }),
    .f({\u2_Display/n1635 ,\u2_Display/n1632 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u784|_al_u787  (
    .b({\u2_Display/n1612 [11],\u2_Display/n1612 [14]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1598 ,\u2_Display/n1595 }),
    .f({\u2_Display/n1633 ,\u2_Display/n1630 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u786|_al_u790  (
    .b({\u2_Display/n1612 [13],\u2_Display/n1612 [17]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1596 ,\u2_Display/n1592 }),
    .f({\u2_Display/n1631 ,\u2_Display/n1627 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u788|_al_u794  (
    .b({\u2_Display/n1612 [15],\u2_Display/n1612 [21]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1594 ,\u2_Display/n1588 }),
    .f({\u2_Display/n1629 ,\u2_Display/n1623 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u789|_al_u791  (
    .b({\u2_Display/n1612 [16],\u2_Display/n1612 [18]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1593 ,\u2_Display/n1591 }),
    .f({\u2_Display/n1628 ,\u2_Display/n1626 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u792|_al_u797  (
    .b({\u2_Display/n1612 [19],\u2_Display/n1612 [24]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1590 ,\u2_Display/n1585 }),
    .f({\u2_Display/n1625 ,\u2_Display/n1620 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u793|_al_u795  (
    .b({\u2_Display/n1612 [20],\u2_Display/n1612 [22]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1589 ,\u2_Display/n1587 }),
    .f({\u2_Display/n1624 ,\u2_Display/n1622 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u796|_al_u799  (
    .b({\u2_Display/n1612 [23],\u2_Display/n1612 [26]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1586 ,\u2_Display/n1583 }),
    .f({\u2_Display/n1621 ,\u2_Display/n1618 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u798|_al_u802  (
    .b({\u2_Display/n1612 [25],\u2_Display/n1612 [29]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1584 ,\u2_Display/n1580 }),
    .f({\u2_Display/n1619 ,\u2_Display/n1615 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u800|_al_u804  (
    .b({\u2_Display/n1612 [27],\u2_Display/n1612 [31]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1582 ,\u2_Display/n1578 }),
    .f({\u2_Display/n1617 ,\u2_Display/n1613 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u801|_al_u803  (
    .b({\u2_Display/n1612 [28],\u2_Display/n1612 [30]}),
    .c({\u2_Display/n1610 ,\u2_Display/n1610 }),
    .d({\u2_Display/n1581 ,\u2_Display/n1579 }),
    .f({\u2_Display/n1616 ,\u2_Display/n1614 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u805|_al_u809  (
    .b({\u2_Display/n2735 [0],\u2_Display/n2735 [4]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2732 ,\u2_Display/n2728 }),
    .f({\u2_Display/n2767 ,\u2_Display/n2763 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u806|_al_u807  (
    .b({\u2_Display/n2735 [1],\u2_Display/n2735 [2]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2731 ,\u2_Display/n2730 }),
    .f({\u2_Display/n2766 ,\u2_Display/n2765 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u808|_al_u811  (
    .b({\u2_Display/n2735 [3],\u2_Display/n2735 [6]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2729 ,\u2_Display/n2726 }),
    .f({\u2_Display/n2764 ,\u2_Display/n2761 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u810|_al_u813  (
    .b({\u2_Display/n2735 [5],\u2_Display/n2735 [8]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2727 ,\u2_Display/n2724 }),
    .f({\u2_Display/n2762 ,\u2_Display/n2759 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u812|_al_u815  (
    .b({\u2_Display/n2735 [7],\u2_Display/n2735 [10]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2725 ,\u2_Display/n2722 }),
    .f({\u2_Display/n2760 ,\u2_Display/n2757 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u814|_al_u817  (
    .b({\u2_Display/n2735 [9],\u2_Display/n2735 [12]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2723 ,\u2_Display/n2720 }),
    .f({\u2_Display/n2758 ,\u2_Display/n2755 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u816|_al_u819  (
    .b({\u2_Display/n2735 [11],\u2_Display/n2735 [14]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2721 ,\u2_Display/n2718 }),
    .f({\u2_Display/n2756 ,\u2_Display/n2753 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u818|_al_u822  (
    .b({\u2_Display/n2735 [13],\u2_Display/n2735 [17]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2719 ,\u2_Display/n2715 }),
    .f({\u2_Display/n2754 ,\u2_Display/n2750 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u820|_al_u826  (
    .b({\u2_Display/n2735 [15],\u2_Display/n2735 [21]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2717 ,\u2_Display/n2711 }),
    .f({\u2_Display/n2752 ,\u2_Display/n2746 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u821|_al_u823  (
    .b({\u2_Display/n2735 [16],\u2_Display/n2735 [18]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2716 ,\u2_Display/n2714 }),
    .f({\u2_Display/n2751 ,\u2_Display/n2749 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u824|_al_u830  (
    .b({\u2_Display/n2735 [19],\u2_Display/n2735 [25]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2713 ,\u2_Display/n2707 }),
    .f({\u2_Display/n2748 ,\u2_Display/n2742 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u825|_al_u827  (
    .b({\u2_Display/n2735 [20],\u2_Display/n2735 [22]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2712 ,\u2_Display/n2710 }),
    .f({\u2_Display/n2747 ,\u2_Display/n2745 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u828|_al_u834  (
    .b({\u2_Display/n2735 [23],\u2_Display/n2735 [29]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2709 ,\u2_Display/n2703 }),
    .f({\u2_Display/n2744 ,\u2_Display/n2738 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u829|_al_u831  (
    .b({\u2_Display/n2735 [24],\u2_Display/n2735 [26]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2708 ,\u2_Display/n2706 }),
    .f({\u2_Display/n2743 ,\u2_Display/n2741 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u832|_al_u836  (
    .b({\u2_Display/n2735 [27],\u2_Display/n2735 [31]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2705 ,\u2_Display/n2701 }),
    .f({\u2_Display/n2740 ,\u2_Display/n2736 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u833|_al_u835  (
    .b({\u2_Display/n2735 [28],\u2_Display/n2735 [30]}),
    .c({\u2_Display/n2733 ,\u2_Display/n2733 }),
    .d({\u2_Display/n2704 ,\u2_Display/n2702 }),
    .f({\u2_Display/n2739 ,\u2_Display/n2737 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u837|_al_u839  (
    .b({\u2_Display/n3893 [0],\u2_Display/n3893 [2]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3890 ,\u2_Display/n3888 }),
    .f({\u2_Display/n3925 ,\u2_Display/n3923 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u838|_al_u842  (
    .b({\u2_Display/n3893 [1],\u2_Display/n3893 [5]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3889 ,\u2_Display/n3885 }),
    .f({\u2_Display/n3924 ,\u2_Display/n3920 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u840|_al_u846  (
    .b({\u2_Display/n3893 [3],\u2_Display/n3893 [9]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3887 ,\u2_Display/n3881 }),
    .f({\u2_Display/n3922 ,\u2_Display/n3916 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u841|_al_u843  (
    .b({\u2_Display/n3893 [4],\u2_Display/n3893 [6]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3886 ,\u2_Display/n3884 }),
    .f({\u2_Display/n3921 ,\u2_Display/n3919 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u844|_al_u849  (
    .b({\u2_Display/n3893 [7],\u2_Display/n3893 [12]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3883 ,\u2_Display/n3878 }),
    .f({\u2_Display/n3918 ,\u2_Display/n3913 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u845|_al_u847  (
    .b({\u2_Display/n3893 [8],\u2_Display/n3893 [10]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3882 ,\u2_Display/n3880 }),
    .f({\u2_Display/n3917 ,\u2_Display/n3915 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u848|_al_u851  (
    .b({\u2_Display/n3893 [11],\u2_Display/n3893 [14]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3879 ,\u2_Display/n3876 }),
    .f({\u2_Display/n3914 ,\u2_Display/n3911 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u850|_al_u854  (
    .b({\u2_Display/n3893 [13],\u2_Display/n3893 [17]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3877 ,\u2_Display/n3873 }),
    .f({\u2_Display/n3912 ,\u2_Display/n3908 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u852|_al_u857  (
    .b({\u2_Display/n3893 [15],\u2_Display/n3893 [20]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3875 ,\u2_Display/n3870 }),
    .f({\u2_Display/n3910 ,\u2_Display/n3905 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u853|_al_u855  (
    .b({\u2_Display/n3893 [16],\u2_Display/n3893 [18]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3874 ,\u2_Display/n3872 }),
    .f({\u2_Display/n3909 ,\u2_Display/n3907 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u856|_al_u859  (
    .b({\u2_Display/n3893 [19],\u2_Display/n3893 [22]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3871 ,\u2_Display/n3868 }),
    .f({\u2_Display/n3906 ,\u2_Display/n3903 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u858|_al_u862  (
    .b({\u2_Display/n3893 [21],\u2_Display/n3893 [25]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3869 ,\u2_Display/n3865 }),
    .f({\u2_Display/n3904 ,\u2_Display/n3900 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u860|_al_u866  (
    .b({\u2_Display/n3893 [23],\u2_Display/n3893 [29]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3867 ,\u2_Display/n3861 }),
    .f({\u2_Display/n3902 ,\u2_Display/n3896 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u861|_al_u863  (
    .b({\u2_Display/n3893 [24],\u2_Display/n3893 [26]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3866 ,\u2_Display/n3864 }),
    .f({\u2_Display/n3901 ,\u2_Display/n3899 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u864|_al_u868  (
    .b({\u2_Display/n3893 [27],\u2_Display/n3893 [31]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3863 ,\u2_Display/n3859 }),
    .f({\u2_Display/n3898 ,\u2_Display/n3894 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u865|_al_u867  (
    .b({\u2_Display/n3893 [28],\u2_Display/n3893 [30]}),
    .c({\u2_Display/n3891 ,\u2_Display/n3891 }),
    .d({\u2_Display/n3862 ,\u2_Display/n3860 }),
    .f({\u2_Display/n3897 ,\u2_Display/n3895 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u869|_al_u871  (
    .b({\u2_Display/n5016 [0],\u2_Display/n5016 [2]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6171 ,\u2_Display/n6169 }),
    .f({\u2_Display/n6206 ,\u2_Display/n6204 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u870|_al_u874  (
    .b({\u2_Display/n5016 [1],\u2_Display/n5016 [5]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6170 ,\u2_Display/n6166 }),
    .f({\u2_Display/n6205 ,\u2_Display/n6201 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u872|_al_u878  (
    .b({\u2_Display/n5016 [3],\u2_Display/n5016 [9]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6168 ,\u2_Display/n6162 }),
    .f({\u2_Display/n6203 ,\u2_Display/n6197 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u873|_al_u875  (
    .b({\u2_Display/n5016 [4],\u2_Display/n5016 [6]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6167 ,\u2_Display/n6165 }),
    .f({\u2_Display/n6202 ,\u2_Display/n6200 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u876|_al_u882  (
    .b({\u2_Display/n5016 [7],\u2_Display/n5016 [13]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6164 ,\u2_Display/n6158 }),
    .f({\u2_Display/n6199 ,\u2_Display/n6193 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u877|_al_u879  (
    .b({\u2_Display/n5016 [8],\u2_Display/n5016 [10]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6163 ,\u2_Display/n6161 }),
    .f({\u2_Display/n6198 ,\u2_Display/n6196 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u880|_al_u886  (
    .b({\u2_Display/n5016 [11],\u2_Display/n5016 [17]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6160 ,\u2_Display/n6154 }),
    .f({\u2_Display/n6195 ,\u2_Display/n6189 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u881|_al_u883  (
    .b({\u2_Display/n5016 [12],\u2_Display/n5016 [14]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6159 ,\u2_Display/n6157 }),
    .f({\u2_Display/n6194 ,\u2_Display/n6192 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u884|_al_u889  (
    .b({\u2_Display/n5016 [15],\u2_Display/n5016 [20]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6156 ,\u2_Display/n6151 }),
    .f({\u2_Display/n6191 ,\u2_Display/n6186 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u885|_al_u887  (
    .b({\u2_Display/n5016 [16],\u2_Display/n5016 [18]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6155 ,\u2_Display/n6153 }),
    .f({\u2_Display/n6190 ,\u2_Display/n6188 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u888|_al_u891  (
    .b({\u2_Display/n5016 [19],\u2_Display/n5016 [22]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6152 ,\u2_Display/n6149 }),
    .f({\u2_Display/n6187 ,\u2_Display/n6184 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u890|_al_u893  (
    .b({\u2_Display/n5016 [21],\u2_Display/n5016 [24]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6150 ,\u2_Display/n6147 }),
    .f({\u2_Display/n6185 ,\u2_Display/n6182 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u892|_al_u895  (
    .b({\u2_Display/n5016 [23],\u2_Display/n5016 [26]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6148 ,\u2_Display/n6145 }),
    .f({\u2_Display/n6183 ,\u2_Display/n6180 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u894|_al_u897  (
    .b({\u2_Display/n5016 [25],\u2_Display/n5016 [28]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6146 ,\u2_Display/n6143 }),
    .f({\u2_Display/n6181 ,\u2_Display/n6178 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u896|_al_u899  (
    .b({\u2_Display/n5016 [27],\u2_Display/n5016 [30]}),
    .c({\u2_Display/n5014 ,\u2_Display/n5014 }),
    .d({\u2_Display/n6144 ,\u2_Display/n6141 }),
    .f({\u2_Display/n6179 ,\u2_Display/n6176 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u898|_al_u900  (
    .b({\u2_Display/n5016 [29],\u2_Display/n5014 }),
    .c({\u2_Display/n5014 ,\u2_Display/n5016 [31]}),
    .d({\u2_Display/n6142 ,\u2_Display/n6140 }),
    .f({\u2_Display/n6177 ,\u2_Display/n6175 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u901|_al_u903  (
    .b({\u2_Display/n524 [0],\u2_Display/n524 [2]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n521 ,\u2_Display/n519 }),
    .f({\u2_Display/n556 ,\u2_Display/n554 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u904|_al_u905  (
    .b({\u2_Display/n524 [3],\u2_Display/n524 [4]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n518 ,\u2_Display/n517 }),
    .f({\u2_Display/n553 ,\u2_Display/n552 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u906|_al_u907  (
    .b({\u2_Display/n524 [5],\u2_Display/n524 [6]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n516 ,\u2_Display/n515 }),
    .f({\u2_Display/n551 ,\u2_Display/n550 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u908|_al_u909  (
    .b({\u2_Display/n524 [7],\u2_Display/n524 [8]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n514 ,\u2_Display/n513 }),
    .f({\u2_Display/n549 ,\u2_Display/n548 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u910|_al_u911  (
    .b({\u2_Display/n524 [9],\u2_Display/n524 [10]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n512 ,\u2_Display/n511 }),
    .f({\u2_Display/n547 ,\u2_Display/n546 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u912|_al_u915  (
    .b({\u2_Display/n524 [11],\u2_Display/n524 [14]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n510 ,\u2_Display/n507 }),
    .f({\u2_Display/n545 ,\u2_Display/n542 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u913|_al_u914  (
    .b({\u2_Display/n524 [12],\u2_Display/n524 [13]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n509 ,\u2_Display/n508 }),
    .f({\u2_Display/n544 ,\u2_Display/n543 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u916|_al_u922  (
    .b({\u2_Display/n524 [15],\u2_Display/n524 [21]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n506 ,\u2_Display/n500 }),
    .f({\u2_Display/n541 ,\u2_Display/n535 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u917|_al_u919  (
    .b({\u2_Display/n524 [16],\u2_Display/n524 [18]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n505 ,\u2_Display/n503 }),
    .f({\u2_Display/n540 ,\u2_Display/n538 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u920|_al_u925  (
    .b({\u2_Display/n524 [19],\u2_Display/n524 [24]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n502 ,\u2_Display/n497 }),
    .f({\u2_Display/n537 ,\u2_Display/n532 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u921|_al_u923  (
    .b({\u2_Display/n524 [20],\u2_Display/n524 [22]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n501 ,\u2_Display/n499 }),
    .f({\u2_Display/n536 ,\u2_Display/n534 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u924|_al_u927  (
    .b({\u2_Display/n524 [23],\u2_Display/n524 [26]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n498 ,\u2_Display/n495 }),
    .f({\u2_Display/n533 ,\u2_Display/n530 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u926|_al_u929  (
    .b({\u2_Display/n524 [25],\u2_Display/n524 [28]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n496 ,\u2_Display/n493 }),
    .f({\u2_Display/n531 ,\u2_Display/n528 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u928|_al_u931  (
    .b({\u2_Display/n524 [27],\u2_Display/n524 [30]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n494 ,\u2_Display/n491 }),
    .f({\u2_Display/n529 ,\u2_Display/n526 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u930|_al_u932  (
    .b({\u2_Display/n524 [29],\u2_Display/n524 [31]}),
    .c({\u2_Display/n522 ,\u2_Display/n522 }),
    .d({\u2_Display/n492 ,\u2_Display/n490 }),
    .f({\u2_Display/n527 ,\u2_Display/n525 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"))
    _al_u933 (
    .b({open_n46183,\u2_Display/n1647 [0]}),
    .c({open_n46184,\u2_Display/n1645 }),
    .d({open_n46187,\u2_Display/n1644 }),
    .f({open_n46205,\u2_Display/n1679 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u934|_al_u935  (
    .b({\u2_Display/n1647 [1],\u2_Display/n1647 [2]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1643 ,\u2_Display/n1642 }),
    .f({\u2_Display/n1678 ,\u2_Display/n1677 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u936|_al_u939  (
    .b({\u2_Display/n1647 [3],\u2_Display/n1647 [6]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1641 ,\u2_Display/n1638 }),
    .f({\u2_Display/n1676 ,\u2_Display/n1673 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u937|_al_u938  (
    .b({\u2_Display/n1647 [4],\u2_Display/n1647 [5]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1640 ,\u2_Display/n1639 }),
    .f({\u2_Display/n1675 ,\u2_Display/n1674 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u940|_al_u941  (
    .b({\u2_Display/n1647 [7],\u2_Display/n1647 [8]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1637 ,\u2_Display/n1636 }),
    .f({\u2_Display/n1672 ,\u2_Display/n1671 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u942|_al_u943  (
    .b({\u2_Display/n1647 [9],\u2_Display/n1647 [10]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1635 ,\u2_Display/n1634 }),
    .f({\u2_Display/n1670 ,\u2_Display/n1669 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u944|_al_u947  (
    .b({\u2_Display/n1647 [11],\u2_Display/n1647 [14]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1633 ,\u2_Display/n1630 }),
    .f({\u2_Display/n1668 ,\u2_Display/n1665 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u945|_al_u946  (
    .b({\u2_Display/n1647 [12],\u2_Display/n1647 [13]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1632 ,\u2_Display/n1631 }),
    .f({\u2_Display/n1667 ,\u2_Display/n1666 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u948|_al_u949  (
    .b({\u2_Display/n1647 [15],\u2_Display/n1647 [16]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1629 ,\u2_Display/n1628 }),
    .f({\u2_Display/n1664 ,\u2_Display/n1663 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u950|_al_u951  (
    .b({\u2_Display/n1647 [17],\u2_Display/n1647 [18]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1627 ,\u2_Display/n1626 }),
    .f({\u2_Display/n1662 ,\u2_Display/n1661 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u952|_al_u953  (
    .b({\u2_Display/n1647 [19],\u2_Display/n1647 [20]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1625 ,\u2_Display/n1624 }),
    .f({\u2_Display/n1660 ,\u2_Display/n1659 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u954|_al_u955  (
    .b({\u2_Display/n1647 [21],\u2_Display/n1647 [22]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1623 ,\u2_Display/n1622 }),
    .f({\u2_Display/n1658 ,\u2_Display/n1657 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u956|_al_u961  (
    .b({\u2_Display/n1647 [23],\u2_Display/n1647 [28]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1621 ,\u2_Display/n1616 }),
    .f({\u2_Display/n1656 ,\u2_Display/n1651 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u957|_al_u959  (
    .b({\u2_Display/n1647 [24],\u2_Display/n1647 [26]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1620 ,\u2_Display/n1618 }),
    .f({\u2_Display/n1655 ,\u2_Display/n1653 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u960|_al_u963  (
    .b({\u2_Display/n1647 [27],\u2_Display/n1647 [30]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1617 ,\u2_Display/n1614 }),
    .f({\u2_Display/n1652 ,\u2_Display/n1649 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u962|_al_u964  (
    .b({\u2_Display/n1647 [29],\u2_Display/n1647 [31]}),
    .c({\u2_Display/n1645 ,\u2_Display/n1645 }),
    .d({\u2_Display/n1615 ,\u2_Display/n1613 }),
    .f({\u2_Display/n1650 ,\u2_Display/n1648 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u965|_al_u969  (
    .b({\u2_Display/n2770 [0],\u2_Display/n2770 [4]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2767 ,\u2_Display/n2763 }),
    .f({\u2_Display/n2802 ,\u2_Display/n2798 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u966|_al_u967  (
    .b({\u2_Display/n2770 [1],\u2_Display/n2770 [2]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2766 ,\u2_Display/n2765 }),
    .f({\u2_Display/n2801 ,\u2_Display/n2800 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u968|_al_u971  (
    .b({\u2_Display/n2770 [3],\u2_Display/n2770 [6]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2764 ,\u2_Display/n2761 }),
    .f({\u2_Display/n2799 ,\u2_Display/n2796 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u970|_al_u974  (
    .b({\u2_Display/n2770 [5],\u2_Display/n2770 [9]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2762 ,\u2_Display/n2758 }),
    .f({\u2_Display/n2797 ,\u2_Display/n2793 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u972|_al_u978  (
    .b({\u2_Display/n2770 [7],\u2_Display/n2770 [13]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2760 ,\u2_Display/n2754 }),
    .f({\u2_Display/n2795 ,\u2_Display/n2789 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u973|_al_u975  (
    .b({\u2_Display/n2770 [8],\u2_Display/n2770 [10]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2759 ,\u2_Display/n2757 }),
    .f({\u2_Display/n2794 ,\u2_Display/n2792 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u976|_al_u982  (
    .b({\u2_Display/n2770 [11],\u2_Display/n2770 [17]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2756 ,\u2_Display/n2750 }),
    .f({\u2_Display/n2791 ,\u2_Display/n2785 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u977|_al_u979  (
    .b({\u2_Display/n2770 [12],\u2_Display/n2770 [14]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2755 ,\u2_Display/n2753 }),
    .f({\u2_Display/n2790 ,\u2_Display/n2788 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u980|_al_u985  (
    .b({\u2_Display/n2770 [15],\u2_Display/n2770 [20]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2752 ,\u2_Display/n2747 }),
    .f({\u2_Display/n2787 ,\u2_Display/n2782 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u981|_al_u983  (
    .b({\u2_Display/n2770 [16],\u2_Display/n2770 [18]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2751 ,\u2_Display/n2749 }),
    .f({\u2_Display/n2786 ,\u2_Display/n2784 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u984|_al_u987  (
    .b({\u2_Display/n2770 [19],\u2_Display/n2770 [22]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2748 ,\u2_Display/n2745 }),
    .f({\u2_Display/n2783 ,\u2_Display/n2780 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u986|_al_u989  (
    .b({\u2_Display/n2770 [21],\u2_Display/n2770 [24]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2746 ,\u2_Display/n2743 }),
    .f({\u2_Display/n2781 ,\u2_Display/n2778 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u988|_al_u991  (
    .b({\u2_Display/n2770 [23],\u2_Display/n2770 [26]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2744 ,\u2_Display/n2741 }),
    .f({\u2_Display/n2779 ,\u2_Display/n2776 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u990|_al_u993  (
    .b({\u2_Display/n2770 [25],\u2_Display/n2770 [28]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2742 ,\u2_Display/n2739 }),
    .f({\u2_Display/n2777 ,\u2_Display/n2774 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u992|_al_u995  (
    .b({\u2_Display/n2770 [27],\u2_Display/n2770 [30]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2740 ,\u2_Display/n2737 }),
    .f({\u2_Display/n2775 ,\u2_Display/n2772 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u994|_al_u996  (
    .b({\u2_Display/n2770 [29],\u2_Display/n2770 [31]}),
    .c({\u2_Display/n2768 ,\u2_Display/n2768 }),
    .d({\u2_Display/n2738 ,\u2_Display/n2736 }),
    .f({\u2_Display/n2773 ,\u2_Display/n2771 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*~C*B*A)"),
    //.LUTF1("(~D*B*C*A)"),
    //.LUTG0("(~1*D*~C*B*A)"),
    //.LUTG1("(~D*B*C*A)"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u997|_al_u998  (
    .a({\u1_Driver/hcnt [0],_al_u997_o}),
    .b({\u1_Driver/hcnt [10],\u1_Driver/hcnt [2]}),
    .c({\u1_Driver/hcnt [1],\u1_Driver/hcnt [3]}),
    .d({\u1_Driver/hcnt [11],\u1_Driver/hcnt [4]}),
    .e({open_n47019,\u1_Driver/hcnt [5]}),
    .f({_al_u997_o,_al_u998_o}));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  EG_PHY_GCLK \u0_PLL/uut/bufg_feedback  (
    .clki(\u0_PLL/uut/clk0_buf ),
    .clko(clk_vga));  // al_ip/PLL.v(34)
  EG_PHY_PLL #(
    //.RID("0X0100"),
    //.WID("0X0100"),
    .CLKC0_CPHASE(8),
    .CLKC0_DIV(9),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(1),
    .CLKC1_DIV(1),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_ENABLE("DISABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(1),
    .CLKC2_DIV(1),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("DISABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(1),
    .CLKC3_DIV(1),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("DISABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(9),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("24.000"),
    .FREQ_LOCK_ACCURACY(2),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .REFCLK_DIV(2),
    .REFCLK_SEL("INTERNAL"),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \u0_PLL/uut/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dwe(1'b0),
    .fbclk(clk_vga),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(clk_24m_pad),
    .reset(\u0_PLL/n0 ),
    .stdby(1'b0),
    .clkc({open_n47088,open_n47089,open_n47090,open_n47091,\u0_PLL/uut/clk0_buf }));  // al_ip/PLL.v(57)
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add0/ucin_al_u5013"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add0/u11_al_u5016  (
    .a({open_n47102,\u1_Driver/hcnt [11]}),
    .c(2'b00),
    .d({open_n47107,1'b0}),
    .fci(\u1_Driver/add0/c11 ),
    .f({open_n47124,\u1_Driver/n2 [11]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add0/ucin_al_u5013"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add0/u3_al_u5014  (
    .a({\u1_Driver/hcnt [5],\u1_Driver/hcnt [3]}),
    .b({\u1_Driver/hcnt [6],\u1_Driver/hcnt [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u1_Driver/add0/c3 ),
    .f({\u1_Driver/n2 [5],\u1_Driver/n2 [3]}),
    .fco(\u1_Driver/add0/c7 ),
    .fx({\u1_Driver/n2 [6],\u1_Driver/n2 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add0/ucin_al_u5013"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add0/u7_al_u5015  (
    .a({\u1_Driver/hcnt [9],\u1_Driver/hcnt [7]}),
    .b({\u1_Driver/hcnt [10],\u1_Driver/hcnt [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u1_Driver/add0/c7 ),
    .f({\u1_Driver/n2 [9],\u1_Driver/n2 [7]}),
    .fco(\u1_Driver/add0/c11 ),
    .fx({\u1_Driver/n2 [10],\u1_Driver/n2 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add0/ucin_al_u5013"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add0/ucin_al_u5013  (
    .a({\u1_Driver/hcnt [1],1'b0}),
    .b({\u1_Driver/hcnt [2],\u1_Driver/hcnt [0]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .f({\u1_Driver/n2 [1],open_n47183}),
    .fco(\u1_Driver/add0/c3 ),
    .fx({\u1_Driver/n2 [2],\u1_Driver/n2 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add1/ucin_al_u5017"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add1/u11_al_u5020  (
    .a({open_n47186,\u1_Driver/vcnt [11]}),
    .c(2'b00),
    .d({open_n47191,1'b0}),
    .fci(\u1_Driver/add1/c11 ),
    .f({open_n47208,\u1_Driver/n7 [11]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add1/ucin_al_u5017"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add1/u3_al_u5018  (
    .a({\u1_Driver/vcnt [5],\u1_Driver/vcnt [3]}),
    .b({\u1_Driver/vcnt [6],\u1_Driver/vcnt [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u1_Driver/add1/c3 ),
    .f({\u1_Driver/n7 [5],\u1_Driver/n7 [3]}),
    .fco(\u1_Driver/add1/c7 ),
    .fx({\u1_Driver/n7 [6],\u1_Driver/n7 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add1/ucin_al_u5017"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add1/u7_al_u5019  (
    .a({\u1_Driver/vcnt [9],\u1_Driver/vcnt [7]}),
    .b({\u1_Driver/vcnt [10],\u1_Driver/vcnt [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u1_Driver/add1/c7 ),
    .f({\u1_Driver/n7 [9],\u1_Driver/n7 [7]}),
    .fco(\u1_Driver/add1/c11 ),
    .fx({\u1_Driver/n7 [10],\u1_Driver/n7 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add1/ucin_al_u5017"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add1/ucin_al_u5017  (
    .a({\u1_Driver/vcnt [1],1'b0}),
    .b({\u1_Driver/vcnt [2],\u1_Driver/vcnt [0]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .f({\u1_Driver/n7 [1],open_n47267}),
    .fco(\u1_Driver/add1/c3 ),
    .fx({\u1_Driver/n7 [2],\u1_Driver/n7 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_0|u1_Driver/lt0_cin  (
    .a({\u1_Driver/hcnt [0],1'b0}),
    .b({1'b1,open_n47270}),
    .fco(\u1_Driver/lt0_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_10|u1_Driver/lt0_9  (
    .a(\u1_Driver/hcnt [10:9]),
    .b(2'b11),
    .fci(\u1_Driver/lt0_c9 ),
    .fco(\u1_Driver/lt0_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_2|u1_Driver/lt0_1  (
    .a(\u1_Driver/hcnt [2:1]),
    .b(2'b11),
    .fci(\u1_Driver/lt0_c1 ),
    .fco(\u1_Driver/lt0_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_4|u1_Driver/lt0_3  (
    .a(\u1_Driver/hcnt [4:3]),
    .b(2'b10),
    .fci(\u1_Driver/lt0_c3 ),
    .fco(\u1_Driver/lt0_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_6|u1_Driver/lt0_5  (
    .a(\u1_Driver/hcnt [6:5]),
    .b(2'b00),
    .fci(\u1_Driver/lt0_c5 ),
    .fco(\u1_Driver/lt0_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_8|u1_Driver/lt0_7  (
    .a(\u1_Driver/hcnt [8:7]),
    .b(2'b01),
    .fci(\u1_Driver/lt0_c7 ),
    .fco(\u1_Driver/lt0_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_cout|u1_Driver/lt0_11  (
    .a({1'b0,\u1_Driver/hcnt [11]}),
    .b(2'b10),
    .fci(\u1_Driver/lt0_c11 ),
    .f({\u1_Driver/n1 ,open_n47434}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_0|u1_Driver/lt1_cin  (
    .a({\u1_Driver/hcnt [0],1'b1}),
    .b({1'b1,open_n47440}),
    .fco(\u1_Driver/lt1_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_10|u1_Driver/lt1_9  (
    .a(\u1_Driver/hcnt [10:9]),
    .b(2'b00),
    .fci(\u1_Driver/lt1_c9 ),
    .fco(\u1_Driver/lt1_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_2|u1_Driver/lt1_1  (
    .a(\u1_Driver/hcnt [2:1]),
    .b(2'b11),
    .fci(\u1_Driver/lt1_c1 ),
    .fco(\u1_Driver/lt1_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_4|u1_Driver/lt1_3  (
    .a(\u1_Driver/hcnt [4:3]),
    .b(2'b01),
    .fci(\u1_Driver/lt1_c3 ),
    .fco(\u1_Driver/lt1_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_6|u1_Driver/lt1_5  (
    .a(\u1_Driver/hcnt [6:5]),
    .b(2'b11),
    .fci(\u1_Driver/lt1_c5 ),
    .fco(\u1_Driver/lt1_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_8|u1_Driver/lt1_7  (
    .a(\u1_Driver/hcnt [8:7]),
    .b(2'b00),
    .fci(\u1_Driver/lt1_c7 ),
    .fco(\u1_Driver/lt1_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_cout|u1_Driver/lt1_11  (
    .a({1'b0,\u1_Driver/hcnt [11]}),
    .b(2'b10),
    .fci(\u1_Driver/lt1_c11 ),
    .f({\u1_Driver/n4 ,open_n47604}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_0|u1_Driver/lt2_cin  (
    .a({\u1_Driver/vcnt [0],1'b1}),
    .b({1'b0,open_n47610}),
    .fco(\u1_Driver/lt2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_10|u1_Driver/lt2_9  (
    .a(\u1_Driver/vcnt [10:9]),
    .b(2'b00),
    .fci(\u1_Driver/lt2_c9 ),
    .fco(\u1_Driver/lt2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_2|u1_Driver/lt2_1  (
    .a(\u1_Driver/vcnt [2:1]),
    .b(2'b01),
    .fci(\u1_Driver/lt2_c1 ),
    .fco(\u1_Driver/lt2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_4|u1_Driver/lt2_3  (
    .a(\u1_Driver/vcnt [4:3]),
    .b(2'b00),
    .fci(\u1_Driver/lt2_c3 ),
    .fco(\u1_Driver/lt2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_6|u1_Driver/lt2_5  (
    .a(\u1_Driver/vcnt [6:5]),
    .b(2'b00),
    .fci(\u1_Driver/lt2_c5 ),
    .fco(\u1_Driver/lt2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_8|u1_Driver/lt2_7  (
    .a(\u1_Driver/vcnt [8:7]),
    .b(2'b00),
    .fci(\u1_Driver/lt2_c7 ),
    .fco(\u1_Driver/lt2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_cout|u1_Driver/lt2_11  (
    .a({1'b0,\u1_Driver/vcnt [11]}),
    .b(2'b10),
    .fci(\u1_Driver/lt2_c11 ),
    .f({\u1_Driver/n10 ,open_n47774}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_0|u1_Driver/lt3_cin  (
    .a(2'b01),
    .b({\u1_Driver/hcnt [0],open_n47780}),
    .fco(\u1_Driver/lt3_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_10|u1_Driver/lt3_9  (
    .a(2'b00),
    .b(\u1_Driver/hcnt [10:9]),
    .fci(\u1_Driver/lt3_c9 ),
    .fco(\u1_Driver/lt3_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_2|u1_Driver/lt3_1  (
    .a(2'b00),
    .b(\u1_Driver/hcnt [2:1]),
    .fci(\u1_Driver/lt3_c1 ),
    .fco(\u1_Driver/lt3_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_4|u1_Driver/lt3_3  (
    .a(2'b01),
    .b(\u1_Driver/hcnt [4:3]),
    .fci(\u1_Driver/lt3_c3 ),
    .fco(\u1_Driver/lt3_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_6|u1_Driver/lt3_5  (
    .a(2'b11),
    .b(\u1_Driver/hcnt [6:5]),
    .fci(\u1_Driver/lt3_c5 ),
    .fco(\u1_Driver/lt3_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_8|u1_Driver/lt3_7  (
    .a(2'b10),
    .b(\u1_Driver/hcnt [8:7]),
    .fci(\u1_Driver/lt3_c7 ),
    .fco(\u1_Driver/lt3_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_cout|u1_Driver/lt3_11  (
    .a(2'b00),
    .b({1'b1,\u1_Driver/hcnt [11]}),
    .fci(\u1_Driver/lt3_c11 ),
    .f({\u1_Driver/n11 ,open_n47944}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_0|u1_Driver/lt4_cin  (
    .a({\u1_Driver/hcnt [0],1'b0}),
    .b({1'b0,open_n47950}),
    .fco(\u1_Driver/lt4_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_10|u1_Driver/lt4_9  (
    .a(\u1_Driver/hcnt [10:9]),
    .b(2'b11),
    .fci(\u1_Driver/lt4_c9 ),
    .fco(\u1_Driver/lt4_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_2|u1_Driver/lt4_1  (
    .a(\u1_Driver/hcnt [2:1]),
    .b(2'b00),
    .fci(\u1_Driver/lt4_c1 ),
    .fco(\u1_Driver/lt4_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_4|u1_Driver/lt4_3  (
    .a(\u1_Driver/hcnt [4:3]),
    .b(2'b01),
    .fci(\u1_Driver/lt4_c3 ),
    .fco(\u1_Driver/lt4_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_6|u1_Driver/lt4_5  (
    .a(\u1_Driver/hcnt [6:5]),
    .b(2'b11),
    .fci(\u1_Driver/lt4_c5 ),
    .fco(\u1_Driver/lt4_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_8|u1_Driver/lt4_7  (
    .a(\u1_Driver/hcnt [8:7]),
    .b(2'b00),
    .fci(\u1_Driver/lt4_c7 ),
    .fco(\u1_Driver/lt4_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_cout|u1_Driver/lt4_11  (
    .a({1'b0,\u1_Driver/hcnt [11]}),
    .b(2'b10),
    .fci(\u1_Driver/lt4_c11 ),
    .f({\u1_Driver/n12 ,open_n48114}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_0|u1_Driver/lt5_cin  (
    .a(2'b11),
    .b({\u1_Driver/vcnt [0],open_n48120}),
    .fco(\u1_Driver/lt5_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_10|u1_Driver/lt5_9  (
    .a(2'b00),
    .b(\u1_Driver/vcnt [10:9]),
    .fci(\u1_Driver/lt5_c9 ),
    .fco(\u1_Driver/lt5_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_2|u1_Driver/lt5_1  (
    .a(2'b00),
    .b(\u1_Driver/vcnt [2:1]),
    .fci(\u1_Driver/lt5_c1 ),
    .fco(\u1_Driver/lt5_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_4|u1_Driver/lt5_3  (
    .a(2'b01),
    .b(\u1_Driver/vcnt [4:3]),
    .fci(\u1_Driver/lt5_c3 ),
    .fco(\u1_Driver/lt5_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_6|u1_Driver/lt5_5  (
    .a(2'b01),
    .b(\u1_Driver/vcnt [6:5]),
    .fci(\u1_Driver/lt5_c5 ),
    .fco(\u1_Driver/lt5_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_8|u1_Driver/lt5_7  (
    .a(2'b00),
    .b(\u1_Driver/vcnt [8:7]),
    .fci(\u1_Driver/lt5_c7 ),
    .fco(\u1_Driver/lt5_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_cout|u1_Driver/lt5_11  (
    .a(2'b00),
    .b({1'b1,\u1_Driver/vcnt [11]}),
    .fci(\u1_Driver/lt5_c11 ),
    .f({\u1_Driver/n14 ,open_n48284}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_0|u1_Driver/lt6_cin  (
    .a({\u1_Driver/vcnt [0],1'b0}),
    .b({1'b1,open_n48290}),
    .fco(\u1_Driver/lt6_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_10|u1_Driver/lt6_9  (
    .a(\u1_Driver/vcnt [10:9]),
    .b(2'b10),
    .fci(\u1_Driver/lt6_c9 ),
    .fco(\u1_Driver/lt6_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_2|u1_Driver/lt6_1  (
    .a(\u1_Driver/vcnt [2:1]),
    .b(2'b00),
    .fci(\u1_Driver/lt6_c1 ),
    .fco(\u1_Driver/lt6_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_4|u1_Driver/lt6_3  (
    .a(\u1_Driver/vcnt [4:3]),
    .b(2'b01),
    .fci(\u1_Driver/lt6_c3 ),
    .fco(\u1_Driver/lt6_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_6|u1_Driver/lt6_5  (
    .a(\u1_Driver/vcnt [6:5]),
    .b(2'b01),
    .fci(\u1_Driver/lt6_c5 ),
    .fco(\u1_Driver/lt6_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_8|u1_Driver/lt6_7  (
    .a(\u1_Driver/vcnt [8:7]),
    .b(2'b00),
    .fci(\u1_Driver/lt6_c7 ),
    .fco(\u1_Driver/lt6_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_cout|u1_Driver/lt6_11  (
    .a({1'b0,\u1_Driver/vcnt [11]}),
    .b(2'b10),
    .fci(\u1_Driver/lt6_c11 ),
    .f({\u1_Driver/n15 ,open_n48454}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_0|u1_Driver/lt7_cin  (
    .a(2'b11),
    .b({\u1_Driver/hcnt [0],open_n48460}),
    .fco(\u1_Driver/lt7_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_10|u1_Driver/lt7_9  (
    .a(2'b00),
    .b(\u1_Driver/hcnt [10:9]),
    .fci(\u1_Driver/lt7_c9 ),
    .fco(\u1_Driver/lt7_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_2|u1_Driver/lt7_1  (
    .a(2'b11),
    .b(\u1_Driver/hcnt [2:1]),
    .fci(\u1_Driver/lt7_c1 ),
    .fco(\u1_Driver/lt7_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_4|u1_Driver/lt7_3  (
    .a(2'b00),
    .b(\u1_Driver/hcnt [4:3]),
    .fci(\u1_Driver/lt7_c3 ),
    .fco(\u1_Driver/lt7_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_6|u1_Driver/lt7_5  (
    .a(2'b11),
    .b(\u1_Driver/hcnt [6:5]),
    .fci(\u1_Driver/lt7_c5 ),
    .fco(\u1_Driver/lt7_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_8|u1_Driver/lt7_7  (
    .a(2'b10),
    .b(\u1_Driver/hcnt [8:7]),
    .fci(\u1_Driver/lt7_c7 ),
    .fco(\u1_Driver/lt7_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_cout|u1_Driver/lt7_11  (
    .a(2'b00),
    .b({1'b1,\u1_Driver/hcnt [11]}),
    .fci(\u1_Driver/lt7_c11 ),
    .f({\u1_Driver/n17 ,open_n48624}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_0|u1_Driver/lt8_cin  (
    .a({\u1_Driver/hcnt [0],1'b0}),
    .b({1'b1,open_n48630}),
    .fco(\u1_Driver/lt8_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_10|u1_Driver/lt8_9  (
    .a(\u1_Driver/hcnt [10:9]),
    .b(2'b11),
    .fci(\u1_Driver/lt8_c9 ),
    .fco(\u1_Driver/lt8_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_2|u1_Driver/lt8_1  (
    .a(\u1_Driver/hcnt [2:1]),
    .b(2'b11),
    .fci(\u1_Driver/lt8_c1 ),
    .fco(\u1_Driver/lt8_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_4|u1_Driver/lt8_3  (
    .a(\u1_Driver/hcnt [4:3]),
    .b(2'b00),
    .fci(\u1_Driver/lt8_c3 ),
    .fco(\u1_Driver/lt8_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_6|u1_Driver/lt8_5  (
    .a(\u1_Driver/hcnt [6:5]),
    .b(2'b11),
    .fci(\u1_Driver/lt8_c5 ),
    .fco(\u1_Driver/lt8_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_8|u1_Driver/lt8_7  (
    .a(\u1_Driver/hcnt [8:7]),
    .b(2'b00),
    .fci(\u1_Driver/lt8_c7 ),
    .fco(\u1_Driver/lt8_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_cout|u1_Driver/lt8_11  (
    .a({1'b0,\u1_Driver/hcnt [11]}),
    .b(2'b10),
    .fci(\u1_Driver/lt8_c11 ),
    .f({\u1_Driver/n18 ,open_n48794}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTG0("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b0  (
    .c({open_n48804,\u1_Driver/n7 [0]}),
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d({open_n48805,\u1_Driver/n6_lutinv }),
    .sr(rst_n_pad),
    .q({open_n48827,\u1_Driver/vcnt [0]}));  // source/rtl/Driver.v(78)
  // source/rtl/Driver.v(78)
  // source/rtl/Driver.v(78)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b10|u1_Driver/reg0_b7  (
    .c({\u1_Driver/n7 [10],\u1_Driver/n7 [7]}),
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d({\u1_Driver/n6_lutinv ,\u1_Driver/n6_lutinv }),
    .sr(rst_n_pad),
    .q({\u1_Driver/vcnt [10],\u1_Driver/vcnt [7]}));  // source/rtl/Driver.v(78)
  // source/rtl/Driver.v(78)
  // source/rtl/Driver.v(78)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b1|u1_Driver/reg0_b11  (
    .c({\u1_Driver/n7 [1],\u1_Driver/n7 [11]}),
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d({\u1_Driver/n6_lutinv ,\u1_Driver/n6_lutinv }),
    .sr(rst_n_pad),
    .q({\u1_Driver/vcnt [1],\u1_Driver/vcnt [11]}));  // source/rtl/Driver.v(78)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*C*B*A)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~1*~D*C*B*A)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b2|_al_u1171  (
    .a({open_n48878,_al_u1170_o}),
    .b({open_n48879,\u1_Driver/vcnt [0]}),
    .c({\u1_Driver/n7 [2],\u1_Driver/vcnt [10]}),
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d({\u1_Driver/n6_lutinv ,\u1_Driver/vcnt [2]}),
    .e({open_n48880,\u1_Driver/vcnt [4]}),
    .sr(rst_n_pad),
    .f({open_n48895,_al_u1171_o}),
    .q({\u1_Driver/vcnt [2],open_n48899}));  // source/rtl/Driver.v(78)
  // source/rtl/Driver.v(78)
  // source/rtl/Driver.v(78)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b3|u1_Driver/reg0_b4  (
    .c({\u1_Driver/n7 [3],\u1_Driver/n7 [4]}),
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d({\u1_Driver/n6_lutinv ,\u1_Driver/n6_lutinv }),
    .sr(rst_n_pad),
    .q({\u1_Driver/vcnt [3],\u1_Driver/vcnt [4]}));  // source/rtl/Driver.v(78)
  // source/rtl/Driver.v(78)
  // source/rtl/Driver.v(78)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b5|u1_Driver/reg0_b6  (
    .c({\u1_Driver/n7 [5],\u1_Driver/n7 [6]}),
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d({\u1_Driver/n6_lutinv ,\u1_Driver/n6_lutinv }),
    .sr(rst_n_pad),
    .q({\u1_Driver/vcnt [5],\u1_Driver/vcnt [6]}));  // source/rtl/Driver.v(78)
  // source/rtl/Driver.v(78)
  // source/rtl/Driver.v(78)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b8|u1_Driver/reg0_b9  (
    .c({\u1_Driver/n7 [8],\u1_Driver/n7 [9]}),
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d({\u1_Driver/n6_lutinv ,\u1_Driver/n6_lutinv }),
    .sr(rst_n_pad),
    .q({\u1_Driver/vcnt [8],\u1_Driver/vcnt [9]}));  // source/rtl/Driver.v(78)
  // source/rtl/Driver.v(62)
  // source/rtl/Driver.v(62)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b0|u1_Driver/reg1_b11  (
    .c({\u1_Driver/n1 ,\u1_Driver/n1 }),
    .clk(clk_vga),
    .d({\u1_Driver/n2 [0],\u1_Driver/n2 [11]}),
    .sr(rst_n_pad),
    .q({\u1_Driver/hcnt [0],\u1_Driver/hcnt [11]}));  // source/rtl/Driver.v(62)
  // source/rtl/Driver.v(62)
  // source/rtl/Driver.v(62)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b10|u1_Driver/reg1_b7  (
    .c({\u1_Driver/n1 ,\u1_Driver/n1 }),
    .clk(clk_vga),
    .d({\u1_Driver/n2 [10],\u1_Driver/n2 [7]}),
    .sr(rst_n_pad),
    .q({\u1_Driver/hcnt [10],\u1_Driver/hcnt [7]}));  // source/rtl/Driver.v(62)
  // source/rtl/Driver.v(62)
  // source/rtl/Driver.v(62)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b1|u1_Driver/reg1_b2  (
    .c({\u1_Driver/n1 ,\u1_Driver/n1 }),
    .clk(clk_vga),
    .d({\u1_Driver/n2 [1],\u1_Driver/n2 [2]}),
    .sr(rst_n_pad),
    .q({\u1_Driver/hcnt [1],\u1_Driver/hcnt [2]}));  // source/rtl/Driver.v(62)
  // source/rtl/Driver.v(62)
  // source/rtl/Driver.v(62)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b3|u1_Driver/reg1_b4  (
    .c({\u1_Driver/n1 ,\u1_Driver/n1 }),
    .clk(clk_vga),
    .d({\u1_Driver/n2 [3],\u1_Driver/n2 [4]}),
    .sr(rst_n_pad),
    .q({\u1_Driver/hcnt [3],\u1_Driver/hcnt [4]}));  // source/rtl/Driver.v(62)
  // source/rtl/Driver.v(62)
  // source/rtl/Driver.v(62)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b5|u1_Driver/reg1_b6  (
    .c({\u1_Driver/n1 ,\u1_Driver/n1 }),
    .clk(clk_vga),
    .d({\u1_Driver/n2 [5],\u1_Driver/n2 [6]}),
    .sr(rst_n_pad),
    .q({\u1_Driver/hcnt [5],\u1_Driver/hcnt [6]}));  // source/rtl/Driver.v(62)
  // source/rtl/Driver.v(62)
  // source/rtl/Driver.v(62)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b8|u1_Driver/reg1_b9  (
    .c({\u1_Driver/n1 ,\u1_Driver/n1 }),
    .clk(clk_vga),
    .d({\u1_Driver/n2 [8],\u1_Driver/n2 [9]}),
    .sr(rst_n_pad),
    .q({\u1_Driver/hcnt [8],\u1_Driver/hcnt [9]}));  // source/rtl/Driver.v(62)
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub0/ucin_al_u5021"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub0/u11_al_u5024  (
    .a({open_n49131,\u1_Driver/hcnt [11]}),
    .c(2'b11),
    .d({open_n49136,1'b0}),
    .fci(\u1_Driver/sub0/c11 ),
    .f({open_n49153,\u1_Driver/n20 [11]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub0/ucin_al_u5021"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub0/u3_al_u5022  (
    .a({\u1_Driver/hcnt [5],\u1_Driver/hcnt [3]}),
    .b({\u1_Driver/hcnt [6],\u1_Driver/hcnt [4]}),
    .c(2'b11),
    .d(2'b10),
    .e(2'b10),
    .fci(\u1_Driver/sub0/c3 ),
    .f({\u1_Driver/n20 [5],\u1_Driver/n20 [3]}),
    .fco(\u1_Driver/sub0/c7 ),
    .fx({\u1_Driver/n20 [6],\u1_Driver/n20 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub0/ucin_al_u5021"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub0/u7_al_u5023  (
    .a({\u1_Driver/hcnt [9],\u1_Driver/hcnt [7]}),
    .b({\u1_Driver/hcnt [10],\u1_Driver/hcnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b01),
    .fci(\u1_Driver/sub0/c7 ),
    .f({\u1_Driver/n20 [9],\u1_Driver/n20 [7]}),
    .fco(\u1_Driver/sub0/c11 ),
    .fx({\u1_Driver/n20 [10],\u1_Driver/n20 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub0/ucin_al_u5021"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub0/ucin_al_u5021  (
    .a({\u1_Driver/hcnt [1],1'b0}),
    .b({\u1_Driver/hcnt [2],\u1_Driver/hcnt [0]}),
    .c(2'b11),
    .d(2'b11),
    .e(2'b11),
    .f({\u1_Driver/n20 [1],open_n49212}),
    .fco(\u1_Driver/sub0/c3 ),
    .fx({\u1_Driver/n20 [2],\u1_Driver/n20 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub1/ucin_al_u5025"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub1/u11_al_u5028  (
    .a({open_n49215,\u1_Driver/vcnt [11]}),
    .c(2'b11),
    .d({open_n49220,1'b0}),
    .fci(\u1_Driver/sub1/c11 ),
    .f({open_n49237,\u1_Driver/n21 [11]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub1/ucin_al_u5025"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub1/u3_al_u5026  (
    .a({\u1_Driver/vcnt [5],\u1_Driver/vcnt [3]}),
    .b({\u1_Driver/vcnt [6],\u1_Driver/vcnt [4]}),
    .c(2'b11),
    .d(2'b11),
    .e(2'b00),
    .fci(\u1_Driver/sub1/c3 ),
    .f({\u1_Driver/n21 [5],\u1_Driver/n21 [3]}),
    .fco(\u1_Driver/sub1/c7 ),
    .fx({\u1_Driver/n21 [6],\u1_Driver/n21 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub1/ucin_al_u5025"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub1/u7_al_u5027  (
    .a({\u1_Driver/vcnt [9],\u1_Driver/vcnt [7]}),
    .b({\u1_Driver/vcnt [10],\u1_Driver/vcnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\u1_Driver/sub1/c7 ),
    .f({\u1_Driver/n21 [9],\u1_Driver/n21 [7]}),
    .fco(\u1_Driver/sub1/c11 ),
    .fx({\u1_Driver/n21 [10],\u1_Driver/n21 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub1/ucin_al_u5025"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub1/ucin_al_u5025  (
    .a({\u1_Driver/vcnt [1],1'b0}),
    .b({\u1_Driver/vcnt [2],\u1_Driver/vcnt [0]}),
    .c(2'b11),
    .d(2'b01),
    .e(2'b01),
    .f({\u1_Driver/n21 [1],open_n49296}),
    .fco(\u1_Driver/sub1/c3 ),
    .fx({\u1_Driver/n21 [2],\u1_Driver/n21 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u11_al_u5008  (
    .a({\u2_Display/n [13],\u2_Display/n [11]}),
    .b({\u2_Display/n [14],\u2_Display/n [12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c11 ),
    .f({\u2_Display/n37 [13],\u2_Display/n37 [11]}),
    .fco(\u2_Display/add0/c15 ),
    .fx({\u2_Display/n37 [14],\u2_Display/n37 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u15_al_u5009  (
    .a({\u2_Display/n [17],\u2_Display/n [15]}),
    .b({\u2_Display/n [18],\u2_Display/n [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c15 ),
    .f({\u2_Display/n37 [17],\u2_Display/n37 [15]}),
    .fco(\u2_Display/add0/c19 ),
    .fx({\u2_Display/n37 [18],\u2_Display/n37 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u19_al_u5010  (
    .a({\u2_Display/n [21],\u2_Display/n [19]}),
    .b({\u2_Display/n [22],\u2_Display/n [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c19 ),
    .f({\u2_Display/n37 [21],\u2_Display/n37 [19]}),
    .fco(\u2_Display/add0/c23 ),
    .fx({\u2_Display/n37 [22],\u2_Display/n37 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u23_al_u5011  (
    .a({\u2_Display/n [25],\u2_Display/n [23]}),
    .b({\u2_Display/n [26],\u2_Display/n [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c23 ),
    .f({\u2_Display/n37 [25],\u2_Display/n37 [23]}),
    .fco(\u2_Display/add0/c27 ),
    .fx({\u2_Display/n37 [26],\u2_Display/n37 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u27_al_u5012  (
    .a({\u2_Display/n [29],\u2_Display/n [27]}),
    .b({\u2_Display/n [30],\u2_Display/n [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c27 ),
    .f({\u2_Display/n37 [29],\u2_Display/n37 [27]}),
    .fx({\u2_Display/n37 [30],\u2_Display/n37 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u3_al_u5006  (
    .a({\u2_Display/n [5],\u2_Display/n [3]}),
    .b({\u2_Display/n [6],\u2_Display/n [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c3 ),
    .f({\u2_Display/n37 [5],\u2_Display/n37 [3]}),
    .fco(\u2_Display/add0/c7 ),
    .fx({\u2_Display/n37 [6],\u2_Display/n37 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u7_al_u5007  (
    .a({\u2_Display/n [9],\u2_Display/n [7]}),
    .b({\u2_Display/n [10],\u2_Display/n [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c7 ),
    .f({\u2_Display/n37 [9],\u2_Display/n37 [7]}),
    .fco(\u2_Display/add0/c11 ),
    .fx({\u2_Display/n37 [10],\u2_Display/n37 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/add0/ucin_al_u5005  (
    .a({\u2_Display/n [1],1'b0}),
    .b({\u2_Display/n [2],\u2_Display/n [0]}),
    .c(2'b00),
    .clk(clk_vga),
    .d(2'b01),
    .e(2'b01),
    .mi(\u2_Display/n37 [5:4]),
    .sr(\u2_Display/n35 ),
    .f({\u2_Display/n37 [1],open_n49439}),
    .fco(\u2_Display/add0/c3 ),
    .fx({\u2_Display/n37 [2],\u2_Display/n37 [0]}),
    .q(\u2_Display/n [5:4]));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u11_al_u4009  (
    .a({\u2_Display/counta [13],\u2_Display/counta [11]}),
    .b({\u2_Display/counta [14],\u2_Display/counta [12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c11 ),
    .f({\u2_Display/n41 [13],\u2_Display/n41 [11]}),
    .fco(\u2_Display/add1/c15 ),
    .fx({\u2_Display/n41 [14],\u2_Display/n41 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u15_al_u4010  (
    .a({\u2_Display/counta [17],\u2_Display/counta [15]}),
    .b({\u2_Display/counta [18],\u2_Display/counta [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c15 ),
    .f({\u2_Display/n41 [17],\u2_Display/n41 [15]}),
    .fco(\u2_Display/add1/c19 ),
    .fx({\u2_Display/n41 [18],\u2_Display/n41 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u19_al_u4011  (
    .a({\u2_Display/counta [21],\u2_Display/counta [19]}),
    .b({\u2_Display/counta [22],\u2_Display/counta [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c19 ),
    .f({\u2_Display/n41 [21],\u2_Display/n41 [19]}),
    .fco(\u2_Display/add1/c23 ),
    .fx({\u2_Display/n41 [22],\u2_Display/n41 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u23_al_u4012  (
    .a({\u2_Display/counta [25],\u2_Display/counta [23]}),
    .b({\u2_Display/counta [26],\u2_Display/counta [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c23 ),
    .f({\u2_Display/n41 [25],\u2_Display/n41 [23]}),
    .fco(\u2_Display/add1/c27 ),
    .fx({\u2_Display/n41 [26],\u2_Display/n41 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u27_al_u4013  (
    .a({\u2_Display/counta [29],\u2_Display/counta [27]}),
    .b({\u2_Display/counta [30],\u2_Display/counta [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c27 ),
    .f({\u2_Display/n41 [29],\u2_Display/n41 [27]}),
    .fco(\u2_Display/add1/c31 ),
    .fx({\u2_Display/n41 [30],\u2_Display/n41 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u31_al_u4014  (
    .a({open_n49530,\u2_Display/counta [31]}),
    .c(2'b00),
    .d({open_n49535,1'b0}),
    .fci(\u2_Display/add1/c31 ),
    .f({open_n49552,\u2_Display/n41 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u3_al_u4007  (
    .a({\u2_Display/counta [5],\u2_Display/counta [3]}),
    .b({\u2_Display/counta [6],\u2_Display/counta [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c3 ),
    .f({\u2_Display/n41 [5],\u2_Display/n41 [3]}),
    .fco(\u2_Display/add1/c7 ),
    .fx({\u2_Display/n41 [6],\u2_Display/n41 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u7_al_u4008  (
    .a({\u2_Display/counta [9],\u2_Display/counta [7]}),
    .b({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c7 ),
    .f({\u2_Display/n41 [9],\u2_Display/n41 [7]}),
    .fco(\u2_Display/add1/c11 ),
    .fx({\u2_Display/n41 [10],\u2_Display/n41 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/add1/ucin_al_u4006  (
    .a({\u2_Display/counta [1],1'b0}),
    .b({\u2_Display/counta [2],\u2_Display/counta [0]}),
    .c(2'b00),
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d(2'b01),
    .e(2'b01),
    .mi(\u2_Display/n41 [6:5]),
    .f({\u2_Display/n41 [1],open_n49607}),
    .fco(\u2_Display/add1/c3 ),
    .fx({\u2_Display/n41 [2],\u2_Display/n41 [0]}),
    .q(\u2_Display/counta [6:5]));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u11_al_u4018  (
    .a({\u2_Display/n3209 ,\u2_Display/n3211 }),
    .b({\u2_Display/n3208 ,\u2_Display/n3210 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add100/c11 ),
    .f({\u2_Display/n3225 [13],\u2_Display/n3225 [11]}),
    .fco(\u2_Display/add100/c15 ),
    .fx({\u2_Display/n3225 [14],\u2_Display/n3225 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u15_al_u4019  (
    .a({\u2_Display/n3205 ,\u2_Display/n3207 }),
    .b({\u2_Display/n3204 ,\u2_Display/n3206 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add100/c15 ),
    .f({\u2_Display/n3225 [17],\u2_Display/n3225 [15]}),
    .fco(\u2_Display/add100/c19 ),
    .fx({\u2_Display/n3225 [18],\u2_Display/n3225 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u19_al_u4020  (
    .a({\u2_Display/n3201 ,\u2_Display/n3203 }),
    .b({\u2_Display/n3200 ,\u2_Display/n3202 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add100/c19 ),
    .f({\u2_Display/n3225 [21],\u2_Display/n3225 [19]}),
    .fco(\u2_Display/add100/c23 ),
    .fx({\u2_Display/n3225 [22],\u2_Display/n3225 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u23_al_u4021  (
    .a({\u2_Display/n3197 ,\u2_Display/n3199 }),
    .b({\u2_Display/n3196 ,\u2_Display/n3198 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add100/c23 ),
    .f({\u2_Display/n3225 [25],\u2_Display/n3225 [23]}),
    .fco(\u2_Display/add100/c27 ),
    .fx({\u2_Display/n3225 [26],\u2_Display/n3225 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u27_al_u4022  (
    .a({\u2_Display/n3193 ,\u2_Display/n3195 }),
    .b({\u2_Display/n3192 ,\u2_Display/n3194 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add100/c27 ),
    .f({\u2_Display/n3225 [29],\u2_Display/n3225 [27]}),
    .fco(\u2_Display/add100/c31 ),
    .fx({\u2_Display/n3225 [30],\u2_Display/n3225 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u31_al_u4023  (
    .a({open_n49698,\u2_Display/n3191 }),
    .c(2'b00),
    .d({open_n49703,1'b1}),
    .fci(\u2_Display/add100/c31 ),
    .f({open_n49720,\u2_Display/n3225 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u3_al_u4016  (
    .a({\u2_Display/n3217 ,\u2_Display/n3219 }),
    .b({\u2_Display/n3216 ,\u2_Display/n3218 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add100/c3 ),
    .f({\u2_Display/n3225 [5],\u2_Display/n3225 [3]}),
    .fco(\u2_Display/add100/c7 ),
    .fx({\u2_Display/n3225 [6],\u2_Display/n3225 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u7_al_u4017  (
    .a({\u2_Display/n3213 ,\u2_Display/n3215 }),
    .b({\u2_Display/n3212 ,\u2_Display/n3214 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add100/c7 ),
    .f({\u2_Display/n3225 [9],\u2_Display/n3225 [7]}),
    .fco(\u2_Display/add100/c11 ),
    .fx({\u2_Display/n3225 [10],\u2_Display/n3225 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/ucin_al_u4015  (
    .a({\u2_Display/n3221 ,1'b1}),
    .b({\u2_Display/n3220 ,\u2_Display/n3222 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3225 [1],open_n49779}),
    .fco(\u2_Display/add100/c3 ),
    .fx({\u2_Display/n3225 [2],\u2_Display/n3225 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u11_al_u4027  (
    .a({\u2_Display/n3244 ,\u2_Display/n3246 }),
    .b({\u2_Display/n3243 ,\u2_Display/n3245 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add101/c11 ),
    .f({\u2_Display/n3260 [13],\u2_Display/n3260 [11]}),
    .fco(\u2_Display/add101/c15 ),
    .fx({\u2_Display/n3260 [14],\u2_Display/n3260 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u15_al_u4028  (
    .a({\u2_Display/n3240 ,\u2_Display/n3242 }),
    .b({\u2_Display/n3239 ,\u2_Display/n3241 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add101/c15 ),
    .f({\u2_Display/n3260 [17],\u2_Display/n3260 [15]}),
    .fco(\u2_Display/add101/c19 ),
    .fx({\u2_Display/n3260 [18],\u2_Display/n3260 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u19_al_u4029  (
    .a({\u2_Display/n3236 ,\u2_Display/n3238 }),
    .b({\u2_Display/n3235 ,\u2_Display/n3237 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add101/c19 ),
    .f({\u2_Display/n3260 [21],\u2_Display/n3260 [19]}),
    .fco(\u2_Display/add101/c23 ),
    .fx({\u2_Display/n3260 [22],\u2_Display/n3260 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u23_al_u4030  (
    .a({\u2_Display/n3232 ,\u2_Display/n3234 }),
    .b({\u2_Display/n3231 ,\u2_Display/n3233 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add101/c23 ),
    .f({\u2_Display/n3260 [25],\u2_Display/n3260 [23]}),
    .fco(\u2_Display/add101/c27 ),
    .fx({\u2_Display/n3260 [26],\u2_Display/n3260 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u27_al_u4031  (
    .a({\u2_Display/n3228 ,\u2_Display/n3230 }),
    .b({\u2_Display/n3227 ,\u2_Display/n3229 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add101/c27 ),
    .f({\u2_Display/n3260 [29],\u2_Display/n3260 [27]}),
    .fco(\u2_Display/add101/c31 ),
    .fx({\u2_Display/n3260 [30],\u2_Display/n3260 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u31_al_u4032  (
    .a({open_n49872,\u2_Display/n3226 }),
    .c(2'b00),
    .d({open_n49877,1'b1}),
    .fci(\u2_Display/add101/c31 ),
    .f({open_n49894,\u2_Display/n3260 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u3_al_u4025  (
    .a({\u2_Display/n3252 ,\u2_Display/n3254 }),
    .b({\u2_Display/n3251 ,\u2_Display/n3253 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add101/c3 ),
    .f({\u2_Display/n3260 [5],\u2_Display/n3260 [3]}),
    .fco(\u2_Display/add101/c7 ),
    .fx({\u2_Display/n3260 [6],\u2_Display/n3260 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u7_al_u4026  (
    .a({\u2_Display/n3248 ,\u2_Display/n3250 }),
    .b({\u2_Display/n3247 ,\u2_Display/n3249 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add101/c7 ),
    .f({\u2_Display/n3260 [9],\u2_Display/n3260 [7]}),
    .fco(\u2_Display/add101/c11 ),
    .fx({\u2_Display/n3260 [10],\u2_Display/n3260 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/ucin_al_u4024  (
    .a({\u2_Display/n3256 ,1'b1}),
    .b({\u2_Display/n3255 ,\u2_Display/n3257 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3260 [1],open_n49953}),
    .fco(\u2_Display/add101/c3 ),
    .fx({\u2_Display/n3260 [2],\u2_Display/n3260 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u11_al_u4036  (
    .a({\u2_Display/n3279 ,\u2_Display/n3281 }),
    .b({\u2_Display/n3278 ,\u2_Display/n3280 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add102/c11 ),
    .f({\u2_Display/n3295 [13],\u2_Display/n3295 [11]}),
    .fco(\u2_Display/add102/c15 ),
    .fx({\u2_Display/n3295 [14],\u2_Display/n3295 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u15_al_u4037  (
    .a({\u2_Display/n3275 ,\u2_Display/n3277 }),
    .b({\u2_Display/n3274 ,\u2_Display/n3276 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add102/c15 ),
    .f({\u2_Display/n3295 [17],\u2_Display/n3295 [15]}),
    .fco(\u2_Display/add102/c19 ),
    .fx({\u2_Display/n3295 [18],\u2_Display/n3295 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u19_al_u4038  (
    .a({\u2_Display/n3271 ,\u2_Display/n3273 }),
    .b({\u2_Display/n3270 ,\u2_Display/n3272 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add102/c19 ),
    .f({\u2_Display/n3295 [21],\u2_Display/n3295 [19]}),
    .fco(\u2_Display/add102/c23 ),
    .fx({\u2_Display/n3295 [22],\u2_Display/n3295 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u23_al_u4039  (
    .a({\u2_Display/n3267 ,\u2_Display/n3269 }),
    .b({\u2_Display/n3266 ,\u2_Display/n3268 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add102/c23 ),
    .f({\u2_Display/n3295 [25],\u2_Display/n3295 [23]}),
    .fco(\u2_Display/add102/c27 ),
    .fx({\u2_Display/n3295 [26],\u2_Display/n3295 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u27_al_u4040  (
    .a({\u2_Display/n3263 ,\u2_Display/n3265 }),
    .b({\u2_Display/n3262 ,\u2_Display/n3264 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add102/c27 ),
    .f({\u2_Display/n3295 [29],\u2_Display/n3295 [27]}),
    .fco(\u2_Display/add102/c31 ),
    .fx({\u2_Display/n3295 [30],\u2_Display/n3295 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u31_al_u4041  (
    .a({open_n50046,\u2_Display/n3261 }),
    .c(2'b00),
    .d({open_n50051,1'b1}),
    .fci(\u2_Display/add102/c31 ),
    .f({open_n50068,\u2_Display/n3295 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u3_al_u4034  (
    .a({\u2_Display/n3287 ,\u2_Display/n3289 }),
    .b({\u2_Display/n3286 ,\u2_Display/n3288 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add102/c3 ),
    .f({\u2_Display/n3295 [5],\u2_Display/n3295 [3]}),
    .fco(\u2_Display/add102/c7 ),
    .fx({\u2_Display/n3295 [6],\u2_Display/n3295 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u7_al_u4035  (
    .a({\u2_Display/n3283 ,\u2_Display/n3285 }),
    .b({\u2_Display/n3282 ,\u2_Display/n3284 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b00),
    .fci(\u2_Display/add102/c7 ),
    .f({\u2_Display/n3295 [9],\u2_Display/n3295 [7]}),
    .fco(\u2_Display/add102/c11 ),
    .fx({\u2_Display/n3295 [10],\u2_Display/n3295 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/ucin_al_u4033  (
    .a({\u2_Display/n3291 ,1'b1}),
    .b({\u2_Display/n3290 ,\u2_Display/n3292 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3295 [1],open_n50127}),
    .fco(\u2_Display/add102/c3 ),
    .fx({\u2_Display/n3295 [2],\u2_Display/n3295 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u11_al_u4045  (
    .a({\u2_Display/n3314 ,\u2_Display/n3316 }),
    .b({\u2_Display/n3313 ,\u2_Display/n3315 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add103/c11 ),
    .f({\u2_Display/n3330 [13],\u2_Display/n3330 [11]}),
    .fco(\u2_Display/add103/c15 ),
    .fx({\u2_Display/n3330 [14],\u2_Display/n3330 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u15_al_u4046  (
    .a({\u2_Display/n3310 ,\u2_Display/n3312 }),
    .b({\u2_Display/n3309 ,\u2_Display/n3311 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add103/c15 ),
    .f({\u2_Display/n3330 [17],\u2_Display/n3330 [15]}),
    .fco(\u2_Display/add103/c19 ),
    .fx({\u2_Display/n3330 [18],\u2_Display/n3330 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u19_al_u4047  (
    .a({\u2_Display/n3306 ,\u2_Display/n3308 }),
    .b({\u2_Display/n3305 ,\u2_Display/n3307 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add103/c19 ),
    .f({\u2_Display/n3330 [21],\u2_Display/n3330 [19]}),
    .fco(\u2_Display/add103/c23 ),
    .fx({\u2_Display/n3330 [22],\u2_Display/n3330 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u23_al_u4048  (
    .a({\u2_Display/n3302 ,\u2_Display/n3304 }),
    .b({\u2_Display/n3301 ,\u2_Display/n3303 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add103/c23 ),
    .f({\u2_Display/n3330 [25],\u2_Display/n3330 [23]}),
    .fco(\u2_Display/add103/c27 ),
    .fx({\u2_Display/n3330 [26],\u2_Display/n3330 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u27_al_u4049  (
    .a({\u2_Display/n3298 ,\u2_Display/n3300 }),
    .b({\u2_Display/n3297 ,\u2_Display/n3299 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add103/c27 ),
    .f({\u2_Display/n3330 [29],\u2_Display/n3330 [27]}),
    .fco(\u2_Display/add103/c31 ),
    .fx({\u2_Display/n3330 [30],\u2_Display/n3330 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u31_al_u4050  (
    .a({open_n50220,\u2_Display/n3296 }),
    .c(2'b00),
    .d({open_n50225,1'b1}),
    .fci(\u2_Display/add103/c31 ),
    .f({open_n50242,\u2_Display/n3330 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u3_al_u4043  (
    .a({\u2_Display/n3322 ,\u2_Display/n3324 }),
    .b({\u2_Display/n3321 ,\u2_Display/n3323 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add103/c3 ),
    .f({\u2_Display/n3330 [5],\u2_Display/n3330 [3]}),
    .fco(\u2_Display/add103/c7 ),
    .fx({\u2_Display/n3330 [6],\u2_Display/n3330 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u7_al_u4044  (
    .a({\u2_Display/n3318 ,\u2_Display/n3320 }),
    .b({\u2_Display/n3317 ,\u2_Display/n3319 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add103/c7 ),
    .f({\u2_Display/n3330 [9],\u2_Display/n3330 [7]}),
    .fco(\u2_Display/add103/c11 ),
    .fx({\u2_Display/n3330 [10],\u2_Display/n3330 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/ucin_al_u4042  (
    .a({\u2_Display/n3326 ,1'b1}),
    .b({\u2_Display/n3325 ,\u2_Display/n3327 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3330 [1],open_n50301}),
    .fco(\u2_Display/add103/c3 ),
    .fx({\u2_Display/n3330 [2],\u2_Display/n3330 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u11_al_u4054  (
    .a({\u2_Display/n3349 ,\u2_Display/n3351 }),
    .b({\u2_Display/n3348 ,\u2_Display/n3350 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add104/c11 ),
    .f({\u2_Display/n3365 [13],\u2_Display/n3365 [11]}),
    .fco(\u2_Display/add104/c15 ),
    .fx({\u2_Display/n3365 [14],\u2_Display/n3365 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u15_al_u4055  (
    .a({\u2_Display/n3345 ,\u2_Display/n3347 }),
    .b({\u2_Display/n3344 ,\u2_Display/n3346 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add104/c15 ),
    .f({\u2_Display/n3365 [17],\u2_Display/n3365 [15]}),
    .fco(\u2_Display/add104/c19 ),
    .fx({\u2_Display/n3365 [18],\u2_Display/n3365 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u19_al_u4056  (
    .a({\u2_Display/n3341 ,\u2_Display/n3343 }),
    .b({\u2_Display/n3340 ,\u2_Display/n3342 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add104/c19 ),
    .f({\u2_Display/n3365 [21],\u2_Display/n3365 [19]}),
    .fco(\u2_Display/add104/c23 ),
    .fx({\u2_Display/n3365 [22],\u2_Display/n3365 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u23_al_u4057  (
    .a({\u2_Display/n3337 ,\u2_Display/n3339 }),
    .b({\u2_Display/n3336 ,\u2_Display/n3338 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add104/c23 ),
    .f({\u2_Display/n3365 [25],\u2_Display/n3365 [23]}),
    .fco(\u2_Display/add104/c27 ),
    .fx({\u2_Display/n3365 [26],\u2_Display/n3365 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u27_al_u4058  (
    .a({\u2_Display/n3333 ,\u2_Display/n3335 }),
    .b({\u2_Display/n3332 ,\u2_Display/n3334 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add104/c27 ),
    .f({\u2_Display/n3365 [29],\u2_Display/n3365 [27]}),
    .fco(\u2_Display/add104/c31 ),
    .fx({\u2_Display/n3365 [30],\u2_Display/n3365 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u31_al_u4059  (
    .a({open_n50394,\u2_Display/n3331 }),
    .c(2'b00),
    .d({open_n50399,1'b1}),
    .fci(\u2_Display/add104/c31 ),
    .f({open_n50416,\u2_Display/n3365 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u3_al_u4052  (
    .a({\u2_Display/n3357 ,\u2_Display/n3359 }),
    .b({\u2_Display/n3356 ,\u2_Display/n3358 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add104/c3 ),
    .f({\u2_Display/n3365 [5],\u2_Display/n3365 [3]}),
    .fco(\u2_Display/add104/c7 ),
    .fx({\u2_Display/n3365 [6],\u2_Display/n3365 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u7_al_u4053  (
    .a({\u2_Display/n3353 ,\u2_Display/n3355 }),
    .b({\u2_Display/n3352 ,\u2_Display/n3354 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add104/c7 ),
    .f({\u2_Display/n3365 [9],\u2_Display/n3365 [7]}),
    .fco(\u2_Display/add104/c11 ),
    .fx({\u2_Display/n3365 [10],\u2_Display/n3365 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/ucin_al_u4051  (
    .a({\u2_Display/n3361 ,1'b1}),
    .b({\u2_Display/n3360 ,\u2_Display/n3362 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3365 [1],open_n50475}),
    .fco(\u2_Display/add104/c3 ),
    .fx({\u2_Display/n3365 [2],\u2_Display/n3365 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u11_al_u4063  (
    .a({\u2_Display/n3384 ,\u2_Display/n3386 }),
    .b({\u2_Display/n3383 ,\u2_Display/n3385 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add105/c11 ),
    .f({\u2_Display/n3400 [13],\u2_Display/n3400 [11]}),
    .fco(\u2_Display/add105/c15 ),
    .fx({\u2_Display/n3400 [14],\u2_Display/n3400 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u15_al_u4064  (
    .a({\u2_Display/n3380 ,\u2_Display/n3382 }),
    .b({\u2_Display/n3379 ,\u2_Display/n3381 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add105/c15 ),
    .f({\u2_Display/n3400 [17],\u2_Display/n3400 [15]}),
    .fco(\u2_Display/add105/c19 ),
    .fx({\u2_Display/n3400 [18],\u2_Display/n3400 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u19_al_u4065  (
    .a({\u2_Display/n3376 ,\u2_Display/n3378 }),
    .b({\u2_Display/n3375 ,\u2_Display/n3377 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add105/c19 ),
    .f({\u2_Display/n3400 [21],\u2_Display/n3400 [19]}),
    .fco(\u2_Display/add105/c23 ),
    .fx({\u2_Display/n3400 [22],\u2_Display/n3400 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u23_al_u4066  (
    .a({\u2_Display/n3372 ,\u2_Display/n3374 }),
    .b({\u2_Display/n3371 ,\u2_Display/n3373 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add105/c23 ),
    .f({\u2_Display/n3400 [25],\u2_Display/n3400 [23]}),
    .fco(\u2_Display/add105/c27 ),
    .fx({\u2_Display/n3400 [26],\u2_Display/n3400 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u27_al_u4067  (
    .a({\u2_Display/n3368 ,\u2_Display/n3370 }),
    .b({\u2_Display/n3367 ,\u2_Display/n3369 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add105/c27 ),
    .f({\u2_Display/n3400 [29],\u2_Display/n3400 [27]}),
    .fco(\u2_Display/add105/c31 ),
    .fx({\u2_Display/n3400 [30],\u2_Display/n3400 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u31_al_u4068  (
    .a({open_n50568,\u2_Display/n3366 }),
    .c(2'b00),
    .d({open_n50573,1'b1}),
    .fci(\u2_Display/add105/c31 ),
    .f({open_n50590,\u2_Display/n3400 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u3_al_u4061  (
    .a({\u2_Display/n3392 ,\u2_Display/n3394 }),
    .b({\u2_Display/n3391 ,\u2_Display/n3393 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add105/c3 ),
    .f({\u2_Display/n3400 [5],\u2_Display/n3400 [3]}),
    .fco(\u2_Display/add105/c7 ),
    .fx({\u2_Display/n3400 [6],\u2_Display/n3400 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u7_al_u4062  (
    .a({\u2_Display/n3388 ,\u2_Display/n3390 }),
    .b({\u2_Display/n3387 ,\u2_Display/n3389 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add105/c7 ),
    .f({\u2_Display/n3400 [9],\u2_Display/n3400 [7]}),
    .fco(\u2_Display/add105/c11 ),
    .fx({\u2_Display/n3400 [10],\u2_Display/n3400 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/ucin_al_u4060  (
    .a({\u2_Display/n3396 ,1'b1}),
    .b({\u2_Display/n3395 ,\u2_Display/n3397 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3400 [1],open_n50649}),
    .fco(\u2_Display/add105/c3 ),
    .fx({\u2_Display/n3400 [2],\u2_Display/n3400 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add106/ucin_al_u5043"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add106/u3_al_u5044  (
    .a({\u2_Display/n3427 ,\u2_Display/n3429 }),
    .b({\u2_Display/n3426 ,\u2_Display/n3428 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b00),
    .fci(\u2_Display/add106/c3 ),
    .f({\u2_Display/n3435 [5],\u2_Display/n3435 [3]}),
    .fco(\u2_Display/add106/c7 ),
    .fx({\u2_Display/n3435 [6],\u2_Display/n3435 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add106/ucin_al_u5043"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add106/u7_al_u5045  (
    .a({\u2_Display/n3423 ,\u2_Display/n3425 }),
    .b({open_n50670,\u2_Display/n3424 }),
    .c(2'b00),
    .d(2'b01),
    .e({open_n50673,1'b1}),
    .fci(\u2_Display/add106/c7 ),
    .f({\u2_Display/n3435 [9],\u2_Display/n3435 [7]}),
    .fx({open_n50689,\u2_Display/n3435 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add106/ucin_al_u5043"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add106/ucin_al_u5043  (
    .a({\u2_Display/n3431 ,1'b1}),
    .b({\u2_Display/n3430 ,\u2_Display/n3432 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3435 [1],open_n50709}),
    .fco(\u2_Display/add106/c3 ),
    .fx({\u2_Display/n3435 [2],\u2_Display/n3435 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u11_al_u4072  (
    .a({\u2_Display/counta [13],\u2_Display/counta [11]}),
    .b({\u2_Display/counta [14],\u2_Display/counta [12]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add117/c11 ),
    .f({\u2_Display/n3788 [13],\u2_Display/n3788 [11]}),
    .fco(\u2_Display/add117/c15 ),
    .fx({\u2_Display/n3788 [14],\u2_Display/n3788 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u15_al_u4073  (
    .a({\u2_Display/counta [17],\u2_Display/counta [15]}),
    .b({\u2_Display/counta [18],\u2_Display/counta [16]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add117/c15 ),
    .f({\u2_Display/n3788 [17],\u2_Display/n3788 [15]}),
    .fco(\u2_Display/add117/c19 ),
    .fx({\u2_Display/n3788 [18],\u2_Display/n3788 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u19_al_u4074  (
    .a({\u2_Display/counta [21],\u2_Display/counta [19]}),
    .b({\u2_Display/counta [22],\u2_Display/counta [20]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add117/c19 ),
    .f({\u2_Display/n3788 [21],\u2_Display/n3788 [19]}),
    .fco(\u2_Display/add117/c23 ),
    .fx({\u2_Display/n3788 [22],\u2_Display/n3788 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u23_al_u4075  (
    .a({\u2_Display/counta [25],\u2_Display/counta [23]}),
    .b({\u2_Display/counta [26],\u2_Display/counta [24]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add117/c23 ),
    .f({\u2_Display/n3788 [25],\u2_Display/n3788 [23]}),
    .fco(\u2_Display/add117/c27 ),
    .fx({\u2_Display/n3788 [26],\u2_Display/n3788 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u27_al_u4076  (
    .a({\u2_Display/counta [29],\u2_Display/counta [27]}),
    .b({\u2_Display/counta [30],\u2_Display/counta [28]}),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add117/c27 ),
    .f({\u2_Display/n3788 [29],\u2_Display/n3788 [27]}),
    .fco(\u2_Display/add117/c31 ),
    .fx({\u2_Display/n3788 [30],\u2_Display/n3788 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u31_al_u4077  (
    .a({open_n50802,\u2_Display/counta [31]}),
    .c(2'b00),
    .d({open_n50807,1'b0}),
    .fci(\u2_Display/add117/c31 ),
    .f({open_n50824,\u2_Display/n3788 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u3_al_u4070  (
    .a({\u2_Display/counta [5],\u2_Display/counta [3]}),
    .b({\u2_Display/counta [6],\u2_Display/counta [4]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add117/c3 ),
    .f({\u2_Display/n3788 [5],\u2_Display/n3788 [3]}),
    .fco(\u2_Display/add117/c7 ),
    .fx({\u2_Display/n3788 [6],\u2_Display/n3788 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u7_al_u4071  (
    .a({\u2_Display/counta [9],\u2_Display/counta [7]}),
    .b({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add117/c7 ),
    .f({\u2_Display/n3788 [9],\u2_Display/n3788 [7]}),
    .fco(\u2_Display/add117/c11 ),
    .fx({\u2_Display/n3788 [10],\u2_Display/n3788 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/ucin_al_u4069  (
    .a({\u2_Display/counta [1],1'b1}),
    .b({\u2_Display/counta [2],\u2_Display/counta [0]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3788 [1],open_n50883}),
    .fco(\u2_Display/add117/c3 ),
    .fx({\u2_Display/n3788 [2],\u2_Display/n3788 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u11_al_u4081  (
    .a({\u2_Display/n3807 ,\u2_Display/n3809 }),
    .b({\u2_Display/n3806 ,\u2_Display/n3808 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add118/c11 ),
    .f({\u2_Display/n3823 [13],\u2_Display/n3823 [11]}),
    .fco(\u2_Display/add118/c15 ),
    .fx({\u2_Display/n3823 [14],\u2_Display/n3823 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u15_al_u4082  (
    .a({\u2_Display/n3803 ,\u2_Display/n3805 }),
    .b({\u2_Display/n3802 ,\u2_Display/n3804 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add118/c15 ),
    .f({\u2_Display/n3823 [17],\u2_Display/n3823 [15]}),
    .fco(\u2_Display/add118/c19 ),
    .fx({\u2_Display/n3823 [18],\u2_Display/n3823 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u19_al_u4083  (
    .a({\u2_Display/n3799 ,\u2_Display/n3801 }),
    .b({\u2_Display/n3798 ,\u2_Display/n3800 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add118/c19 ),
    .f({\u2_Display/n3823 [21],\u2_Display/n3823 [19]}),
    .fco(\u2_Display/add118/c23 ),
    .fx({\u2_Display/n3823 [22],\u2_Display/n3823 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u23_al_u4084  (
    .a({\u2_Display/n3795 ,\u2_Display/n3797 }),
    .b({\u2_Display/n3794 ,\u2_Display/n3796 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add118/c23 ),
    .f({\u2_Display/n3823 [25],\u2_Display/n3823 [23]}),
    .fco(\u2_Display/add118/c27 ),
    .fx({\u2_Display/n3823 [26],\u2_Display/n3823 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u27_al_u4085  (
    .a({\u2_Display/n3791 ,\u2_Display/n3793 }),
    .b({\u2_Display/n3790 ,\u2_Display/n3792 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add118/c27 ),
    .f({\u2_Display/n3823 [29],\u2_Display/n3823 [27]}),
    .fco(\u2_Display/add118/c31 ),
    .fx({\u2_Display/n3823 [30],\u2_Display/n3823 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u31_al_u4086  (
    .a({open_n50976,\u2_Display/n3789 }),
    .c(2'b00),
    .d({open_n50981,1'b1}),
    .fci(\u2_Display/add118/c31 ),
    .f({open_n50998,\u2_Display/n3823 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u3_al_u4079  (
    .a({\u2_Display/n3815 ,\u2_Display/n3817 }),
    .b({\u2_Display/n3814 ,\u2_Display/n3816 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add118/c3 ),
    .f({\u2_Display/n3823 [5],\u2_Display/n3823 [3]}),
    .fco(\u2_Display/add118/c7 ),
    .fx({\u2_Display/n3823 [6],\u2_Display/n3823 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u7_al_u4080  (
    .a({\u2_Display/n3811 ,\u2_Display/n3813 }),
    .b({\u2_Display/n3810 ,\u2_Display/n3812 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add118/c7 ),
    .f({\u2_Display/n3823 [9],\u2_Display/n3823 [7]}),
    .fco(\u2_Display/add118/c11 ),
    .fx({\u2_Display/n3823 [10],\u2_Display/n3823 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/ucin_al_u4078  (
    .a({\u2_Display/n3819 ,1'b1}),
    .b({\u2_Display/n3818 ,\u2_Display/n3820 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3823 [1],open_n51057}),
    .fco(\u2_Display/add118/c3 ),
    .fx({\u2_Display/n3823 [2],\u2_Display/n3823 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u11_al_u4090  (
    .a({\u2_Display/n3842 ,\u2_Display/n3844 }),
    .b({\u2_Display/n3841 ,\u2_Display/n3843 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add119/c11 ),
    .f({\u2_Display/n3858 [13],\u2_Display/n3858 [11]}),
    .fco(\u2_Display/add119/c15 ),
    .fx({\u2_Display/n3858 [14],\u2_Display/n3858 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u15_al_u4091  (
    .a({\u2_Display/n3838 ,\u2_Display/n3840 }),
    .b({\u2_Display/n3837 ,\u2_Display/n3839 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add119/c15 ),
    .f({\u2_Display/n3858 [17],\u2_Display/n3858 [15]}),
    .fco(\u2_Display/add119/c19 ),
    .fx({\u2_Display/n3858 [18],\u2_Display/n3858 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u19_al_u4092  (
    .a({\u2_Display/n3834 ,\u2_Display/n3836 }),
    .b({\u2_Display/n3833 ,\u2_Display/n3835 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add119/c19 ),
    .f({\u2_Display/n3858 [21],\u2_Display/n3858 [19]}),
    .fco(\u2_Display/add119/c23 ),
    .fx({\u2_Display/n3858 [22],\u2_Display/n3858 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u23_al_u4093  (
    .a({\u2_Display/n3830 ,\u2_Display/n3832 }),
    .b({\u2_Display/n3829 ,\u2_Display/n3831 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add119/c23 ),
    .f({\u2_Display/n3858 [25],\u2_Display/n3858 [23]}),
    .fco(\u2_Display/add119/c27 ),
    .fx({\u2_Display/n3858 [26],\u2_Display/n3858 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u27_al_u4094  (
    .a({\u2_Display/n3826 ,\u2_Display/n3828 }),
    .b({\u2_Display/n3825 ,\u2_Display/n3827 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add119/c27 ),
    .f({\u2_Display/n3858 [29],\u2_Display/n3858 [27]}),
    .fco(\u2_Display/add119/c31 ),
    .fx({\u2_Display/n3858 [30],\u2_Display/n3858 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u31_al_u4095  (
    .a({open_n51150,\u2_Display/n3824 }),
    .c(2'b00),
    .d({open_n51155,1'b1}),
    .fci(\u2_Display/add119/c31 ),
    .f({open_n51172,\u2_Display/n3858 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u3_al_u4088  (
    .a({\u2_Display/n3850 ,\u2_Display/n3852 }),
    .b({\u2_Display/n3849 ,\u2_Display/n3851 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add119/c3 ),
    .f({\u2_Display/n3858 [5],\u2_Display/n3858 [3]}),
    .fco(\u2_Display/add119/c7 ),
    .fx({\u2_Display/n3858 [6],\u2_Display/n3858 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u7_al_u4089  (
    .a({\u2_Display/n3846 ,\u2_Display/n3848 }),
    .b({\u2_Display/n3845 ,\u2_Display/n3847 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add119/c7 ),
    .f({\u2_Display/n3858 [9],\u2_Display/n3858 [7]}),
    .fco(\u2_Display/add119/c11 ),
    .fx({\u2_Display/n3858 [10],\u2_Display/n3858 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/ucin_al_u4087  (
    .a({\u2_Display/n3854 ,1'b1}),
    .b({\u2_Display/n3853 ,\u2_Display/n3855 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3858 [1],open_n51231}),
    .fco(\u2_Display/add119/c3 ),
    .fx({\u2_Display/n3858 [2],\u2_Display/n3858 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u11_al_u4099  (
    .a({\u2_Display/n3877 ,\u2_Display/n3879 }),
    .b({\u2_Display/n3876 ,\u2_Display/n3878 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add120/c11 ),
    .f({\u2_Display/n3893 [13],\u2_Display/n3893 [11]}),
    .fco(\u2_Display/add120/c15 ),
    .fx({\u2_Display/n3893 [14],\u2_Display/n3893 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u15_al_u4100  (
    .a({\u2_Display/n3873 ,\u2_Display/n3875 }),
    .b({\u2_Display/n3872 ,\u2_Display/n3874 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add120/c15 ),
    .f({\u2_Display/n3893 [17],\u2_Display/n3893 [15]}),
    .fco(\u2_Display/add120/c19 ),
    .fx({\u2_Display/n3893 [18],\u2_Display/n3893 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u19_al_u4101  (
    .a({\u2_Display/n3869 ,\u2_Display/n3871 }),
    .b({\u2_Display/n3868 ,\u2_Display/n3870 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add120/c19 ),
    .f({\u2_Display/n3893 [21],\u2_Display/n3893 [19]}),
    .fco(\u2_Display/add120/c23 ),
    .fx({\u2_Display/n3893 [22],\u2_Display/n3893 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u23_al_u4102  (
    .a({\u2_Display/n3865 ,\u2_Display/n3867 }),
    .b({\u2_Display/n3864 ,\u2_Display/n3866 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add120/c23 ),
    .f({\u2_Display/n3893 [25],\u2_Display/n3893 [23]}),
    .fco(\u2_Display/add120/c27 ),
    .fx({\u2_Display/n3893 [26],\u2_Display/n3893 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u27_al_u4103  (
    .a({\u2_Display/n3861 ,\u2_Display/n3863 }),
    .b({\u2_Display/n3860 ,\u2_Display/n3862 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add120/c27 ),
    .f({\u2_Display/n3893 [29],\u2_Display/n3893 [27]}),
    .fco(\u2_Display/add120/c31 ),
    .fx({\u2_Display/n3893 [30],\u2_Display/n3893 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u31_al_u4104  (
    .a({open_n51324,\u2_Display/n3859 }),
    .c(2'b00),
    .d({open_n51329,1'b1}),
    .fci(\u2_Display/add120/c31 ),
    .f({open_n51346,\u2_Display/n3893 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u3_al_u4097  (
    .a({\u2_Display/n3885 ,\u2_Display/n3887 }),
    .b({\u2_Display/n3884 ,\u2_Display/n3886 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add120/c3 ),
    .f({\u2_Display/n3893 [5],\u2_Display/n3893 [3]}),
    .fco(\u2_Display/add120/c7 ),
    .fx({\u2_Display/n3893 [6],\u2_Display/n3893 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u7_al_u4098  (
    .a({\u2_Display/n3881 ,\u2_Display/n3883 }),
    .b({\u2_Display/n3880 ,\u2_Display/n3882 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add120/c7 ),
    .f({\u2_Display/n3893 [9],\u2_Display/n3893 [7]}),
    .fco(\u2_Display/add120/c11 ),
    .fx({\u2_Display/n3893 [10],\u2_Display/n3893 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/ucin_al_u4096  (
    .a({\u2_Display/n3889 ,1'b1}),
    .b({\u2_Display/n3888 ,\u2_Display/n3890 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3893 [1],open_n51405}),
    .fco(\u2_Display/add120/c3 ),
    .fx({\u2_Display/n3893 [2],\u2_Display/n3893 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u11_al_u4108  (
    .a({\u2_Display/n3912 ,\u2_Display/n3914 }),
    .b({\u2_Display/n3911 ,\u2_Display/n3913 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add121/c11 ),
    .f({\u2_Display/n3928 [13],\u2_Display/n3928 [11]}),
    .fco(\u2_Display/add121/c15 ),
    .fx({\u2_Display/n3928 [14],\u2_Display/n3928 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u15_al_u4109  (
    .a({\u2_Display/n3908 ,\u2_Display/n3910 }),
    .b({\u2_Display/n3907 ,\u2_Display/n3909 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add121/c15 ),
    .f({\u2_Display/n3928 [17],\u2_Display/n3928 [15]}),
    .fco(\u2_Display/add121/c19 ),
    .fx({\u2_Display/n3928 [18],\u2_Display/n3928 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u19_al_u4110  (
    .a({\u2_Display/n3904 ,\u2_Display/n3906 }),
    .b({\u2_Display/n3903 ,\u2_Display/n3905 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add121/c19 ),
    .f({\u2_Display/n3928 [21],\u2_Display/n3928 [19]}),
    .fco(\u2_Display/add121/c23 ),
    .fx({\u2_Display/n3928 [22],\u2_Display/n3928 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u23_al_u4111  (
    .a({\u2_Display/n3900 ,\u2_Display/n3902 }),
    .b({\u2_Display/n3899 ,\u2_Display/n3901 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add121/c23 ),
    .f({\u2_Display/n3928 [25],\u2_Display/n3928 [23]}),
    .fco(\u2_Display/add121/c27 ),
    .fx({\u2_Display/n3928 [26],\u2_Display/n3928 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u27_al_u4112  (
    .a({\u2_Display/n3896 ,\u2_Display/n3898 }),
    .b({\u2_Display/n3895 ,\u2_Display/n3897 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add121/c27 ),
    .f({\u2_Display/n3928 [29],\u2_Display/n3928 [27]}),
    .fco(\u2_Display/add121/c31 ),
    .fx({\u2_Display/n3928 [30],\u2_Display/n3928 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u31_al_u4113  (
    .a({open_n51498,\u2_Display/n3894 }),
    .c(2'b00),
    .d({open_n51503,1'b1}),
    .fci(\u2_Display/add121/c31 ),
    .f({open_n51520,\u2_Display/n3928 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u3_al_u4106  (
    .a({\u2_Display/n3920 ,\u2_Display/n3922 }),
    .b({\u2_Display/n3919 ,\u2_Display/n3921 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add121/c3 ),
    .f({\u2_Display/n3928 [5],\u2_Display/n3928 [3]}),
    .fco(\u2_Display/add121/c7 ),
    .fx({\u2_Display/n3928 [6],\u2_Display/n3928 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u7_al_u4107  (
    .a({\u2_Display/n3916 ,\u2_Display/n3918 }),
    .b({\u2_Display/n3915 ,\u2_Display/n3917 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add121/c7 ),
    .f({\u2_Display/n3928 [9],\u2_Display/n3928 [7]}),
    .fco(\u2_Display/add121/c11 ),
    .fx({\u2_Display/n3928 [10],\u2_Display/n3928 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/ucin_al_u4105  (
    .a({\u2_Display/n3924 ,1'b1}),
    .b({\u2_Display/n3923 ,\u2_Display/n3925 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3928 [1],open_n51579}),
    .fco(\u2_Display/add121/c3 ),
    .fx({\u2_Display/n3928 [2],\u2_Display/n3928 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u11_al_u4117  (
    .a({\u2_Display/n3947 ,\u2_Display/n3949 }),
    .b({\u2_Display/n3946 ,\u2_Display/n3948 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add122/c11 ),
    .f({\u2_Display/n3963 [13],\u2_Display/n3963 [11]}),
    .fco(\u2_Display/add122/c15 ),
    .fx({\u2_Display/n3963 [14],\u2_Display/n3963 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u15_al_u4118  (
    .a({\u2_Display/n3943 ,\u2_Display/n3945 }),
    .b({\u2_Display/n3942 ,\u2_Display/n3944 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add122/c15 ),
    .f({\u2_Display/n3963 [17],\u2_Display/n3963 [15]}),
    .fco(\u2_Display/add122/c19 ),
    .fx({\u2_Display/n3963 [18],\u2_Display/n3963 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u19_al_u4119  (
    .a({\u2_Display/n3939 ,\u2_Display/n3941 }),
    .b({\u2_Display/n3938 ,\u2_Display/n3940 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add122/c19 ),
    .f({\u2_Display/n3963 [21],\u2_Display/n3963 [19]}),
    .fco(\u2_Display/add122/c23 ),
    .fx({\u2_Display/n3963 [22],\u2_Display/n3963 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u23_al_u4120  (
    .a({\u2_Display/n3935 ,\u2_Display/n3937 }),
    .b({\u2_Display/n3934 ,\u2_Display/n3936 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add122/c23 ),
    .f({\u2_Display/n3963 [25],\u2_Display/n3963 [23]}),
    .fco(\u2_Display/add122/c27 ),
    .fx({\u2_Display/n3963 [26],\u2_Display/n3963 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u27_al_u4121  (
    .a({\u2_Display/n3931 ,\u2_Display/n3933 }),
    .b({\u2_Display/n3930 ,\u2_Display/n3932 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add122/c27 ),
    .f({\u2_Display/n3963 [29],\u2_Display/n3963 [27]}),
    .fco(\u2_Display/add122/c31 ),
    .fx({\u2_Display/n3963 [30],\u2_Display/n3963 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u31_al_u4122  (
    .a({open_n51672,\u2_Display/n3929 }),
    .c(2'b00),
    .d({open_n51677,1'b1}),
    .fci(\u2_Display/add122/c31 ),
    .f({open_n51694,\u2_Display/n3963 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u3_al_u4115  (
    .a({\u2_Display/n3955 ,\u2_Display/n3957 }),
    .b({\u2_Display/n3954 ,\u2_Display/n3956 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add122/c3 ),
    .f({\u2_Display/n3963 [5],\u2_Display/n3963 [3]}),
    .fco(\u2_Display/add122/c7 ),
    .fx({\u2_Display/n3963 [6],\u2_Display/n3963 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u7_al_u4116  (
    .a({\u2_Display/n3951 ,\u2_Display/n3953 }),
    .b({\u2_Display/n3950 ,\u2_Display/n3952 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add122/c7 ),
    .f({\u2_Display/n3963 [9],\u2_Display/n3963 [7]}),
    .fco(\u2_Display/add122/c11 ),
    .fx({\u2_Display/n3963 [10],\u2_Display/n3963 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/ucin_al_u4114  (
    .a({\u2_Display/n3959 ,1'b1}),
    .b({\u2_Display/n3958 ,\u2_Display/n3960 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3963 [1],open_n51753}),
    .fco(\u2_Display/add122/c3 ),
    .fx({\u2_Display/n3963 [2],\u2_Display/n3963 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u11_al_u4126  (
    .a({\u2_Display/n3982 ,\u2_Display/n3984 }),
    .b({\u2_Display/n3981 ,\u2_Display/n3983 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add123/c11 ),
    .f({\u2_Display/n3998 [13],\u2_Display/n3998 [11]}),
    .fco(\u2_Display/add123/c15 ),
    .fx({\u2_Display/n3998 [14],\u2_Display/n3998 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u15_al_u4127  (
    .a({\u2_Display/n3978 ,\u2_Display/n3980 }),
    .b({\u2_Display/n3977 ,\u2_Display/n3979 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add123/c15 ),
    .f({\u2_Display/n3998 [17],\u2_Display/n3998 [15]}),
    .fco(\u2_Display/add123/c19 ),
    .fx({\u2_Display/n3998 [18],\u2_Display/n3998 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u19_al_u4128  (
    .a({\u2_Display/n3974 ,\u2_Display/n3976 }),
    .b({\u2_Display/n3973 ,\u2_Display/n3975 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add123/c19 ),
    .f({\u2_Display/n3998 [21],\u2_Display/n3998 [19]}),
    .fco(\u2_Display/add123/c23 ),
    .fx({\u2_Display/n3998 [22],\u2_Display/n3998 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u23_al_u4129  (
    .a({\u2_Display/n3970 ,\u2_Display/n3972 }),
    .b({\u2_Display/n3969 ,\u2_Display/n3971 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add123/c23 ),
    .f({\u2_Display/n3998 [25],\u2_Display/n3998 [23]}),
    .fco(\u2_Display/add123/c27 ),
    .fx({\u2_Display/n3998 [26],\u2_Display/n3998 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u27_al_u4130  (
    .a({\u2_Display/n3966 ,\u2_Display/n3968 }),
    .b({\u2_Display/n3965 ,\u2_Display/n3967 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add123/c27 ),
    .f({\u2_Display/n3998 [29],\u2_Display/n3998 [27]}),
    .fco(\u2_Display/add123/c31 ),
    .fx({\u2_Display/n3998 [30],\u2_Display/n3998 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u31_al_u4131  (
    .a({open_n51846,\u2_Display/n3964 }),
    .c(2'b00),
    .d({open_n51851,1'b1}),
    .fci(\u2_Display/add123/c31 ),
    .f({open_n51868,\u2_Display/n3998 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u3_al_u4124  (
    .a({\u2_Display/n3990 ,\u2_Display/n3992 }),
    .b({\u2_Display/n3989 ,\u2_Display/n3991 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add123/c3 ),
    .f({\u2_Display/n3998 [5],\u2_Display/n3998 [3]}),
    .fco(\u2_Display/add123/c7 ),
    .fx({\u2_Display/n3998 [6],\u2_Display/n3998 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u7_al_u4125  (
    .a({\u2_Display/n3986 ,\u2_Display/n3988 }),
    .b({\u2_Display/n3985 ,\u2_Display/n3987 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add123/c7 ),
    .f({\u2_Display/n3998 [9],\u2_Display/n3998 [7]}),
    .fco(\u2_Display/add123/c11 ),
    .fx({\u2_Display/n3998 [10],\u2_Display/n3998 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/ucin_al_u4123  (
    .a({\u2_Display/n3994 ,1'b1}),
    .b({\u2_Display/n3993 ,\u2_Display/n3995 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3998 [1],open_n51927}),
    .fco(\u2_Display/add123/c3 ),
    .fx({\u2_Display/n3998 [2],\u2_Display/n3998 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u11_al_u4135  (
    .a({\u2_Display/n4017 ,\u2_Display/n4019 }),
    .b({\u2_Display/n4016 ,\u2_Display/n4018 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add124/c11 ),
    .f({\u2_Display/n4033 [13],\u2_Display/n4033 [11]}),
    .fco(\u2_Display/add124/c15 ),
    .fx({\u2_Display/n4033 [14],\u2_Display/n4033 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u15_al_u4136  (
    .a({\u2_Display/n4013 ,\u2_Display/n4015 }),
    .b({\u2_Display/n4012 ,\u2_Display/n4014 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add124/c15 ),
    .f({\u2_Display/n4033 [17],\u2_Display/n4033 [15]}),
    .fco(\u2_Display/add124/c19 ),
    .fx({\u2_Display/n4033 [18],\u2_Display/n4033 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u19_al_u4137  (
    .a({\u2_Display/n4009 ,\u2_Display/n4011 }),
    .b({\u2_Display/n4008 ,\u2_Display/n4010 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add124/c19 ),
    .f({\u2_Display/n4033 [21],\u2_Display/n4033 [19]}),
    .fco(\u2_Display/add124/c23 ),
    .fx({\u2_Display/n4033 [22],\u2_Display/n4033 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u23_al_u4138  (
    .a({\u2_Display/n4005 ,\u2_Display/n4007 }),
    .b({\u2_Display/n4004 ,\u2_Display/n4006 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add124/c23 ),
    .f({\u2_Display/n4033 [25],\u2_Display/n4033 [23]}),
    .fco(\u2_Display/add124/c27 ),
    .fx({\u2_Display/n4033 [26],\u2_Display/n4033 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u27_al_u4139  (
    .a({\u2_Display/n4001 ,\u2_Display/n4003 }),
    .b({\u2_Display/n4000 ,\u2_Display/n4002 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add124/c27 ),
    .f({\u2_Display/n4033 [29],\u2_Display/n4033 [27]}),
    .fco(\u2_Display/add124/c31 ),
    .fx({\u2_Display/n4033 [30],\u2_Display/n4033 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u31_al_u4140  (
    .a({open_n52020,\u2_Display/n3999 }),
    .c(2'b00),
    .d({open_n52025,1'b1}),
    .fci(\u2_Display/add124/c31 ),
    .f({open_n52042,\u2_Display/n4033 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u3_al_u4133  (
    .a({\u2_Display/n4025 ,\u2_Display/n4027 }),
    .b({\u2_Display/n4024 ,\u2_Display/n4026 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add124/c3 ),
    .f({\u2_Display/n4033 [5],\u2_Display/n4033 [3]}),
    .fco(\u2_Display/add124/c7 ),
    .fx({\u2_Display/n4033 [6],\u2_Display/n4033 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u7_al_u4134  (
    .a({\u2_Display/n4021 ,\u2_Display/n4023 }),
    .b({\u2_Display/n4020 ,\u2_Display/n4022 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add124/c7 ),
    .f({\u2_Display/n4033 [9],\u2_Display/n4033 [7]}),
    .fco(\u2_Display/add124/c11 ),
    .fx({\u2_Display/n4033 [10],\u2_Display/n4033 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/ucin_al_u4132  (
    .a({\u2_Display/n4029 ,1'b1}),
    .b({\u2_Display/n4028 ,\u2_Display/n4030 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4033 [1],open_n52101}),
    .fco(\u2_Display/add124/c3 ),
    .fx({\u2_Display/n4033 [2],\u2_Display/n4033 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u11_al_u4144  (
    .a({\u2_Display/n4052 ,\u2_Display/n4054 }),
    .b({\u2_Display/n4051 ,\u2_Display/n4053 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add125/c11 ),
    .f({\u2_Display/n4068 [13],\u2_Display/n4068 [11]}),
    .fco(\u2_Display/add125/c15 ),
    .fx({\u2_Display/n4068 [14],\u2_Display/n4068 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u15_al_u4145  (
    .a({\u2_Display/n4048 ,\u2_Display/n4050 }),
    .b({\u2_Display/n4047 ,\u2_Display/n4049 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add125/c15 ),
    .f({\u2_Display/n4068 [17],\u2_Display/n4068 [15]}),
    .fco(\u2_Display/add125/c19 ),
    .fx({\u2_Display/n4068 [18],\u2_Display/n4068 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u19_al_u4146  (
    .a({\u2_Display/n4044 ,\u2_Display/n4046 }),
    .b({\u2_Display/n4043 ,\u2_Display/n4045 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add125/c19 ),
    .f({\u2_Display/n4068 [21],\u2_Display/n4068 [19]}),
    .fco(\u2_Display/add125/c23 ),
    .fx({\u2_Display/n4068 [22],\u2_Display/n4068 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u23_al_u4147  (
    .a({\u2_Display/n4040 ,\u2_Display/n4042 }),
    .b({\u2_Display/n4039 ,\u2_Display/n4041 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add125/c23 ),
    .f({\u2_Display/n4068 [25],\u2_Display/n4068 [23]}),
    .fco(\u2_Display/add125/c27 ),
    .fx({\u2_Display/n4068 [26],\u2_Display/n4068 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u27_al_u4148  (
    .a({\u2_Display/n4036 ,\u2_Display/n4038 }),
    .b({\u2_Display/n4035 ,\u2_Display/n4037 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add125/c27 ),
    .f({\u2_Display/n4068 [29],\u2_Display/n4068 [27]}),
    .fco(\u2_Display/add125/c31 ),
    .fx({\u2_Display/n4068 [30],\u2_Display/n4068 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u31_al_u4149  (
    .a({open_n52194,\u2_Display/n4034 }),
    .c(2'b00),
    .d({open_n52199,1'b1}),
    .fci(\u2_Display/add125/c31 ),
    .f({open_n52216,\u2_Display/n4068 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u3_al_u4142  (
    .a({\u2_Display/n4060 ,\u2_Display/n4062 }),
    .b({\u2_Display/n4059 ,\u2_Display/n4061 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add125/c3 ),
    .f({\u2_Display/n4068 [5],\u2_Display/n4068 [3]}),
    .fco(\u2_Display/add125/c7 ),
    .fx({\u2_Display/n4068 [6],\u2_Display/n4068 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u7_al_u4143  (
    .a({\u2_Display/n4056 ,\u2_Display/n4058 }),
    .b({\u2_Display/n4055 ,\u2_Display/n4057 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add125/c7 ),
    .f({\u2_Display/n4068 [9],\u2_Display/n4068 [7]}),
    .fco(\u2_Display/add125/c11 ),
    .fx({\u2_Display/n4068 [10],\u2_Display/n4068 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/ucin_al_u4141  (
    .a({\u2_Display/n4064 ,1'b1}),
    .b({\u2_Display/n4063 ,\u2_Display/n4065 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4068 [1],open_n52275}),
    .fco(\u2_Display/add125/c3 ),
    .fx({\u2_Display/n4068 [2],\u2_Display/n4068 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u11_al_u4153  (
    .a({\u2_Display/n4087 ,\u2_Display/n4089 }),
    .b({\u2_Display/n4086 ,\u2_Display/n4088 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add126/c11 ),
    .f({\u2_Display/n4103 [13],\u2_Display/n4103 [11]}),
    .fco(\u2_Display/add126/c15 ),
    .fx({\u2_Display/n4103 [14],\u2_Display/n4103 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u15_al_u4154  (
    .a({\u2_Display/n4083 ,\u2_Display/n4085 }),
    .b({\u2_Display/n4082 ,\u2_Display/n4084 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add126/c15 ),
    .f({\u2_Display/n4103 [17],\u2_Display/n4103 [15]}),
    .fco(\u2_Display/add126/c19 ),
    .fx({\u2_Display/n4103 [18],\u2_Display/n4103 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u19_al_u4155  (
    .a({\u2_Display/n4079 ,\u2_Display/n4081 }),
    .b({\u2_Display/n4078 ,\u2_Display/n4080 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add126/c19 ),
    .f({\u2_Display/n4103 [21],\u2_Display/n4103 [19]}),
    .fco(\u2_Display/add126/c23 ),
    .fx({\u2_Display/n4103 [22],\u2_Display/n4103 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u23_al_u4156  (
    .a({\u2_Display/n4075 ,\u2_Display/n4077 }),
    .b({\u2_Display/n4074 ,\u2_Display/n4076 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add126/c23 ),
    .f({\u2_Display/n4103 [25],\u2_Display/n4103 [23]}),
    .fco(\u2_Display/add126/c27 ),
    .fx({\u2_Display/n4103 [26],\u2_Display/n4103 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u27_al_u4157  (
    .a({\u2_Display/n4071 ,\u2_Display/n4073 }),
    .b({\u2_Display/n4070 ,\u2_Display/n4072 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add126/c27 ),
    .f({\u2_Display/n4103 [29],\u2_Display/n4103 [27]}),
    .fco(\u2_Display/add126/c31 ),
    .fx({\u2_Display/n4103 [30],\u2_Display/n4103 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u31_al_u4158  (
    .a({open_n52368,\u2_Display/n4069 }),
    .c(2'b00),
    .d({open_n52373,1'b1}),
    .fci(\u2_Display/add126/c31 ),
    .f({open_n52390,\u2_Display/n4103 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u3_al_u4151  (
    .a({\u2_Display/n4095 ,\u2_Display/n4097 }),
    .b({\u2_Display/n4094 ,\u2_Display/n4096 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add126/c3 ),
    .f({\u2_Display/n4103 [5],\u2_Display/n4103 [3]}),
    .fco(\u2_Display/add126/c7 ),
    .fx({\u2_Display/n4103 [6],\u2_Display/n4103 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u7_al_u4152  (
    .a({\u2_Display/n4091 ,\u2_Display/n4093 }),
    .b({\u2_Display/n4090 ,\u2_Display/n4092 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add126/c7 ),
    .f({\u2_Display/n4103 [9],\u2_Display/n4103 [7]}),
    .fco(\u2_Display/add126/c11 ),
    .fx({\u2_Display/n4103 [10],\u2_Display/n4103 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/ucin_al_u4150  (
    .a({\u2_Display/n4099 ,1'b1}),
    .b({\u2_Display/n4098 ,\u2_Display/n4100 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4103 [1],open_n52449}),
    .fco(\u2_Display/add126/c3 ),
    .fx({\u2_Display/n4103 [2],\u2_Display/n4103 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u11_al_u4162  (
    .a({\u2_Display/n4122 ,\u2_Display/n4124 }),
    .b({\u2_Display/n4121 ,\u2_Display/n4123 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add127/c11 ),
    .f({\u2_Display/n4138 [13],\u2_Display/n4138 [11]}),
    .fco(\u2_Display/add127/c15 ),
    .fx({\u2_Display/n4138 [14],\u2_Display/n4138 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u15_al_u4163  (
    .a({\u2_Display/n4118 ,\u2_Display/n4120 }),
    .b({\u2_Display/n4117 ,\u2_Display/n4119 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add127/c15 ),
    .f({\u2_Display/n4138 [17],\u2_Display/n4138 [15]}),
    .fco(\u2_Display/add127/c19 ),
    .fx({\u2_Display/n4138 [18],\u2_Display/n4138 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u19_al_u4164  (
    .a({\u2_Display/n4114 ,\u2_Display/n4116 }),
    .b({\u2_Display/n4113 ,\u2_Display/n4115 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add127/c19 ),
    .f({\u2_Display/n4138 [21],\u2_Display/n4138 [19]}),
    .fco(\u2_Display/add127/c23 ),
    .fx({\u2_Display/n4138 [22],\u2_Display/n4138 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u23_al_u4165  (
    .a({\u2_Display/n4110 ,\u2_Display/n4112 }),
    .b({\u2_Display/n4109 ,\u2_Display/n4111 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add127/c23 ),
    .f({\u2_Display/n4138 [25],\u2_Display/n4138 [23]}),
    .fco(\u2_Display/add127/c27 ),
    .fx({\u2_Display/n4138 [26],\u2_Display/n4138 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u27_al_u4166  (
    .a({\u2_Display/n4106 ,\u2_Display/n4108 }),
    .b({\u2_Display/n4105 ,\u2_Display/n4107 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add127/c27 ),
    .f({\u2_Display/n4138 [29],\u2_Display/n4138 [27]}),
    .fco(\u2_Display/add127/c31 ),
    .fx({\u2_Display/n4138 [30],\u2_Display/n4138 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u31_al_u4167  (
    .a({open_n52542,\u2_Display/n4104 }),
    .c(2'b00),
    .d({open_n52547,1'b1}),
    .fci(\u2_Display/add127/c31 ),
    .f({open_n52564,\u2_Display/n4138 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u3_al_u4160  (
    .a({\u2_Display/n4130 ,\u2_Display/n4132 }),
    .b({\u2_Display/n4129 ,\u2_Display/n4131 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add127/c3 ),
    .f({\u2_Display/n4138 [5],\u2_Display/n4138 [3]}),
    .fco(\u2_Display/add127/c7 ),
    .fx({\u2_Display/n4138 [6],\u2_Display/n4138 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u7_al_u4161  (
    .a({\u2_Display/n4126 ,\u2_Display/n4128 }),
    .b({\u2_Display/n4125 ,\u2_Display/n4127 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add127/c7 ),
    .f({\u2_Display/n4138 [9],\u2_Display/n4138 [7]}),
    .fco(\u2_Display/add127/c11 ),
    .fx({\u2_Display/n4138 [10],\u2_Display/n4138 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/ucin_al_u4159  (
    .a({\u2_Display/n4134 ,1'b1}),
    .b({\u2_Display/n4133 ,\u2_Display/n4135 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4138 [1],open_n52623}),
    .fco(\u2_Display/add127/c3 ),
    .fx({\u2_Display/n4138 [2],\u2_Display/n4138 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u11_al_u4171  (
    .a({\u2_Display/n4157 ,\u2_Display/n4159 }),
    .b({\u2_Display/n4156 ,\u2_Display/n4158 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add128/c11 ),
    .f({\u2_Display/n4173 [13],\u2_Display/n4173 [11]}),
    .fco(\u2_Display/add128/c15 ),
    .fx({\u2_Display/n4173 [14],\u2_Display/n4173 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u15_al_u4172  (
    .a({\u2_Display/n4153 ,\u2_Display/n4155 }),
    .b({\u2_Display/n4152 ,\u2_Display/n4154 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add128/c15 ),
    .f({\u2_Display/n4173 [17],\u2_Display/n4173 [15]}),
    .fco(\u2_Display/add128/c19 ),
    .fx({\u2_Display/n4173 [18],\u2_Display/n4173 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u19_al_u4173  (
    .a({\u2_Display/n4149 ,\u2_Display/n4151 }),
    .b({\u2_Display/n4148 ,\u2_Display/n4150 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add128/c19 ),
    .f({\u2_Display/n4173 [21],\u2_Display/n4173 [19]}),
    .fco(\u2_Display/add128/c23 ),
    .fx({\u2_Display/n4173 [22],\u2_Display/n4173 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u23_al_u4174  (
    .a({\u2_Display/n4145 ,\u2_Display/n4147 }),
    .b({\u2_Display/n4144 ,\u2_Display/n4146 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add128/c23 ),
    .f({\u2_Display/n4173 [25],\u2_Display/n4173 [23]}),
    .fco(\u2_Display/add128/c27 ),
    .fx({\u2_Display/n4173 [26],\u2_Display/n4173 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u27_al_u4175  (
    .a({\u2_Display/n4141 ,\u2_Display/n4143 }),
    .b({\u2_Display/n4140 ,\u2_Display/n4142 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add128/c27 ),
    .f({\u2_Display/n4173 [29],\u2_Display/n4173 [27]}),
    .fco(\u2_Display/add128/c31 ),
    .fx({\u2_Display/n4173 [30],\u2_Display/n4173 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u31_al_u4176  (
    .a({open_n52716,\u2_Display/n4139 }),
    .c(2'b00),
    .d({open_n52721,1'b1}),
    .fci(\u2_Display/add128/c31 ),
    .f({open_n52738,\u2_Display/n4173 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u3_al_u4169  (
    .a({\u2_Display/n4165 ,\u2_Display/n4167 }),
    .b({\u2_Display/n4164 ,\u2_Display/n4166 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add128/c3 ),
    .f({\u2_Display/n4173 [5],\u2_Display/n4173 [3]}),
    .fco(\u2_Display/add128/c7 ),
    .fx({\u2_Display/n4173 [6],\u2_Display/n4173 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u7_al_u4170  (
    .a({\u2_Display/n4161 ,\u2_Display/n4163 }),
    .b({\u2_Display/n4160 ,\u2_Display/n4162 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add128/c7 ),
    .f({\u2_Display/n4173 [9],\u2_Display/n4173 [7]}),
    .fco(\u2_Display/add128/c11 ),
    .fx({\u2_Display/n4173 [10],\u2_Display/n4173 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/ucin_al_u4168  (
    .a({\u2_Display/n4169 ,1'b1}),
    .b({\u2_Display/n4168 ,\u2_Display/n4170 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4173 [1],open_n52797}),
    .fco(\u2_Display/add128/c3 ),
    .fx({\u2_Display/n4173 [2],\u2_Display/n4173 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u11_al_u4180  (
    .a({\u2_Display/n4192 ,\u2_Display/n4194 }),
    .b({\u2_Display/n4191 ,\u2_Display/n4193 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add129/c11 ),
    .f({\u2_Display/n4208 [13],\u2_Display/n4208 [11]}),
    .fco(\u2_Display/add129/c15 ),
    .fx({\u2_Display/n4208 [14],\u2_Display/n4208 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u15_al_u4181  (
    .a({\u2_Display/n4188 ,\u2_Display/n4190 }),
    .b({\u2_Display/n4187 ,\u2_Display/n4189 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add129/c15 ),
    .f({\u2_Display/n4208 [17],\u2_Display/n4208 [15]}),
    .fco(\u2_Display/add129/c19 ),
    .fx({\u2_Display/n4208 [18],\u2_Display/n4208 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u19_al_u4182  (
    .a({\u2_Display/n4184 ,\u2_Display/n4186 }),
    .b({\u2_Display/n4183 ,\u2_Display/n4185 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add129/c19 ),
    .f({\u2_Display/n4208 [21],\u2_Display/n4208 [19]}),
    .fco(\u2_Display/add129/c23 ),
    .fx({\u2_Display/n4208 [22],\u2_Display/n4208 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u23_al_u4183  (
    .a({\u2_Display/n4180 ,\u2_Display/n4182 }),
    .b({\u2_Display/n4179 ,\u2_Display/n4181 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add129/c23 ),
    .f({\u2_Display/n4208 [25],\u2_Display/n4208 [23]}),
    .fco(\u2_Display/add129/c27 ),
    .fx({\u2_Display/n4208 [26],\u2_Display/n4208 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u27_al_u4184  (
    .a({\u2_Display/n4176 ,\u2_Display/n4178 }),
    .b({\u2_Display/n4175 ,\u2_Display/n4177 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add129/c27 ),
    .f({\u2_Display/n4208 [29],\u2_Display/n4208 [27]}),
    .fco(\u2_Display/add129/c31 ),
    .fx({\u2_Display/n4208 [30],\u2_Display/n4208 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u31_al_u4185  (
    .a({open_n52890,\u2_Display/n4174 }),
    .c(2'b00),
    .d({open_n52895,1'b1}),
    .fci(\u2_Display/add129/c31 ),
    .f({open_n52912,\u2_Display/n4208 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u3_al_u4178  (
    .a({\u2_Display/n4200 ,\u2_Display/n4202 }),
    .b({\u2_Display/n4199 ,\u2_Display/n4201 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add129/c3 ),
    .f({\u2_Display/n4208 [5],\u2_Display/n4208 [3]}),
    .fco(\u2_Display/add129/c7 ),
    .fx({\u2_Display/n4208 [6],\u2_Display/n4208 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u7_al_u4179  (
    .a({\u2_Display/n4196 ,\u2_Display/n4198 }),
    .b({\u2_Display/n4195 ,\u2_Display/n4197 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add129/c7 ),
    .f({\u2_Display/n4208 [9],\u2_Display/n4208 [7]}),
    .fco(\u2_Display/add129/c11 ),
    .fx({\u2_Display/n4208 [10],\u2_Display/n4208 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/ucin_al_u4177  (
    .a({\u2_Display/n4204 ,1'b1}),
    .b({\u2_Display/n4203 ,\u2_Display/n4205 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4208 [1],open_n52971}),
    .fco(\u2_Display/add129/c3 ),
    .fx({\u2_Display/n4208 [2],\u2_Display/n4208 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u11_al_u4189  (
    .a({\u2_Display/n4227 ,\u2_Display/n4229 }),
    .b({\u2_Display/n4226 ,\u2_Display/n4228 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add130/c11 ),
    .f({\u2_Display/n4243 [13],\u2_Display/n4243 [11]}),
    .fco(\u2_Display/add130/c15 ),
    .fx({\u2_Display/n4243 [14],\u2_Display/n4243 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u15_al_u4190  (
    .a({\u2_Display/n4223 ,\u2_Display/n4225 }),
    .b({\u2_Display/n4222 ,\u2_Display/n4224 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add130/c15 ),
    .f({\u2_Display/n4243 [17],\u2_Display/n4243 [15]}),
    .fco(\u2_Display/add130/c19 ),
    .fx({\u2_Display/n4243 [18],\u2_Display/n4243 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u19_al_u4191  (
    .a({\u2_Display/n4219 ,\u2_Display/n4221 }),
    .b({\u2_Display/n4218 ,\u2_Display/n4220 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add130/c19 ),
    .f({\u2_Display/n4243 [21],\u2_Display/n4243 [19]}),
    .fco(\u2_Display/add130/c23 ),
    .fx({\u2_Display/n4243 [22],\u2_Display/n4243 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u23_al_u4192  (
    .a({\u2_Display/n4215 ,\u2_Display/n4217 }),
    .b({\u2_Display/n4214 ,\u2_Display/n4216 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add130/c23 ),
    .f({\u2_Display/n4243 [25],\u2_Display/n4243 [23]}),
    .fco(\u2_Display/add130/c27 ),
    .fx({\u2_Display/n4243 [26],\u2_Display/n4243 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u27_al_u4193  (
    .a({\u2_Display/n4211 ,\u2_Display/n4213 }),
    .b({\u2_Display/n4210 ,\u2_Display/n4212 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add130/c27 ),
    .f({\u2_Display/n4243 [29],\u2_Display/n4243 [27]}),
    .fco(\u2_Display/add130/c31 ),
    .fx({\u2_Display/n4243 [30],\u2_Display/n4243 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u31_al_u4194  (
    .a({open_n53064,\u2_Display/n4209 }),
    .c(2'b00),
    .d({open_n53069,1'b1}),
    .fci(\u2_Display/add130/c31 ),
    .f({open_n53086,\u2_Display/n4243 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u3_al_u4187  (
    .a({\u2_Display/n4235 ,\u2_Display/n4237 }),
    .b({\u2_Display/n4234 ,\u2_Display/n4236 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add130/c3 ),
    .f({\u2_Display/n4243 [5],\u2_Display/n4243 [3]}),
    .fco(\u2_Display/add130/c7 ),
    .fx({\u2_Display/n4243 [6],\u2_Display/n4243 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u7_al_u4188  (
    .a({\u2_Display/n4231 ,\u2_Display/n4233 }),
    .b({\u2_Display/n4230 ,\u2_Display/n4232 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add130/c7 ),
    .f({\u2_Display/n4243 [9],\u2_Display/n4243 [7]}),
    .fco(\u2_Display/add130/c11 ),
    .fx({\u2_Display/n4243 [10],\u2_Display/n4243 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/ucin_al_u4186  (
    .a({\u2_Display/n4239 ,1'b1}),
    .b({\u2_Display/n4238 ,\u2_Display/n4240 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4243 [1],open_n53145}),
    .fco(\u2_Display/add130/c3 ),
    .fx({\u2_Display/n4243 [2],\u2_Display/n4243 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u11_al_u4198  (
    .a({\u2_Display/n4262 ,\u2_Display/n4264 }),
    .b({\u2_Display/n4261 ,\u2_Display/n4263 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add131/c11 ),
    .f({\u2_Display/n4278 [13],\u2_Display/n4278 [11]}),
    .fco(\u2_Display/add131/c15 ),
    .fx({\u2_Display/n4278 [14],\u2_Display/n4278 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u15_al_u4199  (
    .a({\u2_Display/n4258 ,\u2_Display/n4260 }),
    .b({\u2_Display/n4257 ,\u2_Display/n4259 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add131/c15 ),
    .f({\u2_Display/n4278 [17],\u2_Display/n4278 [15]}),
    .fco(\u2_Display/add131/c19 ),
    .fx({\u2_Display/n4278 [18],\u2_Display/n4278 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u19_al_u4200  (
    .a({\u2_Display/n4254 ,\u2_Display/n4256 }),
    .b({\u2_Display/n4253 ,\u2_Display/n4255 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add131/c19 ),
    .f({\u2_Display/n4278 [21],\u2_Display/n4278 [19]}),
    .fco(\u2_Display/add131/c23 ),
    .fx({\u2_Display/n4278 [22],\u2_Display/n4278 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u23_al_u4201  (
    .a({\u2_Display/n4250 ,\u2_Display/n4252 }),
    .b({\u2_Display/n4249 ,\u2_Display/n4251 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add131/c23 ),
    .f({\u2_Display/n4278 [25],\u2_Display/n4278 [23]}),
    .fco(\u2_Display/add131/c27 ),
    .fx({\u2_Display/n4278 [26],\u2_Display/n4278 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u27_al_u4202  (
    .a({\u2_Display/n4246 ,\u2_Display/n4248 }),
    .b({\u2_Display/n4245 ,\u2_Display/n4247 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add131/c27 ),
    .f({\u2_Display/n4278 [29],\u2_Display/n4278 [27]}),
    .fco(\u2_Display/add131/c31 ),
    .fx({\u2_Display/n4278 [30],\u2_Display/n4278 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u31_al_u4203  (
    .a({open_n53238,\u2_Display/n4244 }),
    .c(2'b00),
    .d({open_n53243,1'b1}),
    .fci(\u2_Display/add131/c31 ),
    .f({open_n53260,\u2_Display/n4278 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u3_al_u4196  (
    .a({\u2_Display/n4270 ,\u2_Display/n4272 }),
    .b({\u2_Display/n4269 ,\u2_Display/n4271 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add131/c3 ),
    .f({\u2_Display/n4278 [5],\u2_Display/n4278 [3]}),
    .fco(\u2_Display/add131/c7 ),
    .fx({\u2_Display/n4278 [6],\u2_Display/n4278 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u7_al_u4197  (
    .a({\u2_Display/n4266 ,\u2_Display/n4268 }),
    .b({\u2_Display/n4265 ,\u2_Display/n4267 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add131/c7 ),
    .f({\u2_Display/n4278 [9],\u2_Display/n4278 [7]}),
    .fco(\u2_Display/add131/c11 ),
    .fx({\u2_Display/n4278 [10],\u2_Display/n4278 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/ucin_al_u4195  (
    .a({\u2_Display/n4274 ,1'b1}),
    .b({\u2_Display/n4273 ,\u2_Display/n4275 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4278 [1],open_n53319}),
    .fco(\u2_Display/add131/c3 ),
    .fx({\u2_Display/n4278 [2],\u2_Display/n4278 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u11_al_u4207  (
    .a({\u2_Display/n4297 ,\u2_Display/n4299 }),
    .b({\u2_Display/n4296 ,\u2_Display/n4298 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add132/c11 ),
    .f({\u2_Display/n4313 [13],\u2_Display/n4313 [11]}),
    .fco(\u2_Display/add132/c15 ),
    .fx({\u2_Display/n4313 [14],\u2_Display/n4313 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u15_al_u4208  (
    .a({\u2_Display/n4293 ,\u2_Display/n4295 }),
    .b({\u2_Display/n4292 ,\u2_Display/n4294 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add132/c15 ),
    .f({\u2_Display/n4313 [17],\u2_Display/n4313 [15]}),
    .fco(\u2_Display/add132/c19 ),
    .fx({\u2_Display/n4313 [18],\u2_Display/n4313 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u19_al_u4209  (
    .a({\u2_Display/n4289 ,\u2_Display/n4291 }),
    .b({\u2_Display/n4288 ,\u2_Display/n4290 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add132/c19 ),
    .f({\u2_Display/n4313 [21],\u2_Display/n4313 [19]}),
    .fco(\u2_Display/add132/c23 ),
    .fx({\u2_Display/n4313 [22],\u2_Display/n4313 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u23_al_u4210  (
    .a({\u2_Display/n4285 ,\u2_Display/n4287 }),
    .b({\u2_Display/n4284 ,\u2_Display/n4286 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add132/c23 ),
    .f({\u2_Display/n4313 [25],\u2_Display/n4313 [23]}),
    .fco(\u2_Display/add132/c27 ),
    .fx({\u2_Display/n4313 [26],\u2_Display/n4313 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u27_al_u4211  (
    .a({\u2_Display/n4281 ,\u2_Display/n4283 }),
    .b({\u2_Display/n4280 ,\u2_Display/n4282 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add132/c27 ),
    .f({\u2_Display/n4313 [29],\u2_Display/n4313 [27]}),
    .fco(\u2_Display/add132/c31 ),
    .fx({\u2_Display/n4313 [30],\u2_Display/n4313 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u31_al_u4212  (
    .a({open_n53412,\u2_Display/n4279 }),
    .c(2'b00),
    .d({open_n53417,1'b1}),
    .fci(\u2_Display/add132/c31 ),
    .f({open_n53434,\u2_Display/n4313 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u3_al_u4205  (
    .a({\u2_Display/n4305 ,\u2_Display/n4307 }),
    .b({\u2_Display/n4304 ,\u2_Display/n4306 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add132/c3 ),
    .f({\u2_Display/n4313 [5],\u2_Display/n4313 [3]}),
    .fco(\u2_Display/add132/c7 ),
    .fx({\u2_Display/n4313 [6],\u2_Display/n4313 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u7_al_u4206  (
    .a({\u2_Display/n4301 ,\u2_Display/n4303 }),
    .b({\u2_Display/n4300 ,\u2_Display/n4302 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add132/c7 ),
    .f({\u2_Display/n4313 [9],\u2_Display/n4313 [7]}),
    .fco(\u2_Display/add132/c11 ),
    .fx({\u2_Display/n4313 [10],\u2_Display/n4313 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/ucin_al_u4204  (
    .a({\u2_Display/n4309 ,1'b1}),
    .b({\u2_Display/n4308 ,\u2_Display/n4310 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4313 [1],open_n53493}),
    .fco(\u2_Display/add132/c3 ),
    .fx({\u2_Display/n4313 [2],\u2_Display/n4313 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u11_al_u4216  (
    .a({\u2_Display/n4332 ,\u2_Display/n4334 }),
    .b({\u2_Display/n4331 ,\u2_Display/n4333 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add133/c11 ),
    .f({\u2_Display/n4348 [13],\u2_Display/n4348 [11]}),
    .fco(\u2_Display/add133/c15 ),
    .fx({\u2_Display/n4348 [14],\u2_Display/n4348 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u15_al_u4217  (
    .a({\u2_Display/n4328 ,\u2_Display/n4330 }),
    .b({\u2_Display/n4327 ,\u2_Display/n4329 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add133/c15 ),
    .f({\u2_Display/n4348 [17],\u2_Display/n4348 [15]}),
    .fco(\u2_Display/add133/c19 ),
    .fx({\u2_Display/n4348 [18],\u2_Display/n4348 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u19_al_u4218  (
    .a({\u2_Display/n4324 ,\u2_Display/n4326 }),
    .b({\u2_Display/n4323 ,\u2_Display/n4325 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add133/c19 ),
    .f({\u2_Display/n4348 [21],\u2_Display/n4348 [19]}),
    .fco(\u2_Display/add133/c23 ),
    .fx({\u2_Display/n4348 [22],\u2_Display/n4348 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u23_al_u4219  (
    .a({\u2_Display/n4320 ,\u2_Display/n4322 }),
    .b({\u2_Display/n4319 ,\u2_Display/n4321 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add133/c23 ),
    .f({\u2_Display/n4348 [25],\u2_Display/n4348 [23]}),
    .fco(\u2_Display/add133/c27 ),
    .fx({\u2_Display/n4348 [26],\u2_Display/n4348 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u27_al_u4220  (
    .a({\u2_Display/n4316 ,\u2_Display/n4318 }),
    .b({\u2_Display/n4315 ,\u2_Display/n4317 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add133/c27 ),
    .f({\u2_Display/n4348 [29],\u2_Display/n4348 [27]}),
    .fco(\u2_Display/add133/c31 ),
    .fx({\u2_Display/n4348 [30],\u2_Display/n4348 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u31_al_u4221  (
    .a({open_n53586,\u2_Display/n4314 }),
    .c(2'b00),
    .d({open_n53591,1'b1}),
    .fci(\u2_Display/add133/c31 ),
    .f({open_n53608,\u2_Display/n4348 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u3_al_u4214  (
    .a({\u2_Display/n4340 ,\u2_Display/n4342 }),
    .b({\u2_Display/n4339 ,\u2_Display/n4341 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add133/c3 ),
    .f({\u2_Display/n4348 [5],\u2_Display/n4348 [3]}),
    .fco(\u2_Display/add133/c7 ),
    .fx({\u2_Display/n4348 [6],\u2_Display/n4348 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u7_al_u4215  (
    .a({\u2_Display/n4336 ,\u2_Display/n4338 }),
    .b({\u2_Display/n4335 ,\u2_Display/n4337 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add133/c7 ),
    .f({\u2_Display/n4348 [9],\u2_Display/n4348 [7]}),
    .fco(\u2_Display/add133/c11 ),
    .fx({\u2_Display/n4348 [10],\u2_Display/n4348 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/ucin_al_u4213  (
    .a({\u2_Display/n4344 ,1'b1}),
    .b({\u2_Display/n4343 ,\u2_Display/n4345 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4348 [1],open_n53667}),
    .fco(\u2_Display/add133/c3 ),
    .fx({\u2_Display/n4348 [2],\u2_Display/n4348 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u11_al_u4225  (
    .a({\u2_Display/n4367 ,\u2_Display/n4369 }),
    .b({\u2_Display/n4366 ,\u2_Display/n4368 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add134/c11 ),
    .f({\u2_Display/n4383 [13],\u2_Display/n4383 [11]}),
    .fco(\u2_Display/add134/c15 ),
    .fx({\u2_Display/n4383 [14],\u2_Display/n4383 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u15_al_u4226  (
    .a({\u2_Display/n4363 ,\u2_Display/n4365 }),
    .b({\u2_Display/n4362 ,\u2_Display/n4364 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add134/c15 ),
    .f({\u2_Display/n4383 [17],\u2_Display/n4383 [15]}),
    .fco(\u2_Display/add134/c19 ),
    .fx({\u2_Display/n4383 [18],\u2_Display/n4383 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u19_al_u4227  (
    .a({\u2_Display/n4359 ,\u2_Display/n4361 }),
    .b({\u2_Display/n4358 ,\u2_Display/n4360 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add134/c19 ),
    .f({\u2_Display/n4383 [21],\u2_Display/n4383 [19]}),
    .fco(\u2_Display/add134/c23 ),
    .fx({\u2_Display/n4383 [22],\u2_Display/n4383 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u23_al_u4228  (
    .a({\u2_Display/n4355 ,\u2_Display/n4357 }),
    .b({\u2_Display/n4354 ,\u2_Display/n4356 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add134/c23 ),
    .f({\u2_Display/n4383 [25],\u2_Display/n4383 [23]}),
    .fco(\u2_Display/add134/c27 ),
    .fx({\u2_Display/n4383 [26],\u2_Display/n4383 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u27_al_u4229  (
    .a({\u2_Display/n4351 ,\u2_Display/n4353 }),
    .b({\u2_Display/n4350 ,\u2_Display/n4352 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add134/c27 ),
    .f({\u2_Display/n4383 [29],\u2_Display/n4383 [27]}),
    .fco(\u2_Display/add134/c31 ),
    .fx({\u2_Display/n4383 [30],\u2_Display/n4383 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u31_al_u4230  (
    .a({open_n53760,\u2_Display/n4349 }),
    .c(2'b00),
    .d({open_n53765,1'b1}),
    .fci(\u2_Display/add134/c31 ),
    .f({open_n53782,\u2_Display/n4383 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u3_al_u4223  (
    .a({\u2_Display/n4375 ,\u2_Display/n4377 }),
    .b({\u2_Display/n4374 ,\u2_Display/n4376 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add134/c3 ),
    .f({\u2_Display/n4383 [5],\u2_Display/n4383 [3]}),
    .fco(\u2_Display/add134/c7 ),
    .fx({\u2_Display/n4383 [6],\u2_Display/n4383 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u7_al_u4224  (
    .a({\u2_Display/n4371 ,\u2_Display/n4373 }),
    .b({\u2_Display/n4370 ,\u2_Display/n4372 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add134/c7 ),
    .f({\u2_Display/n4383 [9],\u2_Display/n4383 [7]}),
    .fco(\u2_Display/add134/c11 ),
    .fx({\u2_Display/n4383 [10],\u2_Display/n4383 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/ucin_al_u4222  (
    .a({\u2_Display/n4379 ,1'b1}),
    .b({\u2_Display/n4378 ,\u2_Display/n4380 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4383 [1],open_n53841}),
    .fco(\u2_Display/add134/c3 ),
    .fx({\u2_Display/n4383 [2],\u2_Display/n4383 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u11_al_u4234  (
    .a({\u2_Display/n4402 ,\u2_Display/n4404 }),
    .b({\u2_Display/n4401 ,\u2_Display/n4403 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add135/c11 ),
    .f({\u2_Display/n4418 [13],\u2_Display/n4418 [11]}),
    .fco(\u2_Display/add135/c15 ),
    .fx({\u2_Display/n4418 [14],\u2_Display/n4418 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u15_al_u4235  (
    .a({\u2_Display/n4398 ,\u2_Display/n4400 }),
    .b({\u2_Display/n4397 ,\u2_Display/n4399 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add135/c15 ),
    .f({\u2_Display/n4418 [17],\u2_Display/n4418 [15]}),
    .fco(\u2_Display/add135/c19 ),
    .fx({\u2_Display/n4418 [18],\u2_Display/n4418 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u19_al_u4236  (
    .a({\u2_Display/n4394 ,\u2_Display/n4396 }),
    .b({\u2_Display/n4393 ,\u2_Display/n4395 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add135/c19 ),
    .f({\u2_Display/n4418 [21],\u2_Display/n4418 [19]}),
    .fco(\u2_Display/add135/c23 ),
    .fx({\u2_Display/n4418 [22],\u2_Display/n4418 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u23_al_u4237  (
    .a({\u2_Display/n4390 ,\u2_Display/n4392 }),
    .b({\u2_Display/n4389 ,\u2_Display/n4391 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add135/c23 ),
    .f({\u2_Display/n4418 [25],\u2_Display/n4418 [23]}),
    .fco(\u2_Display/add135/c27 ),
    .fx({\u2_Display/n4418 [26],\u2_Display/n4418 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u27_al_u4238  (
    .a({\u2_Display/n4386 ,\u2_Display/n4388 }),
    .b({\u2_Display/n4385 ,\u2_Display/n4387 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add135/c27 ),
    .f({\u2_Display/n4418 [29],\u2_Display/n4418 [27]}),
    .fco(\u2_Display/add135/c31 ),
    .fx({\u2_Display/n4418 [30],\u2_Display/n4418 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u31_al_u4239  (
    .a({open_n53934,\u2_Display/n4384 }),
    .c(2'b00),
    .d({open_n53939,1'b1}),
    .fci(\u2_Display/add135/c31 ),
    .f({open_n53956,\u2_Display/n4418 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u3_al_u4232  (
    .a({\u2_Display/n4410 ,\u2_Display/n4412 }),
    .b({\u2_Display/n4409 ,\u2_Display/n4411 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add135/c3 ),
    .f({\u2_Display/n4418 [5],\u2_Display/n4418 [3]}),
    .fco(\u2_Display/add135/c7 ),
    .fx({\u2_Display/n4418 [6],\u2_Display/n4418 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u7_al_u4233  (
    .a({\u2_Display/n4406 ,\u2_Display/n4408 }),
    .b({\u2_Display/n4405 ,\u2_Display/n4407 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add135/c7 ),
    .f({\u2_Display/n4418 [9],\u2_Display/n4418 [7]}),
    .fco(\u2_Display/add135/c11 ),
    .fx({\u2_Display/n4418 [10],\u2_Display/n4418 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/ucin_al_u4231  (
    .a({\u2_Display/n4414 ,1'b1}),
    .b({\u2_Display/n4413 ,\u2_Display/n4415 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4418 [1],open_n54015}),
    .fco(\u2_Display/add135/c3 ),
    .fx({\u2_Display/n4418 [2],\u2_Display/n4418 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u11_al_u4243  (
    .a({\u2_Display/n4437 ,\u2_Display/n4439 }),
    .b({\u2_Display/n4436 ,\u2_Display/n4438 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add136/c11 ),
    .f({\u2_Display/n4453 [13],\u2_Display/n4453 [11]}),
    .fco(\u2_Display/add136/c15 ),
    .fx({\u2_Display/n4453 [14],\u2_Display/n4453 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u15_al_u4244  (
    .a({\u2_Display/n4433 ,\u2_Display/n4435 }),
    .b({\u2_Display/n4432 ,\u2_Display/n4434 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add136/c15 ),
    .f({\u2_Display/n4453 [17],\u2_Display/n4453 [15]}),
    .fco(\u2_Display/add136/c19 ),
    .fx({\u2_Display/n4453 [18],\u2_Display/n4453 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u19_al_u4245  (
    .a({\u2_Display/n4429 ,\u2_Display/n4431 }),
    .b({\u2_Display/n4428 ,\u2_Display/n4430 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add136/c19 ),
    .f({\u2_Display/n4453 [21],\u2_Display/n4453 [19]}),
    .fco(\u2_Display/add136/c23 ),
    .fx({\u2_Display/n4453 [22],\u2_Display/n4453 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u23_al_u4246  (
    .a({\u2_Display/n4425 ,\u2_Display/n4427 }),
    .b({\u2_Display/n4424 ,\u2_Display/n4426 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add136/c23 ),
    .f({\u2_Display/n4453 [25],\u2_Display/n4453 [23]}),
    .fco(\u2_Display/add136/c27 ),
    .fx({\u2_Display/n4453 [26],\u2_Display/n4453 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u27_al_u4247  (
    .a({\u2_Display/n4421 ,\u2_Display/n4423 }),
    .b({\u2_Display/n4420 ,\u2_Display/n4422 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add136/c27 ),
    .f({\u2_Display/n4453 [29],\u2_Display/n4453 [27]}),
    .fco(\u2_Display/add136/c31 ),
    .fx({\u2_Display/n4453 [30],\u2_Display/n4453 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u31_al_u4248  (
    .a({open_n54108,\u2_Display/n4419 }),
    .c(2'b00),
    .d({open_n54113,1'b1}),
    .fci(\u2_Display/add136/c31 ),
    .f({open_n54130,\u2_Display/n4453 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u3_al_u4241  (
    .a({\u2_Display/n4445 ,\u2_Display/n4447 }),
    .b({\u2_Display/n4444 ,\u2_Display/n4446 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add136/c3 ),
    .f({\u2_Display/n4453 [5],\u2_Display/n4453 [3]}),
    .fco(\u2_Display/add136/c7 ),
    .fx({\u2_Display/n4453 [6],\u2_Display/n4453 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u7_al_u4242  (
    .a({\u2_Display/n4441 ,\u2_Display/n4443 }),
    .b({\u2_Display/n4440 ,\u2_Display/n4442 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add136/c7 ),
    .f({\u2_Display/n4453 [9],\u2_Display/n4453 [7]}),
    .fco(\u2_Display/add136/c11 ),
    .fx({\u2_Display/n4453 [10],\u2_Display/n4453 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/ucin_al_u4240  (
    .a({\u2_Display/n4449 ,1'b1}),
    .b({\u2_Display/n4448 ,\u2_Display/n4450 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4453 [1],open_n54189}),
    .fco(\u2_Display/add136/c3 ),
    .fx({\u2_Display/n4453 [2],\u2_Display/n4453 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u11_al_u4252  (
    .a({\u2_Display/n4472 ,\u2_Display/n4474 }),
    .b({\u2_Display/n4471 ,\u2_Display/n4473 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add137/c11 ),
    .f({\u2_Display/n4488 [13],\u2_Display/n4488 [11]}),
    .fco(\u2_Display/add137/c15 ),
    .fx({\u2_Display/n4488 [14],\u2_Display/n4488 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u15_al_u4253  (
    .a({\u2_Display/n4468 ,\u2_Display/n4470 }),
    .b({\u2_Display/n4467 ,\u2_Display/n4469 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add137/c15 ),
    .f({\u2_Display/n4488 [17],\u2_Display/n4488 [15]}),
    .fco(\u2_Display/add137/c19 ),
    .fx({\u2_Display/n4488 [18],\u2_Display/n4488 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u19_al_u4254  (
    .a({\u2_Display/n4464 ,\u2_Display/n4466 }),
    .b({\u2_Display/n4463 ,\u2_Display/n4465 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add137/c19 ),
    .f({\u2_Display/n4488 [21],\u2_Display/n4488 [19]}),
    .fco(\u2_Display/add137/c23 ),
    .fx({\u2_Display/n4488 [22],\u2_Display/n4488 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u23_al_u4255  (
    .a({\u2_Display/n4460 ,\u2_Display/n4462 }),
    .b({\u2_Display/n4459 ,\u2_Display/n4461 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add137/c23 ),
    .f({\u2_Display/n4488 [25],\u2_Display/n4488 [23]}),
    .fco(\u2_Display/add137/c27 ),
    .fx({\u2_Display/n4488 [26],\u2_Display/n4488 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u27_al_u4256  (
    .a({\u2_Display/n4456 ,\u2_Display/n4458 }),
    .b({\u2_Display/n4455 ,\u2_Display/n4457 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add137/c27 ),
    .f({\u2_Display/n4488 [29],\u2_Display/n4488 [27]}),
    .fco(\u2_Display/add137/c31 ),
    .fx({\u2_Display/n4488 [30],\u2_Display/n4488 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u31_al_u4257  (
    .a({open_n54282,\u2_Display/n4454 }),
    .c(2'b00),
    .d({open_n54287,1'b1}),
    .fci(\u2_Display/add137/c31 ),
    .f({open_n54304,\u2_Display/n4488 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u3_al_u4250  (
    .a({\u2_Display/n4480 ,\u2_Display/n4482 }),
    .b({\u2_Display/n4479 ,\u2_Display/n4481 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add137/c3 ),
    .f({\u2_Display/n4488 [5],\u2_Display/n4488 [3]}),
    .fco(\u2_Display/add137/c7 ),
    .fx({\u2_Display/n4488 [6],\u2_Display/n4488 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u7_al_u4251  (
    .a({\u2_Display/n4476 ,\u2_Display/n4478 }),
    .b({\u2_Display/n4475 ,\u2_Display/n4477 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add137/c7 ),
    .f({\u2_Display/n4488 [9],\u2_Display/n4488 [7]}),
    .fco(\u2_Display/add137/c11 ),
    .fx({\u2_Display/n4488 [10],\u2_Display/n4488 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/ucin_al_u4249  (
    .a({\u2_Display/n4484 ,1'b1}),
    .b({\u2_Display/n4483 ,\u2_Display/n4485 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4488 [1],open_n54363}),
    .fco(\u2_Display/add137/c3 ),
    .fx({\u2_Display/n4488 [2],\u2_Display/n4488 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u11_al_u4261  (
    .a({\u2_Display/n4507 ,\u2_Display/n4509 }),
    .b({\u2_Display/n4506 ,\u2_Display/n4508 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add138/c11 ),
    .f({\u2_Display/n4523 [13],\u2_Display/n4523 [11]}),
    .fco(\u2_Display/add138/c15 ),
    .fx({\u2_Display/n4523 [14],\u2_Display/n4523 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u15_al_u4262  (
    .a({\u2_Display/n4503 ,\u2_Display/n4505 }),
    .b({\u2_Display/n4502 ,\u2_Display/n4504 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add138/c15 ),
    .f({\u2_Display/n4523 [17],\u2_Display/n4523 [15]}),
    .fco(\u2_Display/add138/c19 ),
    .fx({\u2_Display/n4523 [18],\u2_Display/n4523 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u19_al_u4263  (
    .a({\u2_Display/n4499 ,\u2_Display/n4501 }),
    .b({\u2_Display/n4498 ,\u2_Display/n4500 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add138/c19 ),
    .f({\u2_Display/n4523 [21],\u2_Display/n4523 [19]}),
    .fco(\u2_Display/add138/c23 ),
    .fx({\u2_Display/n4523 [22],\u2_Display/n4523 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u23_al_u4264  (
    .a({\u2_Display/n4495 ,\u2_Display/n4497 }),
    .b({\u2_Display/n4494 ,\u2_Display/n4496 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add138/c23 ),
    .f({\u2_Display/n4523 [25],\u2_Display/n4523 [23]}),
    .fco(\u2_Display/add138/c27 ),
    .fx({\u2_Display/n4523 [26],\u2_Display/n4523 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u27_al_u4265  (
    .a({\u2_Display/n4491 ,\u2_Display/n4493 }),
    .b({\u2_Display/n4490 ,\u2_Display/n4492 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add138/c27 ),
    .f({\u2_Display/n4523 [29],\u2_Display/n4523 [27]}),
    .fco(\u2_Display/add138/c31 ),
    .fx({\u2_Display/n4523 [30],\u2_Display/n4523 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u31_al_u4266  (
    .a({open_n54456,\u2_Display/n4489 }),
    .c(2'b00),
    .d({open_n54461,1'b1}),
    .fci(\u2_Display/add138/c31 ),
    .f({open_n54478,\u2_Display/n4523 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u3_al_u4259  (
    .a({\u2_Display/n4515 ,\u2_Display/n4517 }),
    .b({\u2_Display/n4514 ,\u2_Display/n4516 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add138/c3 ),
    .f({\u2_Display/n4523 [5],\u2_Display/n4523 [3]}),
    .fco(\u2_Display/add138/c7 ),
    .fx({\u2_Display/n4523 [6],\u2_Display/n4523 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u7_al_u4260  (
    .a({\u2_Display/n4511 ,\u2_Display/n4513 }),
    .b({\u2_Display/n4510 ,\u2_Display/n4512 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add138/c7 ),
    .f({\u2_Display/n4523 [9],\u2_Display/n4523 [7]}),
    .fco(\u2_Display/add138/c11 ),
    .fx({\u2_Display/n4523 [10],\u2_Display/n4523 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/ucin_al_u4258  (
    .a({\u2_Display/n4519 ,1'b1}),
    .b({\u2_Display/n4518 ,\u2_Display/n4520 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4523 [1],open_n54537}),
    .fco(\u2_Display/add138/c3 ),
    .fx({\u2_Display/n4523 [2],\u2_Display/n4523 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add139/ucin_al_u5046"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add139/u3_al_u5047  (
    .a({\u2_Display/n4550 ,\u2_Display/n4552 }),
    .b({\u2_Display/n4549 ,\u2_Display/n4551 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add139/c3 ),
    .f({\u2_Display/n4558 [5],\u2_Display/n4558 [3]}),
    .fco(\u2_Display/add139/c7 ),
    .fx({\u2_Display/n4558 [6],\u2_Display/n4558 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add139/ucin_al_u5046"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add139/u7_al_u5048  (
    .a({\u2_Display/n4546 ,\u2_Display/n4548 }),
    .b({open_n54558,\u2_Display/n4547 }),
    .c(2'b00),
    .d(2'b01),
    .e({open_n54561,1'b0}),
    .fci(\u2_Display/add139/c7 ),
    .f({\u2_Display/n4558 [9],\u2_Display/n4558 [7]}),
    .fx({open_n54577,\u2_Display/n4558 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add139/ucin_al_u5046"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add139/ucin_al_u5046  (
    .a({\u2_Display/n4554 ,1'b1}),
    .b({\u2_Display/n4553 ,\u2_Display/n4555 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4558 [1],open_n54597}),
    .fco(\u2_Display/add139/c3 ),
    .fx({\u2_Display/n4558 [2],\u2_Display/n4558 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u11_al_u4270  (
    .a({\u2_Display/counta [13],\u2_Display/counta [11]}),
    .b({\u2_Display/counta [14],\u2_Display/counta [12]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add14/c11 ),
    .f({\u2_Display/n4911 [13],\u2_Display/n4911 [11]}),
    .fco(\u2_Display/add14/c15 ),
    .fx({\u2_Display/n4911 [14],\u2_Display/n4911 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u15_al_u4271  (
    .a({\u2_Display/counta [17],\u2_Display/counta [15]}),
    .b({\u2_Display/counta [18],\u2_Display/counta [16]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add14/c15 ),
    .f({\u2_Display/n4911 [17],\u2_Display/n4911 [15]}),
    .fco(\u2_Display/add14/c19 ),
    .fx({\u2_Display/n4911 [18],\u2_Display/n4911 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u19_al_u4272  (
    .a({\u2_Display/counta [21],\u2_Display/counta [19]}),
    .b({\u2_Display/counta [22],\u2_Display/counta [20]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add14/c19 ),
    .f({\u2_Display/n4911 [21],\u2_Display/n4911 [19]}),
    .fco(\u2_Display/add14/c23 ),
    .fx({\u2_Display/n4911 [22],\u2_Display/n4911 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u23_al_u4273  (
    .a({\u2_Display/counta [25],\u2_Display/counta [23]}),
    .b({\u2_Display/counta [26],\u2_Display/counta [24]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add14/c23 ),
    .f({\u2_Display/n4911 [25],\u2_Display/n4911 [23]}),
    .fco(\u2_Display/add14/c27 ),
    .fx({\u2_Display/n4911 [26],\u2_Display/n4911 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u27_al_u4274  (
    .a({\u2_Display/counta [29],\u2_Display/counta [27]}),
    .b({\u2_Display/counta [30],\u2_Display/counta [28]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add14/c27 ),
    .f({\u2_Display/n4911 [29],\u2_Display/n4911 [27]}),
    .fco(\u2_Display/add14/c31 ),
    .fx({\u2_Display/n4911 [30],\u2_Display/n4911 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u31_al_u4275  (
    .a({open_n54690,\u2_Display/counta [31]}),
    .c(2'b00),
    .d({open_n54695,1'b0}),
    .fci(\u2_Display/add14/c31 ),
    .f({open_n54712,\u2_Display/n4911 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u3_al_u4268  (
    .a({\u2_Display/counta [5],\u2_Display/counta [3]}),
    .b({\u2_Display/counta [6],\u2_Display/counta [4]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add14/c3 ),
    .f({\u2_Display/n4911 [5],\u2_Display/n4911 [3]}),
    .fco(\u2_Display/add14/c7 ),
    .fx({\u2_Display/n4911 [6],\u2_Display/n4911 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u7_al_u4269  (
    .a({\u2_Display/counta [9],\u2_Display/counta [7]}),
    .b({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add14/c7 ),
    .f({\u2_Display/n4911 [9],\u2_Display/n4911 [7]}),
    .fco(\u2_Display/add14/c11 ),
    .fx({\u2_Display/n4911 [10],\u2_Display/n4911 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/ucin_al_u4267  (
    .a({\u2_Display/counta [1],1'b1}),
    .b({\u2_Display/counta [2],\u2_Display/counta [0]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4911 [1],open_n54771}),
    .fco(\u2_Display/add14/c3 ),
    .fx({\u2_Display/n4911 [2],\u2_Display/n4911 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u11_al_u4279  (
    .a({\u2_Display/n6088 ,\u2_Display/n6090 }),
    .b({\u2_Display/n6087 ,\u2_Display/n6089 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add151/c11 ),
    .f({\u2_Display/n4946 [13],\u2_Display/n4946 [11]}),
    .fco(\u2_Display/add151/c15 ),
    .fx({\u2_Display/n4946 [14],\u2_Display/n4946 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u15_al_u4280  (
    .a({\u2_Display/n6084 ,\u2_Display/n6086 }),
    .b({\u2_Display/n6083 ,\u2_Display/n6085 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add151/c15 ),
    .f({\u2_Display/n4946 [17],\u2_Display/n4946 [15]}),
    .fco(\u2_Display/add151/c19 ),
    .fx({\u2_Display/n4946 [18],\u2_Display/n4946 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u19_al_u4281  (
    .a({\u2_Display/n6080 ,\u2_Display/n6082 }),
    .b({\u2_Display/n6079 ,\u2_Display/n6081 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add151/c19 ),
    .f({\u2_Display/n4946 [21],\u2_Display/n4946 [19]}),
    .fco(\u2_Display/add151/c23 ),
    .fx({\u2_Display/n4946 [22],\u2_Display/n4946 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u23_al_u4282  (
    .a({\u2_Display/n6076 ,\u2_Display/n6078 }),
    .b({\u2_Display/n6075 ,\u2_Display/n6077 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add151/c23 ),
    .f({\u2_Display/n4946 [25],\u2_Display/n4946 [23]}),
    .fco(\u2_Display/add151/c27 ),
    .fx({\u2_Display/n4946 [26],\u2_Display/n4946 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u27_al_u4283  (
    .a({\u2_Display/n6072 ,\u2_Display/n6074 }),
    .b({\u2_Display/n6071 ,\u2_Display/n6073 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add151/c27 ),
    .f({\u2_Display/n4946 [29],\u2_Display/n4946 [27]}),
    .fco(\u2_Display/add151/c31 ),
    .fx({\u2_Display/n4946 [30],\u2_Display/n4946 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u31_al_u4284  (
    .a({open_n54864,\u2_Display/n6070 }),
    .c(2'b00),
    .d({open_n54869,1'b1}),
    .fci(\u2_Display/add151/c31 ),
    .f({open_n54886,\u2_Display/n4946 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u3_al_u4277  (
    .a({\u2_Display/n6096 ,\u2_Display/n6098 }),
    .b({\u2_Display/n6095 ,\u2_Display/n6097 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add151/c3 ),
    .f({\u2_Display/n4946 [5],\u2_Display/n4946 [3]}),
    .fco(\u2_Display/add151/c7 ),
    .fx({\u2_Display/n4946 [6],\u2_Display/n4946 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u7_al_u4278  (
    .a({\u2_Display/n6092 ,\u2_Display/n6094 }),
    .b({\u2_Display/n6091 ,\u2_Display/n6093 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add151/c7 ),
    .f({\u2_Display/n4946 [9],\u2_Display/n4946 [7]}),
    .fco(\u2_Display/add151/c11 ),
    .fx({\u2_Display/n4946 [10],\u2_Display/n4946 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/ucin_al_u4276  (
    .a({\u2_Display/n6100 ,1'b1}),
    .b({\u2_Display/n6099 ,\u2_Display/n6101 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4946 [1],open_n54945}),
    .fco(\u2_Display/add151/c3 ),
    .fx({\u2_Display/n4946 [2],\u2_Display/n4946 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u11_al_u4288  (
    .a({\u2_Display/n6123 ,\u2_Display/n6125 }),
    .b({\u2_Display/n6122 ,\u2_Display/n6124 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add152/c11 ),
    .f({\u2_Display/n4981 [13],\u2_Display/n4981 [11]}),
    .fco(\u2_Display/add152/c15 ),
    .fx({\u2_Display/n4981 [14],\u2_Display/n4981 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u15_al_u4289  (
    .a({\u2_Display/n6119 ,\u2_Display/n6121 }),
    .b({\u2_Display/n6118 ,\u2_Display/n6120 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add152/c15 ),
    .f({\u2_Display/n4981 [17],\u2_Display/n4981 [15]}),
    .fco(\u2_Display/add152/c19 ),
    .fx({\u2_Display/n4981 [18],\u2_Display/n4981 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u19_al_u4290  (
    .a({\u2_Display/n6115 ,\u2_Display/n6117 }),
    .b({\u2_Display/n6114 ,\u2_Display/n6116 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add152/c19 ),
    .f({\u2_Display/n4981 [21],\u2_Display/n4981 [19]}),
    .fco(\u2_Display/add152/c23 ),
    .fx({\u2_Display/n4981 [22],\u2_Display/n4981 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u23_al_u4291  (
    .a({\u2_Display/n6111 ,\u2_Display/n6113 }),
    .b({\u2_Display/n6110 ,\u2_Display/n6112 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add152/c23 ),
    .f({\u2_Display/n4981 [25],\u2_Display/n4981 [23]}),
    .fco(\u2_Display/add152/c27 ),
    .fx({\u2_Display/n4981 [26],\u2_Display/n4981 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u27_al_u4292  (
    .a({\u2_Display/n6107 ,\u2_Display/n6109 }),
    .b({\u2_Display/n6106 ,\u2_Display/n6108 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add152/c27 ),
    .f({\u2_Display/n4981 [29],\u2_Display/n4981 [27]}),
    .fco(\u2_Display/add152/c31 ),
    .fx({\u2_Display/n4981 [30],\u2_Display/n4981 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u31_al_u4293  (
    .a({open_n55038,\u2_Display/n6105 }),
    .c(2'b00),
    .d({open_n55043,1'b1}),
    .fci(\u2_Display/add152/c31 ),
    .f({open_n55060,\u2_Display/n4981 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u3_al_u4286  (
    .a({\u2_Display/n6131 ,\u2_Display/n6133 }),
    .b({\u2_Display/n6130 ,\u2_Display/n6132 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add152/c3 ),
    .f({\u2_Display/n4981 [5],\u2_Display/n4981 [3]}),
    .fco(\u2_Display/add152/c7 ),
    .fx({\u2_Display/n4981 [6],\u2_Display/n4981 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u7_al_u4287  (
    .a({\u2_Display/n6127 ,\u2_Display/n6129 }),
    .b({\u2_Display/n6126 ,\u2_Display/n6128 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add152/c7 ),
    .f({\u2_Display/n4981 [9],\u2_Display/n4981 [7]}),
    .fco(\u2_Display/add152/c11 ),
    .fx({\u2_Display/n4981 [10],\u2_Display/n4981 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/ucin_al_u4285  (
    .a({\u2_Display/n6135 ,1'b1}),
    .b({\u2_Display/n6134 ,\u2_Display/n6136 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4981 [1],open_n55119}),
    .fco(\u2_Display/add152/c3 ),
    .fx({\u2_Display/n4981 [2],\u2_Display/n4981 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u11_al_u4297  (
    .a({\u2_Display/n6158 ,\u2_Display/n6160 }),
    .b({\u2_Display/n6157 ,\u2_Display/n6159 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add153/c11 ),
    .f({\u2_Display/n5016 [13],\u2_Display/n5016 [11]}),
    .fco(\u2_Display/add153/c15 ),
    .fx({\u2_Display/n5016 [14],\u2_Display/n5016 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u15_al_u4298  (
    .a({\u2_Display/n6154 ,\u2_Display/n6156 }),
    .b({\u2_Display/n6153 ,\u2_Display/n6155 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add153/c15 ),
    .f({\u2_Display/n5016 [17],\u2_Display/n5016 [15]}),
    .fco(\u2_Display/add153/c19 ),
    .fx({\u2_Display/n5016 [18],\u2_Display/n5016 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u19_al_u4299  (
    .a({\u2_Display/n6150 ,\u2_Display/n6152 }),
    .b({\u2_Display/n6149 ,\u2_Display/n6151 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add153/c19 ),
    .f({\u2_Display/n5016 [21],\u2_Display/n5016 [19]}),
    .fco(\u2_Display/add153/c23 ),
    .fx({\u2_Display/n5016 [22],\u2_Display/n5016 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u23_al_u4300  (
    .a({\u2_Display/n6146 ,\u2_Display/n6148 }),
    .b({\u2_Display/n6145 ,\u2_Display/n6147 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add153/c23 ),
    .f({\u2_Display/n5016 [25],\u2_Display/n5016 [23]}),
    .fco(\u2_Display/add153/c27 ),
    .fx({\u2_Display/n5016 [26],\u2_Display/n5016 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u27_al_u4301  (
    .a({\u2_Display/n6142 ,\u2_Display/n6144 }),
    .b({\u2_Display/n6141 ,\u2_Display/n6143 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add153/c27 ),
    .f({\u2_Display/n5016 [29],\u2_Display/n5016 [27]}),
    .fco(\u2_Display/add153/c31 ),
    .fx({\u2_Display/n5016 [30],\u2_Display/n5016 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u31_al_u4302  (
    .a({open_n55212,\u2_Display/n6140 }),
    .c(2'b00),
    .d({open_n55217,1'b1}),
    .fci(\u2_Display/add153/c31 ),
    .f({open_n55234,\u2_Display/n5016 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u3_al_u4295  (
    .a({\u2_Display/n6166 ,\u2_Display/n6168 }),
    .b({\u2_Display/n6165 ,\u2_Display/n6167 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add153/c3 ),
    .f({\u2_Display/n5016 [5],\u2_Display/n5016 [3]}),
    .fco(\u2_Display/add153/c7 ),
    .fx({\u2_Display/n5016 [6],\u2_Display/n5016 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u7_al_u4296  (
    .a({\u2_Display/n6162 ,\u2_Display/n6164 }),
    .b({\u2_Display/n6161 ,\u2_Display/n6163 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add153/c7 ),
    .f({\u2_Display/n5016 [9],\u2_Display/n5016 [7]}),
    .fco(\u2_Display/add153/c11 ),
    .fx({\u2_Display/n5016 [10],\u2_Display/n5016 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/ucin_al_u4294  (
    .a({\u2_Display/n6170 ,1'b1}),
    .b({\u2_Display/n6169 ,\u2_Display/n6171 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5016 [1],open_n55293}),
    .fco(\u2_Display/add153/c3 ),
    .fx({\u2_Display/n5016 [2],\u2_Display/n5016 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u11_al_u4306  (
    .a({\u2_Display/n6193 ,\u2_Display/n6195 }),
    .b({\u2_Display/n6192 ,\u2_Display/n6194 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add154/c11 ),
    .f({\u2_Display/n5051 [13],\u2_Display/n5051 [11]}),
    .fco(\u2_Display/add154/c15 ),
    .fx({\u2_Display/n5051 [14],\u2_Display/n5051 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u15_al_u4307  (
    .a({\u2_Display/n6189 ,\u2_Display/n6191 }),
    .b({\u2_Display/n6188 ,\u2_Display/n6190 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add154/c15 ),
    .f({\u2_Display/n5051 [17],\u2_Display/n5051 [15]}),
    .fco(\u2_Display/add154/c19 ),
    .fx({\u2_Display/n5051 [18],\u2_Display/n5051 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u19_al_u4308  (
    .a({\u2_Display/n6185 ,\u2_Display/n6187 }),
    .b({\u2_Display/n6184 ,\u2_Display/n6186 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add154/c19 ),
    .f({\u2_Display/n5051 [21],\u2_Display/n5051 [19]}),
    .fco(\u2_Display/add154/c23 ),
    .fx({\u2_Display/n5051 [22],\u2_Display/n5051 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u23_al_u4309  (
    .a({\u2_Display/n6181 ,\u2_Display/n6183 }),
    .b({\u2_Display/n6180 ,\u2_Display/n6182 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add154/c23 ),
    .f({\u2_Display/n5051 [25],\u2_Display/n5051 [23]}),
    .fco(\u2_Display/add154/c27 ),
    .fx({\u2_Display/n5051 [26],\u2_Display/n5051 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u27_al_u4310  (
    .a({\u2_Display/n6177 ,\u2_Display/n6179 }),
    .b({\u2_Display/n6176 ,\u2_Display/n6178 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add154/c27 ),
    .f({\u2_Display/n5051 [29],\u2_Display/n5051 [27]}),
    .fco(\u2_Display/add154/c31 ),
    .fx({\u2_Display/n5051 [30],\u2_Display/n5051 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u31_al_u4311  (
    .a({open_n55386,\u2_Display/n6175 }),
    .c(2'b00),
    .d({open_n55391,1'b1}),
    .fci(\u2_Display/add154/c31 ),
    .f({open_n55408,\u2_Display/n5051 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u3_al_u4304  (
    .a({\u2_Display/n6201 ,\u2_Display/n6203 }),
    .b({\u2_Display/n6200 ,\u2_Display/n6202 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add154/c3 ),
    .f({\u2_Display/n5051 [5],\u2_Display/n5051 [3]}),
    .fco(\u2_Display/add154/c7 ),
    .fx({\u2_Display/n5051 [6],\u2_Display/n5051 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u7_al_u4305  (
    .a({\u2_Display/n6197 ,\u2_Display/n6199 }),
    .b({\u2_Display/n6196 ,\u2_Display/n6198 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add154/c7 ),
    .f({\u2_Display/n5051 [9],\u2_Display/n5051 [7]}),
    .fco(\u2_Display/add154/c11 ),
    .fx({\u2_Display/n5051 [10],\u2_Display/n5051 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/ucin_al_u4303  (
    .a({\u2_Display/n6205 ,1'b1}),
    .b({\u2_Display/n6204 ,\u2_Display/n6206 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5051 [1],open_n55467}),
    .fco(\u2_Display/add154/c3 ),
    .fx({\u2_Display/n5051 [2],\u2_Display/n5051 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u11_al_u4315  (
    .a({\u2_Display/n6228 ,\u2_Display/n6230 }),
    .b({\u2_Display/n6227 ,\u2_Display/n6229 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add155/c11 ),
    .f({\u2_Display/n5086 [13],\u2_Display/n5086 [11]}),
    .fco(\u2_Display/add155/c15 ),
    .fx({\u2_Display/n5086 [14],\u2_Display/n5086 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u15_al_u4316  (
    .a({\u2_Display/n6224 ,\u2_Display/n6226 }),
    .b({\u2_Display/n6223 ,\u2_Display/n6225 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add155/c15 ),
    .f({\u2_Display/n5086 [17],\u2_Display/n5086 [15]}),
    .fco(\u2_Display/add155/c19 ),
    .fx({\u2_Display/n5086 [18],\u2_Display/n5086 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u19_al_u4317  (
    .a({\u2_Display/n6220 ,\u2_Display/n6222 }),
    .b({\u2_Display/n6219 ,\u2_Display/n6221 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add155/c19 ),
    .f({\u2_Display/n5086 [21],\u2_Display/n5086 [19]}),
    .fco(\u2_Display/add155/c23 ),
    .fx({\u2_Display/n5086 [22],\u2_Display/n5086 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u23_al_u4318  (
    .a({\u2_Display/n6216 ,\u2_Display/n6218 }),
    .b({\u2_Display/n6215 ,\u2_Display/n6217 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add155/c23 ),
    .f({\u2_Display/n5086 [25],\u2_Display/n5086 [23]}),
    .fco(\u2_Display/add155/c27 ),
    .fx({\u2_Display/n5086 [26],\u2_Display/n5086 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u27_al_u4319  (
    .a({\u2_Display/n6212 ,\u2_Display/n6214 }),
    .b({\u2_Display/n6211 ,\u2_Display/n6213 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add155/c27 ),
    .f({\u2_Display/n5086 [29],\u2_Display/n5086 [27]}),
    .fco(\u2_Display/add155/c31 ),
    .fx({\u2_Display/n5086 [30],\u2_Display/n5086 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u31_al_u4320  (
    .a({open_n55560,\u2_Display/n6210 }),
    .c(2'b00),
    .d({open_n55565,1'b1}),
    .fci(\u2_Display/add155/c31 ),
    .f({open_n55582,\u2_Display/n5086 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u3_al_u4313  (
    .a({\u2_Display/n6236 ,\u2_Display/n6238 }),
    .b({\u2_Display/n6235 ,\u2_Display/n6237 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add155/c3 ),
    .f({\u2_Display/n5086 [5],\u2_Display/n5086 [3]}),
    .fco(\u2_Display/add155/c7 ),
    .fx({\u2_Display/n5086 [6],\u2_Display/n5086 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u7_al_u4314  (
    .a({\u2_Display/n6232 ,\u2_Display/n6234 }),
    .b({\u2_Display/n6231 ,\u2_Display/n6233 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add155/c7 ),
    .f({\u2_Display/n5086 [9],\u2_Display/n5086 [7]}),
    .fco(\u2_Display/add155/c11 ),
    .fx({\u2_Display/n5086 [10],\u2_Display/n5086 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/ucin_al_u4312  (
    .a({\u2_Display/n6240 ,1'b1}),
    .b({\u2_Display/n6239 ,\u2_Display/n6241 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5086 [1],open_n55641}),
    .fco(\u2_Display/add155/c3 ),
    .fx({\u2_Display/n5086 [2],\u2_Display/n5086 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u11_al_u4324  (
    .a({\u2_Display/n6263 ,\u2_Display/n6265 }),
    .b({\u2_Display/n6262 ,\u2_Display/n6264 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add156/c11 ),
    .f({\u2_Display/n5121 [13],\u2_Display/n5121 [11]}),
    .fco(\u2_Display/add156/c15 ),
    .fx({\u2_Display/n5121 [14],\u2_Display/n5121 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u15_al_u4325  (
    .a({\u2_Display/n6259 ,\u2_Display/n6261 }),
    .b({\u2_Display/n6258 ,\u2_Display/n6260 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add156/c15 ),
    .f({\u2_Display/n5121 [17],\u2_Display/n5121 [15]}),
    .fco(\u2_Display/add156/c19 ),
    .fx({\u2_Display/n5121 [18],\u2_Display/n5121 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u19_al_u4326  (
    .a({\u2_Display/n6255 ,\u2_Display/n6257 }),
    .b({\u2_Display/n6254 ,\u2_Display/n6256 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add156/c19 ),
    .f({\u2_Display/n5121 [21],\u2_Display/n5121 [19]}),
    .fco(\u2_Display/add156/c23 ),
    .fx({\u2_Display/n5121 [22],\u2_Display/n5121 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u23_al_u4327  (
    .a({\u2_Display/n6251 ,\u2_Display/n6253 }),
    .b({\u2_Display/n6250 ,\u2_Display/n6252 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add156/c23 ),
    .f({\u2_Display/n5121 [25],\u2_Display/n5121 [23]}),
    .fco(\u2_Display/add156/c27 ),
    .fx({\u2_Display/n5121 [26],\u2_Display/n5121 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u27_al_u4328  (
    .a({\u2_Display/n6247 ,\u2_Display/n6249 }),
    .b({\u2_Display/n6246 ,\u2_Display/n6248 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add156/c27 ),
    .f({\u2_Display/n5121 [29],\u2_Display/n5121 [27]}),
    .fco(\u2_Display/add156/c31 ),
    .fx({\u2_Display/n5121 [30],\u2_Display/n5121 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u31_al_u4329  (
    .a({open_n55734,\u2_Display/n6245 }),
    .c(2'b00),
    .d({open_n55739,1'b1}),
    .fci(\u2_Display/add156/c31 ),
    .f({open_n55756,\u2_Display/n5121 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u3_al_u4322  (
    .a({\u2_Display/n6271 ,\u2_Display/n6273 }),
    .b({\u2_Display/n6270 ,\u2_Display/n6272 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add156/c3 ),
    .f({\u2_Display/n5121 [5],\u2_Display/n5121 [3]}),
    .fco(\u2_Display/add156/c7 ),
    .fx({\u2_Display/n5121 [6],\u2_Display/n5121 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u7_al_u4323  (
    .a({\u2_Display/n6267 ,\u2_Display/n6269 }),
    .b({\u2_Display/n6266 ,\u2_Display/n6268 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add156/c7 ),
    .f({\u2_Display/n5121 [9],\u2_Display/n5121 [7]}),
    .fco(\u2_Display/add156/c11 ),
    .fx({\u2_Display/n5121 [10],\u2_Display/n5121 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/ucin_al_u4321  (
    .a({\u2_Display/n6275 ,1'b1}),
    .b({\u2_Display/n6274 ,\u2_Display/n6276 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5121 [1],open_n55815}),
    .fco(\u2_Display/add156/c3 ),
    .fx({\u2_Display/n5121 [2],\u2_Display/n5121 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u11_al_u4333  (
    .a({\u2_Display/n6298 ,\u2_Display/n6300 }),
    .b({\u2_Display/n6297 ,\u2_Display/n6299 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add157/c11 ),
    .f({\u2_Display/n5156 [13],\u2_Display/n5156 [11]}),
    .fco(\u2_Display/add157/c15 ),
    .fx({\u2_Display/n5156 [14],\u2_Display/n5156 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u15_al_u4334  (
    .a({\u2_Display/n6294 ,\u2_Display/n6296 }),
    .b({\u2_Display/n6293 ,\u2_Display/n6295 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add157/c15 ),
    .f({\u2_Display/n5156 [17],\u2_Display/n5156 [15]}),
    .fco(\u2_Display/add157/c19 ),
    .fx({\u2_Display/n5156 [18],\u2_Display/n5156 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u19_al_u4335  (
    .a({\u2_Display/n6290 ,\u2_Display/n6292 }),
    .b({\u2_Display/n6289 ,\u2_Display/n6291 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add157/c19 ),
    .f({\u2_Display/n5156 [21],\u2_Display/n5156 [19]}),
    .fco(\u2_Display/add157/c23 ),
    .fx({\u2_Display/n5156 [22],\u2_Display/n5156 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u23_al_u4336  (
    .a({\u2_Display/n6286 ,\u2_Display/n6288 }),
    .b({\u2_Display/n6285 ,\u2_Display/n6287 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add157/c23 ),
    .f({\u2_Display/n5156 [25],\u2_Display/n5156 [23]}),
    .fco(\u2_Display/add157/c27 ),
    .fx({\u2_Display/n5156 [26],\u2_Display/n5156 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u27_al_u4337  (
    .a({\u2_Display/n6282 ,\u2_Display/n6284 }),
    .b({\u2_Display/n6281 ,\u2_Display/n6283 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add157/c27 ),
    .f({\u2_Display/n5156 [29],\u2_Display/n5156 [27]}),
    .fco(\u2_Display/add157/c31 ),
    .fx({\u2_Display/n5156 [30],\u2_Display/n5156 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u31_al_u4338  (
    .a({open_n55908,\u2_Display/n6280 }),
    .c(2'b00),
    .d({open_n55913,1'b1}),
    .fci(\u2_Display/add157/c31 ),
    .f({open_n55930,\u2_Display/n5156 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u3_al_u4331  (
    .a({\u2_Display/n6306 ,\u2_Display/n6308 }),
    .b({\u2_Display/n6305 ,\u2_Display/n6307 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add157/c3 ),
    .f({\u2_Display/n5156 [5],\u2_Display/n5156 [3]}),
    .fco(\u2_Display/add157/c7 ),
    .fx({\u2_Display/n5156 [6],\u2_Display/n5156 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u7_al_u4332  (
    .a({\u2_Display/n6302 ,\u2_Display/n6304 }),
    .b({\u2_Display/n6301 ,\u2_Display/n6303 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add157/c7 ),
    .f({\u2_Display/n5156 [9],\u2_Display/n5156 [7]}),
    .fco(\u2_Display/add157/c11 ),
    .fx({\u2_Display/n5156 [10],\u2_Display/n5156 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/ucin_al_u4330  (
    .a({\u2_Display/n6310 ,1'b1}),
    .b({\u2_Display/n6309 ,\u2_Display/n6311 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5156 [1],open_n55989}),
    .fco(\u2_Display/add157/c3 ),
    .fx({\u2_Display/n5156 [2],\u2_Display/n5156 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u11_al_u4342  (
    .a({\u2_Display/n6333 ,\u2_Display/n6335 }),
    .b({\u2_Display/n6332 ,\u2_Display/n6334 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add158/c11 ),
    .f({\u2_Display/n5191 [13],\u2_Display/n5191 [11]}),
    .fco(\u2_Display/add158/c15 ),
    .fx({\u2_Display/n5191 [14],\u2_Display/n5191 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u15_al_u4343  (
    .a({\u2_Display/n6329 ,\u2_Display/n6331 }),
    .b({\u2_Display/n6328 ,\u2_Display/n6330 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add158/c15 ),
    .f({\u2_Display/n5191 [17],\u2_Display/n5191 [15]}),
    .fco(\u2_Display/add158/c19 ),
    .fx({\u2_Display/n5191 [18],\u2_Display/n5191 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u19_al_u4344  (
    .a({\u2_Display/n6325 ,\u2_Display/n6327 }),
    .b({\u2_Display/n6324 ,\u2_Display/n6326 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add158/c19 ),
    .f({\u2_Display/n5191 [21],\u2_Display/n5191 [19]}),
    .fco(\u2_Display/add158/c23 ),
    .fx({\u2_Display/n5191 [22],\u2_Display/n5191 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u23_al_u4345  (
    .a({\u2_Display/n6321 ,\u2_Display/n6323 }),
    .b({\u2_Display/n6320 ,\u2_Display/n6322 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add158/c23 ),
    .f({\u2_Display/n5191 [25],\u2_Display/n5191 [23]}),
    .fco(\u2_Display/add158/c27 ),
    .fx({\u2_Display/n5191 [26],\u2_Display/n5191 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u27_al_u4346  (
    .a({\u2_Display/n6317 ,\u2_Display/n6319 }),
    .b({\u2_Display/n6316 ,\u2_Display/n6318 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add158/c27 ),
    .f({\u2_Display/n5191 [29],\u2_Display/n5191 [27]}),
    .fco(\u2_Display/add158/c31 ),
    .fx({\u2_Display/n5191 [30],\u2_Display/n5191 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u31_al_u4347  (
    .a({open_n56082,\u2_Display/n6315 }),
    .c(2'b00),
    .d({open_n56087,1'b1}),
    .fci(\u2_Display/add158/c31 ),
    .f({open_n56104,\u2_Display/n5191 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u3_al_u4340  (
    .a({\u2_Display/n6341 ,\u2_Display/n6343 }),
    .b({\u2_Display/n6340 ,\u2_Display/n6342 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add158/c3 ),
    .f({\u2_Display/n5191 [5],\u2_Display/n5191 [3]}),
    .fco(\u2_Display/add158/c7 ),
    .fx({\u2_Display/n5191 [6],\u2_Display/n5191 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u7_al_u4341  (
    .a({\u2_Display/n6337 ,\u2_Display/n6339 }),
    .b({\u2_Display/n6336 ,\u2_Display/n6338 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add158/c7 ),
    .f({\u2_Display/n5191 [9],\u2_Display/n5191 [7]}),
    .fco(\u2_Display/add158/c11 ),
    .fx({\u2_Display/n5191 [10],\u2_Display/n5191 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/ucin_al_u4339  (
    .a({\u2_Display/n6345 ,1'b1}),
    .b({\u2_Display/n6344 ,\u2_Display/n6346 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5191 [1],open_n56163}),
    .fco(\u2_Display/add158/c3 ),
    .fx({\u2_Display/n5191 [2],\u2_Display/n5191 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u11_al_u4351  (
    .a({\u2_Display/n5210 ,\u2_Display/n5212 }),
    .b({\u2_Display/n5209 ,\u2_Display/n5211 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add159/c11 ),
    .f({\u2_Display/n5226 [13],\u2_Display/n5226 [11]}),
    .fco(\u2_Display/add159/c15 ),
    .fx({\u2_Display/n5226 [14],\u2_Display/n5226 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u15_al_u4352  (
    .a({\u2_Display/n5206 ,\u2_Display/n5208 }),
    .b({\u2_Display/n5205 ,\u2_Display/n5207 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add159/c15 ),
    .f({\u2_Display/n5226 [17],\u2_Display/n5226 [15]}),
    .fco(\u2_Display/add159/c19 ),
    .fx({\u2_Display/n5226 [18],\u2_Display/n5226 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u19_al_u4353  (
    .a({\u2_Display/n5202 ,\u2_Display/n5204 }),
    .b({\u2_Display/n5201 ,\u2_Display/n5203 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add159/c19 ),
    .f({\u2_Display/n5226 [21],\u2_Display/n5226 [19]}),
    .fco(\u2_Display/add159/c23 ),
    .fx({\u2_Display/n5226 [22],\u2_Display/n5226 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u23_al_u4354  (
    .a({\u2_Display/n5198 ,\u2_Display/n5200 }),
    .b({\u2_Display/n5197 ,\u2_Display/n5199 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add159/c23 ),
    .f({\u2_Display/n5226 [25],\u2_Display/n5226 [23]}),
    .fco(\u2_Display/add159/c27 ),
    .fx({\u2_Display/n5226 [26],\u2_Display/n5226 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u27_al_u4355  (
    .a({\u2_Display/n6352 ,\u2_Display/n5196 }),
    .b({\u2_Display/n6351 ,\u2_Display/n6353 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add159/c27 ),
    .f({\u2_Display/n5226 [29],\u2_Display/n5226 [27]}),
    .fco(\u2_Display/add159/c31 ),
    .fx({\u2_Display/n5226 [30],\u2_Display/n5226 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u31_al_u4356  (
    .a({open_n56256,\u2_Display/n6350 }),
    .c(2'b00),
    .d({open_n56261,1'b1}),
    .fci(\u2_Display/add159/c31 ),
    .f({open_n56278,\u2_Display/n5226 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u3_al_u4349  (
    .a({\u2_Display/n5218 ,\u2_Display/n5220 }),
    .b({\u2_Display/n5217 ,\u2_Display/n5219 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add159/c3 ),
    .f({\u2_Display/n5226 [5],\u2_Display/n5226 [3]}),
    .fco(\u2_Display/add159/c7 ),
    .fx({\u2_Display/n5226 [6],\u2_Display/n5226 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u7_al_u4350  (
    .a({\u2_Display/n5214 ,\u2_Display/n5216 }),
    .b({\u2_Display/n5213 ,\u2_Display/n5215 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add159/c7 ),
    .f({\u2_Display/n5226 [9],\u2_Display/n5226 [7]}),
    .fco(\u2_Display/add159/c11 ),
    .fx({\u2_Display/n5226 [10],\u2_Display/n5226 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/ucin_al_u4348  (
    .a({\u2_Display/n5222 ,1'b1}),
    .b({\u2_Display/n5221 ,\u2_Display/n5223 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5226 [1],open_n56337}),
    .fco(\u2_Display/add159/c3 ),
    .fx({\u2_Display/n5226 [2],\u2_Display/n5226 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u11_al_u4360  (
    .a({\u2_Display/n5245 ,\u2_Display/n5247 }),
    .b({\u2_Display/n5244 ,\u2_Display/n5246 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add160/c11 ),
    .f({\u2_Display/n5261 [13],\u2_Display/n5261 [11]}),
    .fco(\u2_Display/add160/c15 ),
    .fx({\u2_Display/n5261 [14],\u2_Display/n5261 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u15_al_u4361  (
    .a({\u2_Display/n5241 ,\u2_Display/n5243 }),
    .b({\u2_Display/n5240 ,\u2_Display/n5242 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add160/c15 ),
    .f({\u2_Display/n5261 [17],\u2_Display/n5261 [15]}),
    .fco(\u2_Display/add160/c19 ),
    .fx({\u2_Display/n5261 [18],\u2_Display/n5261 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u19_al_u4362  (
    .a({\u2_Display/n5237 ,\u2_Display/n5239 }),
    .b({\u2_Display/n5236 ,\u2_Display/n5238 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add160/c19 ),
    .f({\u2_Display/n5261 [21],\u2_Display/n5261 [19]}),
    .fco(\u2_Display/add160/c23 ),
    .fx({\u2_Display/n5261 [22],\u2_Display/n5261 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u23_al_u4363  (
    .a({\u2_Display/n5233 ,\u2_Display/n5235 }),
    .b({\u2_Display/n5232 ,\u2_Display/n5234 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add160/c23 ),
    .f({\u2_Display/n5261 [25],\u2_Display/n5261 [23]}),
    .fco(\u2_Display/add160/c27 ),
    .fx({\u2_Display/n5261 [26],\u2_Display/n5261 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u27_al_u4364  (
    .a({\u2_Display/n5229 ,\u2_Display/n5231 }),
    .b({\u2_Display/n5228 ,\u2_Display/n5230 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add160/c27 ),
    .f({\u2_Display/n5261 [29],\u2_Display/n5261 [27]}),
    .fco(\u2_Display/add160/c31 ),
    .fx({\u2_Display/n5261 [30],\u2_Display/n5261 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u31_al_u4365  (
    .a({open_n56430,\u2_Display/n5227 }),
    .c(2'b00),
    .d({open_n56435,1'b1}),
    .fci(\u2_Display/add160/c31 ),
    .f({open_n56452,\u2_Display/n5261 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u3_al_u4358  (
    .a({\u2_Display/n5253 ,\u2_Display/n5255 }),
    .b({\u2_Display/n5252 ,\u2_Display/n5254 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add160/c3 ),
    .f({\u2_Display/n5261 [5],\u2_Display/n5261 [3]}),
    .fco(\u2_Display/add160/c7 ),
    .fx({\u2_Display/n5261 [6],\u2_Display/n5261 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u7_al_u4359  (
    .a({\u2_Display/n5249 ,\u2_Display/n5251 }),
    .b({\u2_Display/n5248 ,\u2_Display/n5250 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add160/c7 ),
    .f({\u2_Display/n5261 [9],\u2_Display/n5261 [7]}),
    .fco(\u2_Display/add160/c11 ),
    .fx({\u2_Display/n5261 [10],\u2_Display/n5261 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/ucin_al_u4357  (
    .a({\u2_Display/n5257 ,1'b1}),
    .b({\u2_Display/n5256 ,\u2_Display/n5258 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5261 [1],open_n56511}),
    .fco(\u2_Display/add160/c3 ),
    .fx({\u2_Display/n5261 [2],\u2_Display/n5261 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u11_al_u4369  (
    .a({\u2_Display/n5280 ,\u2_Display/n5282 }),
    .b({\u2_Display/n5279 ,\u2_Display/n5281 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add161/c11 ),
    .f({\u2_Display/n5296 [13],\u2_Display/n5296 [11]}),
    .fco(\u2_Display/add161/c15 ),
    .fx({\u2_Display/n5296 [14],\u2_Display/n5296 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u15_al_u4370  (
    .a({\u2_Display/n5276 ,\u2_Display/n5278 }),
    .b({\u2_Display/n5275 ,\u2_Display/n5277 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add161/c15 ),
    .f({\u2_Display/n5296 [17],\u2_Display/n5296 [15]}),
    .fco(\u2_Display/add161/c19 ),
    .fx({\u2_Display/n5296 [18],\u2_Display/n5296 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u19_al_u4371  (
    .a({\u2_Display/n5272 ,\u2_Display/n5274 }),
    .b({\u2_Display/n5271 ,\u2_Display/n5273 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add161/c19 ),
    .f({\u2_Display/n5296 [21],\u2_Display/n5296 [19]}),
    .fco(\u2_Display/add161/c23 ),
    .fx({\u2_Display/n5296 [22],\u2_Display/n5296 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u23_al_u4372  (
    .a({\u2_Display/n5268 ,\u2_Display/n5270 }),
    .b({\u2_Display/n5267 ,\u2_Display/n5269 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add161/c23 ),
    .f({\u2_Display/n5296 [25],\u2_Display/n5296 [23]}),
    .fco(\u2_Display/add161/c27 ),
    .fx({\u2_Display/n5296 [26],\u2_Display/n5296 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u27_al_u4373  (
    .a({\u2_Display/n5264 ,\u2_Display/n5266 }),
    .b({\u2_Display/n5263 ,\u2_Display/n5265 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add161/c27 ),
    .f({\u2_Display/n5296 [29],\u2_Display/n5296 [27]}),
    .fco(\u2_Display/add161/c31 ),
    .fx({\u2_Display/n5296 [30],\u2_Display/n5296 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u31_al_u4374  (
    .a({open_n56604,\u2_Display/n5262 }),
    .c(2'b00),
    .d({open_n56609,1'b1}),
    .fci(\u2_Display/add161/c31 ),
    .f({open_n56626,\u2_Display/n5296 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u3_al_u4367  (
    .a({\u2_Display/n5288 ,\u2_Display/n5290 }),
    .b({\u2_Display/n5287 ,\u2_Display/n5289 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add161/c3 ),
    .f({\u2_Display/n5296 [5],\u2_Display/n5296 [3]}),
    .fco(\u2_Display/add161/c7 ),
    .fx({\u2_Display/n5296 [6],\u2_Display/n5296 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u7_al_u4368  (
    .a({\u2_Display/n5284 ,\u2_Display/n5286 }),
    .b({\u2_Display/n5283 ,\u2_Display/n5285 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add161/c7 ),
    .f({\u2_Display/n5296 [9],\u2_Display/n5296 [7]}),
    .fco(\u2_Display/add161/c11 ),
    .fx({\u2_Display/n5296 [10],\u2_Display/n5296 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/ucin_al_u4366  (
    .a({\u2_Display/n5292 ,1'b1}),
    .b({\u2_Display/n5291 ,\u2_Display/n5293 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5296 [1],open_n56685}),
    .fco(\u2_Display/add161/c3 ),
    .fx({\u2_Display/n5296 [2],\u2_Display/n5296 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u11_al_u4378  (
    .a({\u2_Display/n5315 ,\u2_Display/n5317 }),
    .b({\u2_Display/n5314 ,\u2_Display/n5316 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add162/c11 ),
    .f({\u2_Display/n5331 [13],\u2_Display/n5331 [11]}),
    .fco(\u2_Display/add162/c15 ),
    .fx({\u2_Display/n5331 [14],\u2_Display/n5331 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u15_al_u4379  (
    .a({\u2_Display/n5311 ,\u2_Display/n5313 }),
    .b({\u2_Display/n5310 ,\u2_Display/n5312 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add162/c15 ),
    .f({\u2_Display/n5331 [17],\u2_Display/n5331 [15]}),
    .fco(\u2_Display/add162/c19 ),
    .fx({\u2_Display/n5331 [18],\u2_Display/n5331 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u19_al_u4380  (
    .a({\u2_Display/n5307 ,\u2_Display/n5309 }),
    .b({\u2_Display/n5306 ,\u2_Display/n5308 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add162/c19 ),
    .f({\u2_Display/n5331 [21],\u2_Display/n5331 [19]}),
    .fco(\u2_Display/add162/c23 ),
    .fx({\u2_Display/n5331 [22],\u2_Display/n5331 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u23_al_u4381  (
    .a({\u2_Display/n5303 ,\u2_Display/n5305 }),
    .b({\u2_Display/n5302 ,\u2_Display/n5304 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add162/c23 ),
    .f({\u2_Display/n5331 [25],\u2_Display/n5331 [23]}),
    .fco(\u2_Display/add162/c27 ),
    .fx({\u2_Display/n5331 [26],\u2_Display/n5331 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u27_al_u4382  (
    .a({\u2_Display/n5299 ,\u2_Display/n5301 }),
    .b({\u2_Display/n5298 ,\u2_Display/n5300 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add162/c27 ),
    .f({\u2_Display/n5331 [29],\u2_Display/n5331 [27]}),
    .fco(\u2_Display/add162/c31 ),
    .fx({\u2_Display/n5331 [30],\u2_Display/n5331 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u31_al_u4383  (
    .a({open_n56778,\u2_Display/n5297 }),
    .c(2'b00),
    .d({open_n56783,1'b1}),
    .fci(\u2_Display/add162/c31 ),
    .f({open_n56800,\u2_Display/n5331 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u3_al_u4376  (
    .a({\u2_Display/n5323 ,\u2_Display/n5325 }),
    .b({\u2_Display/n5322 ,\u2_Display/n5324 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add162/c3 ),
    .f({\u2_Display/n5331 [5],\u2_Display/n5331 [3]}),
    .fco(\u2_Display/add162/c7 ),
    .fx({\u2_Display/n5331 [6],\u2_Display/n5331 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u7_al_u4377  (
    .a({\u2_Display/n5319 ,\u2_Display/n5321 }),
    .b({\u2_Display/n5318 ,\u2_Display/n5320 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add162/c7 ),
    .f({\u2_Display/n5331 [9],\u2_Display/n5331 [7]}),
    .fco(\u2_Display/add162/c11 ),
    .fx({\u2_Display/n5331 [10],\u2_Display/n5331 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/ucin_al_u4375  (
    .a({\u2_Display/n5327 ,1'b1}),
    .b({\u2_Display/n5326 ,\u2_Display/n5328 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5331 [1],open_n56859}),
    .fco(\u2_Display/add162/c3 ),
    .fx({\u2_Display/n5331 [2],\u2_Display/n5331 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u11_al_u4387  (
    .a({\u2_Display/n5350 ,\u2_Display/n5352 }),
    .b({\u2_Display/n5349 ,\u2_Display/n5351 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add163/c11 ),
    .f({\u2_Display/n5366 [13],\u2_Display/n5366 [11]}),
    .fco(\u2_Display/add163/c15 ),
    .fx({\u2_Display/n5366 [14],\u2_Display/n5366 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u15_al_u4388  (
    .a({\u2_Display/n5346 ,\u2_Display/n5348 }),
    .b({\u2_Display/n5345 ,\u2_Display/n5347 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add163/c15 ),
    .f({\u2_Display/n5366 [17],\u2_Display/n5366 [15]}),
    .fco(\u2_Display/add163/c19 ),
    .fx({\u2_Display/n5366 [18],\u2_Display/n5366 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u19_al_u4389  (
    .a({\u2_Display/n5342 ,\u2_Display/n5344 }),
    .b({\u2_Display/n5341 ,\u2_Display/n5343 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add163/c19 ),
    .f({\u2_Display/n5366 [21],\u2_Display/n5366 [19]}),
    .fco(\u2_Display/add163/c23 ),
    .fx({\u2_Display/n5366 [22],\u2_Display/n5366 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u23_al_u4390  (
    .a({\u2_Display/n5338 ,\u2_Display/n5340 }),
    .b({\u2_Display/n5337 ,\u2_Display/n5339 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add163/c23 ),
    .f({\u2_Display/n5366 [25],\u2_Display/n5366 [23]}),
    .fco(\u2_Display/add163/c27 ),
    .fx({\u2_Display/n5366 [26],\u2_Display/n5366 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u27_al_u4391  (
    .a({\u2_Display/n5334 ,\u2_Display/n5336 }),
    .b({\u2_Display/n5333 ,\u2_Display/n5335 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add163/c27 ),
    .f({\u2_Display/n5366 [29],\u2_Display/n5366 [27]}),
    .fco(\u2_Display/add163/c31 ),
    .fx({\u2_Display/n5366 [30],\u2_Display/n5366 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u31_al_u4392  (
    .a({open_n56952,\u2_Display/n5332 }),
    .c(2'b00),
    .d({open_n56957,1'b1}),
    .fci(\u2_Display/add163/c31 ),
    .f({open_n56974,\u2_Display/n5366 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u3_al_u4385  (
    .a({\u2_Display/n5358 ,\u2_Display/n5360 }),
    .b({\u2_Display/n5357 ,\u2_Display/n5359 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add163/c3 ),
    .f({\u2_Display/n5366 [5],\u2_Display/n5366 [3]}),
    .fco(\u2_Display/add163/c7 ),
    .fx({\u2_Display/n5366 [6],\u2_Display/n5366 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u7_al_u4386  (
    .a({\u2_Display/n5354 ,\u2_Display/n5356 }),
    .b({\u2_Display/n5353 ,\u2_Display/n5355 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add163/c7 ),
    .f({\u2_Display/n5366 [9],\u2_Display/n5366 [7]}),
    .fco(\u2_Display/add163/c11 ),
    .fx({\u2_Display/n5366 [10],\u2_Display/n5366 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/ucin_al_u4384  (
    .a({\u2_Display/n5362 ,1'b1}),
    .b({\u2_Display/n5361 ,\u2_Display/n5363 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5366 [1],open_n57033}),
    .fco(\u2_Display/add163/c3 ),
    .fx({\u2_Display/n5366 [2],\u2_Display/n5366 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u11_al_u4396  (
    .a({\u2_Display/n5385 ,\u2_Display/n5387 }),
    .b({\u2_Display/n5384 ,\u2_Display/n5386 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add164/c11 ),
    .f({\u2_Display/n5401 [13],\u2_Display/n5401 [11]}),
    .fco(\u2_Display/add164/c15 ),
    .fx({\u2_Display/n5401 [14],\u2_Display/n5401 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u15_al_u4397  (
    .a({\u2_Display/n5381 ,\u2_Display/n5383 }),
    .b({\u2_Display/n5380 ,\u2_Display/n5382 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add164/c15 ),
    .f({\u2_Display/n5401 [17],\u2_Display/n5401 [15]}),
    .fco(\u2_Display/add164/c19 ),
    .fx({\u2_Display/n5401 [18],\u2_Display/n5401 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u19_al_u4398  (
    .a({\u2_Display/n5377 ,\u2_Display/n5379 }),
    .b({\u2_Display/n5376 ,\u2_Display/n5378 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add164/c19 ),
    .f({\u2_Display/n5401 [21],\u2_Display/n5401 [19]}),
    .fco(\u2_Display/add164/c23 ),
    .fx({\u2_Display/n5401 [22],\u2_Display/n5401 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u23_al_u4399  (
    .a({\u2_Display/n5373 ,\u2_Display/n5375 }),
    .b({\u2_Display/n5372 ,\u2_Display/n5374 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add164/c23 ),
    .f({\u2_Display/n5401 [25],\u2_Display/n5401 [23]}),
    .fco(\u2_Display/add164/c27 ),
    .fx({\u2_Display/n5401 [26],\u2_Display/n5401 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u27_al_u4400  (
    .a({\u2_Display/n5369 ,\u2_Display/n5371 }),
    .b({\u2_Display/n5368 ,\u2_Display/n5370 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add164/c27 ),
    .f({\u2_Display/n5401 [29],\u2_Display/n5401 [27]}),
    .fco(\u2_Display/add164/c31 ),
    .fx({\u2_Display/n5401 [30],\u2_Display/n5401 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u31_al_u4401  (
    .a({open_n57126,\u2_Display/n5367 }),
    .c(2'b00),
    .d({open_n57131,1'b1}),
    .fci(\u2_Display/add164/c31 ),
    .f({open_n57148,\u2_Display/n5401 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u3_al_u4394  (
    .a({\u2_Display/n5393 ,\u2_Display/n5395 }),
    .b({\u2_Display/n5392 ,\u2_Display/n5394 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add164/c3 ),
    .f({\u2_Display/n5401 [5],\u2_Display/n5401 [3]}),
    .fco(\u2_Display/add164/c7 ),
    .fx({\u2_Display/n5401 [6],\u2_Display/n5401 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u7_al_u4395  (
    .a({\u2_Display/n5389 ,\u2_Display/n5391 }),
    .b({\u2_Display/n5388 ,\u2_Display/n5390 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add164/c7 ),
    .f({\u2_Display/n5401 [9],\u2_Display/n5401 [7]}),
    .fco(\u2_Display/add164/c11 ),
    .fx({\u2_Display/n5401 [10],\u2_Display/n5401 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/ucin_al_u4393  (
    .a({\u2_Display/n5397 ,1'b1}),
    .b({\u2_Display/n5396 ,\u2_Display/n5398 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5401 [1],open_n57207}),
    .fco(\u2_Display/add164/c3 ),
    .fx({\u2_Display/n5401 [2],\u2_Display/n5401 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u11_al_u4405  (
    .a({\u2_Display/n5420 ,\u2_Display/n5422 }),
    .b({\u2_Display/n5419 ,\u2_Display/n5421 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add165/c11 ),
    .f({\u2_Display/n5436 [13],\u2_Display/n5436 [11]}),
    .fco(\u2_Display/add165/c15 ),
    .fx({\u2_Display/n5436 [14],\u2_Display/n5436 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u15_al_u4406  (
    .a({\u2_Display/n5416 ,\u2_Display/n5418 }),
    .b({\u2_Display/n5415 ,\u2_Display/n5417 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add165/c15 ),
    .f({\u2_Display/n5436 [17],\u2_Display/n5436 [15]}),
    .fco(\u2_Display/add165/c19 ),
    .fx({\u2_Display/n5436 [18],\u2_Display/n5436 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u19_al_u4407  (
    .a({\u2_Display/n5412 ,\u2_Display/n5414 }),
    .b({\u2_Display/n5411 ,\u2_Display/n5413 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add165/c19 ),
    .f({\u2_Display/n5436 [21],\u2_Display/n5436 [19]}),
    .fco(\u2_Display/add165/c23 ),
    .fx({\u2_Display/n5436 [22],\u2_Display/n5436 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u23_al_u4408  (
    .a({\u2_Display/n5408 ,\u2_Display/n5410 }),
    .b({\u2_Display/n5407 ,\u2_Display/n5409 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add165/c23 ),
    .f({\u2_Display/n5436 [25],\u2_Display/n5436 [23]}),
    .fco(\u2_Display/add165/c27 ),
    .fx({\u2_Display/n5436 [26],\u2_Display/n5436 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u27_al_u4409  (
    .a({\u2_Display/n5404 ,\u2_Display/n5406 }),
    .b({\u2_Display/n5403 ,\u2_Display/n5405 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add165/c27 ),
    .f({\u2_Display/n5436 [29],\u2_Display/n5436 [27]}),
    .fco(\u2_Display/add165/c31 ),
    .fx({\u2_Display/n5436 [30],\u2_Display/n5436 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u31_al_u4410  (
    .a({open_n57300,\u2_Display/n5402 }),
    .c(2'b00),
    .d({open_n57305,1'b1}),
    .fci(\u2_Display/add165/c31 ),
    .f({open_n57322,\u2_Display/n5436 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u3_al_u4403  (
    .a({\u2_Display/n5428 ,\u2_Display/n5430 }),
    .b({\u2_Display/n5427 ,\u2_Display/n5429 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add165/c3 ),
    .f({\u2_Display/n5436 [5],\u2_Display/n5436 [3]}),
    .fco(\u2_Display/add165/c7 ),
    .fx({\u2_Display/n5436 [6],\u2_Display/n5436 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u7_al_u4404  (
    .a({\u2_Display/n5424 ,\u2_Display/n5426 }),
    .b({\u2_Display/n5423 ,\u2_Display/n5425 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add165/c7 ),
    .f({\u2_Display/n5436 [9],\u2_Display/n5436 [7]}),
    .fco(\u2_Display/add165/c11 ),
    .fx({\u2_Display/n5436 [10],\u2_Display/n5436 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/ucin_al_u4402  (
    .a({\u2_Display/n5432 ,1'b1}),
    .b({\u2_Display/n5431 ,\u2_Display/n5433 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5436 [1],open_n57381}),
    .fco(\u2_Display/add165/c3 ),
    .fx({\u2_Display/n5436 [2],\u2_Display/n5436 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u11_al_u4414  (
    .a({\u2_Display/n5455 ,\u2_Display/n5457 }),
    .b({\u2_Display/n5454 ,\u2_Display/n5456 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add166/c11 ),
    .f({\u2_Display/n5471 [13],\u2_Display/n5471 [11]}),
    .fco(\u2_Display/add166/c15 ),
    .fx({\u2_Display/n5471 [14],\u2_Display/n5471 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u15_al_u4415  (
    .a({\u2_Display/n5451 ,\u2_Display/n5453 }),
    .b({\u2_Display/n5450 ,\u2_Display/n5452 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add166/c15 ),
    .f({\u2_Display/n5471 [17],\u2_Display/n5471 [15]}),
    .fco(\u2_Display/add166/c19 ),
    .fx({\u2_Display/n5471 [18],\u2_Display/n5471 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u19_al_u4416  (
    .a({\u2_Display/n5447 ,\u2_Display/n5449 }),
    .b({\u2_Display/n5446 ,\u2_Display/n5448 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add166/c19 ),
    .f({\u2_Display/n5471 [21],\u2_Display/n5471 [19]}),
    .fco(\u2_Display/add166/c23 ),
    .fx({\u2_Display/n5471 [22],\u2_Display/n5471 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u23_al_u4417  (
    .a({\u2_Display/n5443 ,\u2_Display/n5445 }),
    .b({\u2_Display/n5442 ,\u2_Display/n5444 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add166/c23 ),
    .f({\u2_Display/n5471 [25],\u2_Display/n5471 [23]}),
    .fco(\u2_Display/add166/c27 ),
    .fx({\u2_Display/n5471 [26],\u2_Display/n5471 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u27_al_u4418  (
    .a({\u2_Display/n5439 ,\u2_Display/n5441 }),
    .b({\u2_Display/n5438 ,\u2_Display/n5440 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add166/c27 ),
    .f({\u2_Display/n5471 [29],\u2_Display/n5471 [27]}),
    .fco(\u2_Display/add166/c31 ),
    .fx({\u2_Display/n5471 [30],\u2_Display/n5471 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u31_al_u4419  (
    .a({open_n57474,\u2_Display/n5437 }),
    .c(2'b00),
    .d({open_n57479,1'b1}),
    .fci(\u2_Display/add166/c31 ),
    .f({open_n57496,\u2_Display/n5471 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u3_al_u4412  (
    .a({\u2_Display/n5463 ,\u2_Display/n5465 }),
    .b({\u2_Display/n5462 ,\u2_Display/n5464 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add166/c3 ),
    .f({\u2_Display/n5471 [5],\u2_Display/n5471 [3]}),
    .fco(\u2_Display/add166/c7 ),
    .fx({\u2_Display/n5471 [6],\u2_Display/n5471 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u7_al_u4413  (
    .a({\u2_Display/n5459 ,\u2_Display/n5461 }),
    .b({\u2_Display/n5458 ,\u2_Display/n5460 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add166/c7 ),
    .f({\u2_Display/n5471 [9],\u2_Display/n5471 [7]}),
    .fco(\u2_Display/add166/c11 ),
    .fx({\u2_Display/n5471 [10],\u2_Display/n5471 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/ucin_al_u4411  (
    .a({\u2_Display/n5467 ,1'b1}),
    .b({\u2_Display/n5466 ,\u2_Display/n5468 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5471 [1],open_n57555}),
    .fco(\u2_Display/add166/c3 ),
    .fx({\u2_Display/n5471 [2],\u2_Display/n5471 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u11_al_u4423  (
    .a({\u2_Display/n5490 ,\u2_Display/n5492 }),
    .b({\u2_Display/n5489 ,\u2_Display/n5491 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add167/c11 ),
    .f({\u2_Display/n5506 [13],\u2_Display/n5506 [11]}),
    .fco(\u2_Display/add167/c15 ),
    .fx({\u2_Display/n5506 [14],\u2_Display/n5506 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u15_al_u4424  (
    .a({\u2_Display/n5486 ,\u2_Display/n5488 }),
    .b({\u2_Display/n5485 ,\u2_Display/n5487 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add167/c15 ),
    .f({\u2_Display/n5506 [17],\u2_Display/n5506 [15]}),
    .fco(\u2_Display/add167/c19 ),
    .fx({\u2_Display/n5506 [18],\u2_Display/n5506 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u19_al_u4425  (
    .a({\u2_Display/n5482 ,\u2_Display/n5484 }),
    .b({\u2_Display/n5481 ,\u2_Display/n5483 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add167/c19 ),
    .f({\u2_Display/n5506 [21],\u2_Display/n5506 [19]}),
    .fco(\u2_Display/add167/c23 ),
    .fx({\u2_Display/n5506 [22],\u2_Display/n5506 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u23_al_u4426  (
    .a({\u2_Display/n5478 ,\u2_Display/n5480 }),
    .b({\u2_Display/n5477 ,\u2_Display/n5479 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add167/c23 ),
    .f({\u2_Display/n5506 [25],\u2_Display/n5506 [23]}),
    .fco(\u2_Display/add167/c27 ),
    .fx({\u2_Display/n5506 [26],\u2_Display/n5506 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u27_al_u4427  (
    .a({\u2_Display/n5474 ,\u2_Display/n5476 }),
    .b({\u2_Display/n5473 ,\u2_Display/n5475 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add167/c27 ),
    .f({\u2_Display/n5506 [29],\u2_Display/n5506 [27]}),
    .fco(\u2_Display/add167/c31 ),
    .fx({\u2_Display/n5506 [30],\u2_Display/n5506 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u31_al_u4428  (
    .a({open_n57648,\u2_Display/n5472 }),
    .c(2'b00),
    .d({open_n57653,1'b1}),
    .fci(\u2_Display/add167/c31 ),
    .f({open_n57670,\u2_Display/n5506 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u3_al_u4421  (
    .a({\u2_Display/n5498 ,\u2_Display/n5500 }),
    .b({\u2_Display/n5497 ,\u2_Display/n5499 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add167/c3 ),
    .f({\u2_Display/n5506 [5],\u2_Display/n5506 [3]}),
    .fco(\u2_Display/add167/c7 ),
    .fx({\u2_Display/n5506 [6],\u2_Display/n5506 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u7_al_u4422  (
    .a({\u2_Display/n5494 ,\u2_Display/n5496 }),
    .b({\u2_Display/n5493 ,\u2_Display/n5495 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add167/c7 ),
    .f({\u2_Display/n5506 [9],\u2_Display/n5506 [7]}),
    .fco(\u2_Display/add167/c11 ),
    .fx({\u2_Display/n5506 [10],\u2_Display/n5506 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/ucin_al_u4420  (
    .a({\u2_Display/n5502 ,1'b1}),
    .b({\u2_Display/n5501 ,\u2_Display/n5503 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5506 [1],open_n57729}),
    .fco(\u2_Display/add167/c3 ),
    .fx({\u2_Display/n5506 [2],\u2_Display/n5506 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u11_al_u4432  (
    .a({\u2_Display/n5525 ,\u2_Display/n5527 }),
    .b({\u2_Display/n5524 ,\u2_Display/n5526 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add168/c11 ),
    .f({\u2_Display/n5541 [13],\u2_Display/n5541 [11]}),
    .fco(\u2_Display/add168/c15 ),
    .fx({\u2_Display/n5541 [14],\u2_Display/n5541 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u15_al_u4433  (
    .a({\u2_Display/n5521 ,\u2_Display/n5523 }),
    .b({\u2_Display/n5520 ,\u2_Display/n5522 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add168/c15 ),
    .f({\u2_Display/n5541 [17],\u2_Display/n5541 [15]}),
    .fco(\u2_Display/add168/c19 ),
    .fx({\u2_Display/n5541 [18],\u2_Display/n5541 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u19_al_u4434  (
    .a({\u2_Display/n5517 ,\u2_Display/n5519 }),
    .b({\u2_Display/n5516 ,\u2_Display/n5518 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add168/c19 ),
    .f({\u2_Display/n5541 [21],\u2_Display/n5541 [19]}),
    .fco(\u2_Display/add168/c23 ),
    .fx({\u2_Display/n5541 [22],\u2_Display/n5541 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u23_al_u4435  (
    .a({\u2_Display/n5513 ,\u2_Display/n5515 }),
    .b({\u2_Display/n5512 ,\u2_Display/n5514 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add168/c23 ),
    .f({\u2_Display/n5541 [25],\u2_Display/n5541 [23]}),
    .fco(\u2_Display/add168/c27 ),
    .fx({\u2_Display/n5541 [26],\u2_Display/n5541 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u27_al_u4436  (
    .a({\u2_Display/n5509 ,\u2_Display/n5511 }),
    .b({\u2_Display/n5508 ,\u2_Display/n5510 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add168/c27 ),
    .f({\u2_Display/n5541 [29],\u2_Display/n5541 [27]}),
    .fco(\u2_Display/add168/c31 ),
    .fx({\u2_Display/n5541 [30],\u2_Display/n5541 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u31_al_u4437  (
    .a({open_n57822,\u2_Display/n5507 }),
    .c(2'b00),
    .d({open_n57827,1'b1}),
    .fci(\u2_Display/add168/c31 ),
    .f({open_n57844,\u2_Display/n5541 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u3_al_u4430  (
    .a({\u2_Display/n5533 ,\u2_Display/n5535 }),
    .b({\u2_Display/n5532 ,\u2_Display/n5534 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add168/c3 ),
    .f({\u2_Display/n5541 [5],\u2_Display/n5541 [3]}),
    .fco(\u2_Display/add168/c7 ),
    .fx({\u2_Display/n5541 [6],\u2_Display/n5541 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u7_al_u4431  (
    .a({\u2_Display/n5529 ,\u2_Display/n5531 }),
    .b({\u2_Display/n5528 ,\u2_Display/n5530 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add168/c7 ),
    .f({\u2_Display/n5541 [9],\u2_Display/n5541 [7]}),
    .fco(\u2_Display/add168/c11 ),
    .fx({\u2_Display/n5541 [10],\u2_Display/n5541 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/ucin_al_u4429  (
    .a({\u2_Display/n5537 ,1'b1}),
    .b({\u2_Display/n5536 ,\u2_Display/n5538 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5541 [1],open_n57903}),
    .fco(\u2_Display/add168/c3 ),
    .fx({\u2_Display/n5541 [2],\u2_Display/n5541 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u11_al_u4441  (
    .a({\u2_Display/n5560 ,\u2_Display/n5562 }),
    .b({\u2_Display/n5559 ,\u2_Display/n5561 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add169/c11 ),
    .f({\u2_Display/n5576 [13],\u2_Display/n5576 [11]}),
    .fco(\u2_Display/add169/c15 ),
    .fx({\u2_Display/n5576 [14],\u2_Display/n5576 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u15_al_u4442  (
    .a({\u2_Display/n5556 ,\u2_Display/n5558 }),
    .b({\u2_Display/n5555 ,\u2_Display/n5557 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add169/c15 ),
    .f({\u2_Display/n5576 [17],\u2_Display/n5576 [15]}),
    .fco(\u2_Display/add169/c19 ),
    .fx({\u2_Display/n5576 [18],\u2_Display/n5576 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u19_al_u4443  (
    .a({\u2_Display/n5552 ,\u2_Display/n5554 }),
    .b({\u2_Display/n5551 ,\u2_Display/n5553 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add169/c19 ),
    .f({\u2_Display/n5576 [21],\u2_Display/n5576 [19]}),
    .fco(\u2_Display/add169/c23 ),
    .fx({\u2_Display/n5576 [22],\u2_Display/n5576 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u23_al_u4444  (
    .a({\u2_Display/n5548 ,\u2_Display/n5550 }),
    .b({\u2_Display/n5547 ,\u2_Display/n5549 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add169/c23 ),
    .f({\u2_Display/n5576 [25],\u2_Display/n5576 [23]}),
    .fco(\u2_Display/add169/c27 ),
    .fx({\u2_Display/n5576 [26],\u2_Display/n5576 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u27_al_u4445  (
    .a({\u2_Display/n5544 ,\u2_Display/n5546 }),
    .b({\u2_Display/n5543 ,\u2_Display/n5545 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add169/c27 ),
    .f({\u2_Display/n5576 [29],\u2_Display/n5576 [27]}),
    .fco(\u2_Display/add169/c31 ),
    .fx({\u2_Display/n5576 [30],\u2_Display/n5576 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u31_al_u4446  (
    .a({open_n57996,\u2_Display/n5542 }),
    .c(2'b00),
    .d({open_n58001,1'b1}),
    .fci(\u2_Display/add169/c31 ),
    .f({open_n58018,\u2_Display/n5576 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u3_al_u4439  (
    .a({\u2_Display/n5568 ,\u2_Display/n5570 }),
    .b({\u2_Display/n5567 ,\u2_Display/n5569 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add169/c3 ),
    .f({\u2_Display/n5576 [5],\u2_Display/n5576 [3]}),
    .fco(\u2_Display/add169/c7 ),
    .fx({\u2_Display/n5576 [6],\u2_Display/n5576 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u7_al_u4440  (
    .a({\u2_Display/n5564 ,\u2_Display/n5566 }),
    .b({\u2_Display/n5563 ,\u2_Display/n5565 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add169/c7 ),
    .f({\u2_Display/n5576 [9],\u2_Display/n5576 [7]}),
    .fco(\u2_Display/add169/c11 ),
    .fx({\u2_Display/n5576 [10],\u2_Display/n5576 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/ucin_al_u4438  (
    .a({\u2_Display/n5572 ,1'b1}),
    .b({\u2_Display/n5571 ,\u2_Display/n5573 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5576 [1],open_n58077}),
    .fco(\u2_Display/add169/c3 ),
    .fx({\u2_Display/n5576 [2],\u2_Display/n5576 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u11_al_u4450  (
    .a({\u2_Display/n5595 ,\u2_Display/n5597 }),
    .b({\u2_Display/n5594 ,\u2_Display/n5596 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add170/c11 ),
    .f({\u2_Display/n5611 [13],\u2_Display/n5611 [11]}),
    .fco(\u2_Display/add170/c15 ),
    .fx({\u2_Display/n5611 [14],\u2_Display/n5611 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u15_al_u4451  (
    .a({\u2_Display/n5591 ,\u2_Display/n5593 }),
    .b({\u2_Display/n5590 ,\u2_Display/n5592 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add170/c15 ),
    .f({\u2_Display/n5611 [17],\u2_Display/n5611 [15]}),
    .fco(\u2_Display/add170/c19 ),
    .fx({\u2_Display/n5611 [18],\u2_Display/n5611 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u19_al_u4452  (
    .a({\u2_Display/n5587 ,\u2_Display/n5589 }),
    .b({\u2_Display/n5586 ,\u2_Display/n5588 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add170/c19 ),
    .f({\u2_Display/n5611 [21],\u2_Display/n5611 [19]}),
    .fco(\u2_Display/add170/c23 ),
    .fx({\u2_Display/n5611 [22],\u2_Display/n5611 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u23_al_u4453  (
    .a({\u2_Display/n5583 ,\u2_Display/n5585 }),
    .b({\u2_Display/n5582 ,\u2_Display/n5584 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add170/c23 ),
    .f({\u2_Display/n5611 [25],\u2_Display/n5611 [23]}),
    .fco(\u2_Display/add170/c27 ),
    .fx({\u2_Display/n5611 [26],\u2_Display/n5611 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u27_al_u4454  (
    .a({\u2_Display/n5579 ,\u2_Display/n5581 }),
    .b({\u2_Display/n5578 ,\u2_Display/n5580 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add170/c27 ),
    .f({\u2_Display/n5611 [29],\u2_Display/n5611 [27]}),
    .fco(\u2_Display/add170/c31 ),
    .fx({\u2_Display/n5611 [30],\u2_Display/n5611 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u31_al_u4455  (
    .a({open_n58170,\u2_Display/n5577 }),
    .c(2'b00),
    .d({open_n58175,1'b1}),
    .fci(\u2_Display/add170/c31 ),
    .f({open_n58192,\u2_Display/n5611 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u3_al_u4448  (
    .a({\u2_Display/n5603 ,\u2_Display/n5605 }),
    .b({\u2_Display/n5602 ,\u2_Display/n5604 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add170/c3 ),
    .f({\u2_Display/n5611 [5],\u2_Display/n5611 [3]}),
    .fco(\u2_Display/add170/c7 ),
    .fx({\u2_Display/n5611 [6],\u2_Display/n5611 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u7_al_u4449  (
    .a({\u2_Display/n5599 ,\u2_Display/n5601 }),
    .b({\u2_Display/n5598 ,\u2_Display/n5600 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add170/c7 ),
    .f({\u2_Display/n5611 [9],\u2_Display/n5611 [7]}),
    .fco(\u2_Display/add170/c11 ),
    .fx({\u2_Display/n5611 [10],\u2_Display/n5611 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/ucin_al_u4447  (
    .a({\u2_Display/n5607 ,1'b1}),
    .b({\u2_Display/n5606 ,\u2_Display/n5608 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5611 [1],open_n58251}),
    .fco(\u2_Display/add170/c3 ),
    .fx({\u2_Display/n5611 [2],\u2_Display/n5611 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u11_al_u4459  (
    .a({\u2_Display/n5630 ,\u2_Display/n5632 }),
    .b({\u2_Display/n5629 ,\u2_Display/n5631 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add171/c11 ),
    .f({\u2_Display/n5646 [13],\u2_Display/n5646 [11]}),
    .fco(\u2_Display/add171/c15 ),
    .fx({\u2_Display/n5646 [14],\u2_Display/n5646 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u15_al_u4460  (
    .a({\u2_Display/n5626 ,\u2_Display/n5628 }),
    .b({\u2_Display/n5625 ,\u2_Display/n5627 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add171/c15 ),
    .f({\u2_Display/n5646 [17],\u2_Display/n5646 [15]}),
    .fco(\u2_Display/add171/c19 ),
    .fx({\u2_Display/n5646 [18],\u2_Display/n5646 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u19_al_u4461  (
    .a({\u2_Display/n5622 ,\u2_Display/n5624 }),
    .b({\u2_Display/n5621 ,\u2_Display/n5623 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add171/c19 ),
    .f({\u2_Display/n5646 [21],\u2_Display/n5646 [19]}),
    .fco(\u2_Display/add171/c23 ),
    .fx({\u2_Display/n5646 [22],\u2_Display/n5646 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u23_al_u4462  (
    .a({\u2_Display/n5618 ,\u2_Display/n5620 }),
    .b({\u2_Display/n5617 ,\u2_Display/n5619 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add171/c23 ),
    .f({\u2_Display/n5646 [25],\u2_Display/n5646 [23]}),
    .fco(\u2_Display/add171/c27 ),
    .fx({\u2_Display/n5646 [26],\u2_Display/n5646 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u27_al_u4463  (
    .a({\u2_Display/n5614 ,\u2_Display/n5616 }),
    .b({\u2_Display/n5613 ,\u2_Display/n5615 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add171/c27 ),
    .f({\u2_Display/n5646 [29],\u2_Display/n5646 [27]}),
    .fco(\u2_Display/add171/c31 ),
    .fx({\u2_Display/n5646 [30],\u2_Display/n5646 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u31_al_u4464  (
    .a({open_n58344,\u2_Display/n5612 }),
    .c(2'b00),
    .d({open_n58349,1'b1}),
    .fci(\u2_Display/add171/c31 ),
    .f({open_n58366,\u2_Display/n5646 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u3_al_u4457  (
    .a({\u2_Display/n5638 ,\u2_Display/n5640 }),
    .b({\u2_Display/n5637 ,\u2_Display/n5639 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add171/c3 ),
    .f({\u2_Display/n5646 [5],\u2_Display/n5646 [3]}),
    .fco(\u2_Display/add171/c7 ),
    .fx({\u2_Display/n5646 [6],\u2_Display/n5646 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u7_al_u4458  (
    .a({\u2_Display/n5634 ,\u2_Display/n5636 }),
    .b({\u2_Display/n5633 ,\u2_Display/n5635 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add171/c7 ),
    .f({\u2_Display/n5646 [9],\u2_Display/n5646 [7]}),
    .fco(\u2_Display/add171/c11 ),
    .fx({\u2_Display/n5646 [10],\u2_Display/n5646 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/ucin_al_u4456  (
    .a({\u2_Display/n5642 ,1'b1}),
    .b({\u2_Display/n5641 ,\u2_Display/n5643 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5646 [1],open_n58425}),
    .fco(\u2_Display/add171/c3 ),
    .fx({\u2_Display/n5646 [2],\u2_Display/n5646 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add172/ucin_al_u5049"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add172/u3_al_u5050  (
    .a({\u2_Display/n5673 ,\u2_Display/n5675 }),
    .b({\u2_Display/n5672 ,\u2_Display/n5674 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add172/c3 ),
    .f({\u2_Display/n5681 [5],\u2_Display/n5681 [3]}),
    .fco(\u2_Display/add172/c7 ),
    .fx({\u2_Display/n5681 [6],\u2_Display/n5681 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add172/ucin_al_u5049"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add172/u7_al_u5051  (
    .a({\u2_Display/n5669 ,\u2_Display/n5671 }),
    .b({open_n58446,\u2_Display/n5670 }),
    .c(2'b00),
    .d(2'b00),
    .e({open_n58449,1'b1}),
    .fci(\u2_Display/add172/c7 ),
    .f({\u2_Display/n5681 [9],\u2_Display/n5681 [7]}),
    .fx({open_n58465,\u2_Display/n5681 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add172/ucin_al_u5049"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add172/ucin_al_u5049  (
    .a({\u2_Display/n5677 ,1'b1}),
    .b({\u2_Display/n5676 ,\u2_Display/n5678 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5681 [1],open_n58485}),
    .fco(\u2_Display/add172/c3 ),
    .fx({\u2_Display/n5681 [2],\u2_Display/n5681 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u11_al_u4468  (
    .a({\u2_Display/counta [13],\u2_Display/counta [11]}),
    .b({\u2_Display/counta [14],\u2_Display/counta [12]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add18/c11 ),
    .f({\u2_Display/n419 [13],\u2_Display/n419 [11]}),
    .fco(\u2_Display/add18/c15 ),
    .fx({\u2_Display/n419 [14],\u2_Display/n419 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u15_al_u4469  (
    .a({\u2_Display/counta [17],\u2_Display/counta [15]}),
    .b({\u2_Display/counta [18],\u2_Display/counta [16]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add18/c15 ),
    .f({\u2_Display/n419 [17],\u2_Display/n419 [15]}),
    .fco(\u2_Display/add18/c19 ),
    .fx({\u2_Display/n419 [18],\u2_Display/n419 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u19_al_u4470  (
    .a({\u2_Display/counta [21],\u2_Display/counta [19]}),
    .b({\u2_Display/counta [22],\u2_Display/counta [20]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add18/c19 ),
    .f({\u2_Display/n419 [21],\u2_Display/n419 [19]}),
    .fco(\u2_Display/add18/c23 ),
    .fx({\u2_Display/n419 [22],\u2_Display/n419 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u23_al_u4471  (
    .a({\u2_Display/counta [25],\u2_Display/counta [23]}),
    .b({\u2_Display/counta [26],\u2_Display/counta [24]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add18/c23 ),
    .f({\u2_Display/n419 [25],\u2_Display/n419 [23]}),
    .fco(\u2_Display/add18/c27 ),
    .fx({\u2_Display/n419 [26],\u2_Display/n419 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u27_al_u4472  (
    .a({\u2_Display/counta [29],\u2_Display/counta [27]}),
    .b({\u2_Display/counta [30],\u2_Display/counta [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add18/c27 ),
    .f({\u2_Display/n419 [29],\u2_Display/n419 [27]}),
    .fco(\u2_Display/add18/c31 ),
    .fx({\u2_Display/n419 [30],\u2_Display/n419 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u31_al_u4473  (
    .a({open_n58578,\u2_Display/counta [31]}),
    .c(2'b00),
    .d({open_n58583,1'b0}),
    .fci(\u2_Display/add18/c31 ),
    .f({open_n58600,\u2_Display/n419 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u3_al_u4466  (
    .a({\u2_Display/counta [5],\u2_Display/counta [3]}),
    .b({\u2_Display/counta [6],\u2_Display/counta [4]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add18/c3 ),
    .f({\u2_Display/n419 [5],\u2_Display/n419 [3]}),
    .fco(\u2_Display/add18/c7 ),
    .fx({\u2_Display/n419 [6],\u2_Display/n419 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u7_al_u4467  (
    .a({\u2_Display/counta [9],\u2_Display/counta [7]}),
    .b({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add18/c7 ),
    .f({\u2_Display/n419 [9],\u2_Display/n419 [7]}),
    .fco(\u2_Display/add18/c11 ),
    .fx({\u2_Display/n419 [10],\u2_Display/n419 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/ucin_al_u4465  (
    .a({\u2_Display/counta [1],1'b1}),
    .b({\u2_Display/counta [2],\u2_Display/counta [0]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n419 [1],open_n58659}),
    .fco(\u2_Display/add18/c3 ),
    .fx({\u2_Display/n419 [2],\u2_Display/n419 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u11_al_u4477  (
    .a({\u2_Display/n438 ,\u2_Display/n440 }),
    .b({\u2_Display/n437 ,\u2_Display/n439 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add19/c11 ),
    .f({\u2_Display/n454 [13],\u2_Display/n454 [11]}),
    .fco(\u2_Display/add19/c15 ),
    .fx({\u2_Display/n454 [14],\u2_Display/n454 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u15_al_u4478  (
    .a({\u2_Display/n434 ,\u2_Display/n436 }),
    .b({\u2_Display/n433 ,\u2_Display/n435 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add19/c15 ),
    .f({\u2_Display/n454 [17],\u2_Display/n454 [15]}),
    .fco(\u2_Display/add19/c19 ),
    .fx({\u2_Display/n454 [18],\u2_Display/n454 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u19_al_u4479  (
    .a({\u2_Display/n430 ,\u2_Display/n432 }),
    .b({\u2_Display/n429 ,\u2_Display/n431 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add19/c19 ),
    .f({\u2_Display/n454 [21],\u2_Display/n454 [19]}),
    .fco(\u2_Display/add19/c23 ),
    .fx({\u2_Display/n454 [22],\u2_Display/n454 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u23_al_u4480  (
    .a({\u2_Display/n426 ,\u2_Display/n428 }),
    .b({\u2_Display/n425 ,\u2_Display/n427 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add19/c23 ),
    .f({\u2_Display/n454 [25],\u2_Display/n454 [23]}),
    .fco(\u2_Display/add19/c27 ),
    .fx({\u2_Display/n454 [26],\u2_Display/n454 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u27_al_u4481  (
    .a({\u2_Display/n422 ,\u2_Display/n424 }),
    .b({\u2_Display/n421 ,\u2_Display/n423 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add19/c27 ),
    .f({\u2_Display/n454 [29],\u2_Display/n454 [27]}),
    .fco(\u2_Display/add19/c31 ),
    .fx({\u2_Display/n454 [30],\u2_Display/n454 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u31_al_u4482  (
    .a({open_n58752,\u2_Display/n420 }),
    .c(2'b00),
    .d({open_n58757,1'b1}),
    .fci(\u2_Display/add19/c31 ),
    .f({open_n58774,\u2_Display/n454 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u3_al_u4475  (
    .a({\u2_Display/n446 ,\u2_Display/n448 }),
    .b({\u2_Display/n445 ,\u2_Display/n447 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add19/c3 ),
    .f({\u2_Display/n454 [5],\u2_Display/n454 [3]}),
    .fco(\u2_Display/add19/c7 ),
    .fx({\u2_Display/n454 [6],\u2_Display/n454 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u7_al_u4476  (
    .a({\u2_Display/n442 ,\u2_Display/n444 }),
    .b({\u2_Display/n441 ,\u2_Display/n443 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add19/c7 ),
    .f({\u2_Display/n454 [9],\u2_Display/n454 [7]}),
    .fco(\u2_Display/add19/c11 ),
    .fx({\u2_Display/n454 [10],\u2_Display/n454 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/ucin_al_u4474  (
    .a({\u2_Display/n450 ,1'b1}),
    .b({\u2_Display/n449 ,\u2_Display/n451 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n454 [1],open_n58833}),
    .fco(\u2_Display/add19/c3 ),
    .fx({\u2_Display/n454 [2],\u2_Display/n454 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u11_al_u4486  (
    .a({\u2_Display/n473 ,\u2_Display/n475 }),
    .b({\u2_Display/n472 ,\u2_Display/n474 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add20/c11 ),
    .f({\u2_Display/n489 [13],\u2_Display/n489 [11]}),
    .fco(\u2_Display/add20/c15 ),
    .fx({\u2_Display/n489 [14],\u2_Display/n489 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u15_al_u4487  (
    .a({\u2_Display/n469 ,\u2_Display/n471 }),
    .b({\u2_Display/n468 ,\u2_Display/n470 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add20/c15 ),
    .f({\u2_Display/n489 [17],\u2_Display/n489 [15]}),
    .fco(\u2_Display/add20/c19 ),
    .fx({\u2_Display/n489 [18],\u2_Display/n489 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u19_al_u4488  (
    .a({\u2_Display/n465 ,\u2_Display/n467 }),
    .b({\u2_Display/n464 ,\u2_Display/n466 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add20/c19 ),
    .f({\u2_Display/n489 [21],\u2_Display/n489 [19]}),
    .fco(\u2_Display/add20/c23 ),
    .fx({\u2_Display/n489 [22],\u2_Display/n489 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u23_al_u4489  (
    .a({\u2_Display/n461 ,\u2_Display/n463 }),
    .b({\u2_Display/n460 ,\u2_Display/n462 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b01),
    .fci(\u2_Display/add20/c23 ),
    .f({\u2_Display/n489 [25],\u2_Display/n489 [23]}),
    .fco(\u2_Display/add20/c27 ),
    .fx({\u2_Display/n489 [26],\u2_Display/n489 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u27_al_u4490  (
    .a({\u2_Display/n457 ,\u2_Display/n459 }),
    .b({\u2_Display/n456 ,\u2_Display/n458 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add20/c27 ),
    .f({\u2_Display/n489 [29],\u2_Display/n489 [27]}),
    .fco(\u2_Display/add20/c31 ),
    .fx({\u2_Display/n489 [30],\u2_Display/n489 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u31_al_u4491  (
    .a({open_n58926,\u2_Display/n455 }),
    .c(2'b00),
    .d({open_n58931,1'b1}),
    .fci(\u2_Display/add20/c31 ),
    .f({open_n58948,\u2_Display/n489 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u3_al_u4484  (
    .a({\u2_Display/n481 ,\u2_Display/n483 }),
    .b({\u2_Display/n480 ,\u2_Display/n482 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add20/c3 ),
    .f({\u2_Display/n489 [5],\u2_Display/n489 [3]}),
    .fco(\u2_Display/add20/c7 ),
    .fx({\u2_Display/n489 [6],\u2_Display/n489 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u7_al_u4485  (
    .a({\u2_Display/n477 ,\u2_Display/n479 }),
    .b({\u2_Display/n476 ,\u2_Display/n478 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add20/c7 ),
    .f({\u2_Display/n489 [9],\u2_Display/n489 [7]}),
    .fco(\u2_Display/add20/c11 ),
    .fx({\u2_Display/n489 [10],\u2_Display/n489 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/ucin_al_u4483  (
    .a({\u2_Display/n485 ,1'b1}),
    .b({\u2_Display/n484 ,\u2_Display/n486 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n489 [1],open_n59007}),
    .fco(\u2_Display/add20/c3 ),
    .fx({\u2_Display/n489 [2],\u2_Display/n489 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u11_al_u4495  (
    .a({\u2_Display/n508 ,\u2_Display/n510 }),
    .b({\u2_Display/n507 ,\u2_Display/n509 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add21/c11 ),
    .f({\u2_Display/n524 [13],\u2_Display/n524 [11]}),
    .fco(\u2_Display/add21/c15 ),
    .fx({\u2_Display/n524 [14],\u2_Display/n524 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u15_al_u4496  (
    .a({\u2_Display/n504 ,\u2_Display/n506 }),
    .b({\u2_Display/n503 ,\u2_Display/n505 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add21/c15 ),
    .f({\u2_Display/n524 [17],\u2_Display/n524 [15]}),
    .fco(\u2_Display/add21/c19 ),
    .fx({\u2_Display/n524 [18],\u2_Display/n524 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u19_al_u4497  (
    .a({\u2_Display/n500 ,\u2_Display/n502 }),
    .b({\u2_Display/n499 ,\u2_Display/n501 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add21/c19 ),
    .f({\u2_Display/n524 [21],\u2_Display/n524 [19]}),
    .fco(\u2_Display/add21/c23 ),
    .fx({\u2_Display/n524 [22],\u2_Display/n524 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u23_al_u4498  (
    .a({\u2_Display/n496 ,\u2_Display/n498 }),
    .b({\u2_Display/n495 ,\u2_Display/n497 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add21/c23 ),
    .f({\u2_Display/n524 [25],\u2_Display/n524 [23]}),
    .fco(\u2_Display/add21/c27 ),
    .fx({\u2_Display/n524 [26],\u2_Display/n524 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u27_al_u4499  (
    .a({\u2_Display/n492 ,\u2_Display/n494 }),
    .b({\u2_Display/n491 ,\u2_Display/n493 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add21/c27 ),
    .f({\u2_Display/n524 [29],\u2_Display/n524 [27]}),
    .fco(\u2_Display/add21/c31 ),
    .fx({\u2_Display/n524 [30],\u2_Display/n524 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u31_al_u4500  (
    .a({open_n59100,\u2_Display/n490 }),
    .c(2'b00),
    .d({open_n59105,1'b1}),
    .fci(\u2_Display/add21/c31 ),
    .f({open_n59122,\u2_Display/n524 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u3_al_u4493  (
    .a({\u2_Display/n516 ,\u2_Display/n518 }),
    .b({\u2_Display/n515 ,\u2_Display/n517 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add21/c3 ),
    .f({\u2_Display/n524 [5],\u2_Display/n524 [3]}),
    .fco(\u2_Display/add21/c7 ),
    .fx({\u2_Display/n524 [6],\u2_Display/n524 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u7_al_u4494  (
    .a({\u2_Display/n512 ,\u2_Display/n514 }),
    .b({\u2_Display/n511 ,\u2_Display/n513 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add21/c7 ),
    .f({\u2_Display/n524 [9],\u2_Display/n524 [7]}),
    .fco(\u2_Display/add21/c11 ),
    .fx({\u2_Display/n524 [10],\u2_Display/n524 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/ucin_al_u4492  (
    .a({\u2_Display/n520 ,1'b1}),
    .b({\u2_Display/n519 ,\u2_Display/n521 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n524 [1],open_n59181}),
    .fco(\u2_Display/add21/c3 ),
    .fx({\u2_Display/n524 [2],\u2_Display/n524 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u11_al_u4504  (
    .a({\u2_Display/n543 ,\u2_Display/n545 }),
    .b({\u2_Display/n542 ,\u2_Display/n544 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add22/c11 ),
    .f({\u2_Display/n559 [13],\u2_Display/n559 [11]}),
    .fco(\u2_Display/add22/c15 ),
    .fx({\u2_Display/n559 [14],\u2_Display/n559 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u15_al_u4505  (
    .a({\u2_Display/n539 ,\u2_Display/n541 }),
    .b({\u2_Display/n538 ,\u2_Display/n540 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add22/c15 ),
    .f({\u2_Display/n559 [17],\u2_Display/n559 [15]}),
    .fco(\u2_Display/add22/c19 ),
    .fx({\u2_Display/n559 [18],\u2_Display/n559 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u19_al_u4506  (
    .a({\u2_Display/n535 ,\u2_Display/n537 }),
    .b({\u2_Display/n534 ,\u2_Display/n536 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add22/c19 ),
    .f({\u2_Display/n559 [21],\u2_Display/n559 [19]}),
    .fco(\u2_Display/add22/c23 ),
    .fx({\u2_Display/n559 [22],\u2_Display/n559 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u23_al_u4507  (
    .a({\u2_Display/n531 ,\u2_Display/n533 }),
    .b({\u2_Display/n530 ,\u2_Display/n532 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add22/c23 ),
    .f({\u2_Display/n559 [25],\u2_Display/n559 [23]}),
    .fco(\u2_Display/add22/c27 ),
    .fx({\u2_Display/n559 [26],\u2_Display/n559 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u27_al_u4508  (
    .a({\u2_Display/n527 ,\u2_Display/n529 }),
    .b({\u2_Display/n526 ,\u2_Display/n528 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add22/c27 ),
    .f({\u2_Display/n559 [29],\u2_Display/n559 [27]}),
    .fco(\u2_Display/add22/c31 ),
    .fx({\u2_Display/n559 [30],\u2_Display/n559 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u31_al_u4509  (
    .a({open_n59274,\u2_Display/n525 }),
    .c(2'b00),
    .d({open_n59279,1'b1}),
    .fci(\u2_Display/add22/c31 ),
    .f({open_n59296,\u2_Display/n559 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u3_al_u4502  (
    .a({\u2_Display/n551 ,\u2_Display/n553 }),
    .b({\u2_Display/n550 ,\u2_Display/n552 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add22/c3 ),
    .f({\u2_Display/n559 [5],\u2_Display/n559 [3]}),
    .fco(\u2_Display/add22/c7 ),
    .fx({\u2_Display/n559 [6],\u2_Display/n559 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u7_al_u4503  (
    .a({\u2_Display/n547 ,\u2_Display/n549 }),
    .b({\u2_Display/n546 ,\u2_Display/n548 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add22/c7 ),
    .f({\u2_Display/n559 [9],\u2_Display/n559 [7]}),
    .fco(\u2_Display/add22/c11 ),
    .fx({\u2_Display/n559 [10],\u2_Display/n559 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/ucin_al_u4501  (
    .a({\u2_Display/n555 ,1'b1}),
    .b({\u2_Display/n554 ,\u2_Display/n556 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n559 [1],open_n59355}),
    .fco(\u2_Display/add22/c3 ),
    .fx({\u2_Display/n559 [2],\u2_Display/n559 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u11_al_u4513  (
    .a({\u2_Display/n578 ,\u2_Display/n580 }),
    .b({\u2_Display/n577 ,\u2_Display/n579 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add23/c11 ),
    .f({\u2_Display/n594 [13],\u2_Display/n594 [11]}),
    .fco(\u2_Display/add23/c15 ),
    .fx({\u2_Display/n594 [14],\u2_Display/n594 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u15_al_u4514  (
    .a({\u2_Display/n574 ,\u2_Display/n576 }),
    .b({\u2_Display/n573 ,\u2_Display/n575 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add23/c15 ),
    .f({\u2_Display/n594 [17],\u2_Display/n594 [15]}),
    .fco(\u2_Display/add23/c19 ),
    .fx({\u2_Display/n594 [18],\u2_Display/n594 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u19_al_u4515  (
    .a({\u2_Display/n570 ,\u2_Display/n572 }),
    .b({\u2_Display/n569 ,\u2_Display/n571 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add23/c19 ),
    .f({\u2_Display/n594 [21],\u2_Display/n594 [19]}),
    .fco(\u2_Display/add23/c23 ),
    .fx({\u2_Display/n594 [22],\u2_Display/n594 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u23_al_u4516  (
    .a({\u2_Display/n566 ,\u2_Display/n568 }),
    .b({\u2_Display/n565 ,\u2_Display/n567 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add23/c23 ),
    .f({\u2_Display/n594 [25],\u2_Display/n594 [23]}),
    .fco(\u2_Display/add23/c27 ),
    .fx({\u2_Display/n594 [26],\u2_Display/n594 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u27_al_u4517  (
    .a({\u2_Display/n562 ,\u2_Display/n564 }),
    .b({\u2_Display/n561 ,\u2_Display/n563 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add23/c27 ),
    .f({\u2_Display/n594 [29],\u2_Display/n594 [27]}),
    .fco(\u2_Display/add23/c31 ),
    .fx({\u2_Display/n594 [30],\u2_Display/n594 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u31_al_u4518  (
    .a({open_n59448,\u2_Display/n560 }),
    .c(2'b00),
    .d({open_n59453,1'b1}),
    .fci(\u2_Display/add23/c31 ),
    .f({open_n59470,\u2_Display/n594 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u3_al_u4511  (
    .a({\u2_Display/n586 ,\u2_Display/n588 }),
    .b({\u2_Display/n585 ,\u2_Display/n587 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add23/c3 ),
    .f({\u2_Display/n594 [5],\u2_Display/n594 [3]}),
    .fco(\u2_Display/add23/c7 ),
    .fx({\u2_Display/n594 [6],\u2_Display/n594 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u7_al_u4512  (
    .a({\u2_Display/n582 ,\u2_Display/n584 }),
    .b({\u2_Display/n581 ,\u2_Display/n583 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add23/c7 ),
    .f({\u2_Display/n594 [9],\u2_Display/n594 [7]}),
    .fco(\u2_Display/add23/c11 ),
    .fx({\u2_Display/n594 [10],\u2_Display/n594 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/ucin_al_u4510  (
    .a({\u2_Display/n590 ,1'b1}),
    .b({\u2_Display/n589 ,\u2_Display/n591 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n594 [1],open_n59529}),
    .fco(\u2_Display/add23/c3 ),
    .fx({\u2_Display/n594 [2],\u2_Display/n594 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u11_al_u4522  (
    .a({\u2_Display/n613 ,\u2_Display/n615 }),
    .b({\u2_Display/n612 ,\u2_Display/n614 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add24/c11 ),
    .f({\u2_Display/n629 [13],\u2_Display/n629 [11]}),
    .fco(\u2_Display/add24/c15 ),
    .fx({\u2_Display/n629 [14],\u2_Display/n629 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u15_al_u4523  (
    .a({\u2_Display/n609 ,\u2_Display/n611 }),
    .b({\u2_Display/n608 ,\u2_Display/n610 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add24/c15 ),
    .f({\u2_Display/n629 [17],\u2_Display/n629 [15]}),
    .fco(\u2_Display/add24/c19 ),
    .fx({\u2_Display/n629 [18],\u2_Display/n629 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u19_al_u4524  (
    .a({\u2_Display/n605 ,\u2_Display/n607 }),
    .b({\u2_Display/n604 ,\u2_Display/n606 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b01),
    .fci(\u2_Display/add24/c19 ),
    .f({\u2_Display/n629 [21],\u2_Display/n629 [19]}),
    .fco(\u2_Display/add24/c23 ),
    .fx({\u2_Display/n629 [22],\u2_Display/n629 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u23_al_u4525  (
    .a({\u2_Display/n601 ,\u2_Display/n603 }),
    .b({\u2_Display/n600 ,\u2_Display/n602 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add24/c23 ),
    .f({\u2_Display/n629 [25],\u2_Display/n629 [23]}),
    .fco(\u2_Display/add24/c27 ),
    .fx({\u2_Display/n629 [26],\u2_Display/n629 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u27_al_u4526  (
    .a({\u2_Display/n597 ,\u2_Display/n599 }),
    .b({\u2_Display/n596 ,\u2_Display/n598 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add24/c27 ),
    .f({\u2_Display/n629 [29],\u2_Display/n629 [27]}),
    .fco(\u2_Display/add24/c31 ),
    .fx({\u2_Display/n629 [30],\u2_Display/n629 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u31_al_u4527  (
    .a({open_n59622,\u2_Display/n595 }),
    .c(2'b00),
    .d({open_n59627,1'b1}),
    .fci(\u2_Display/add24/c31 ),
    .f({open_n59644,\u2_Display/n629 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u3_al_u4520  (
    .a({\u2_Display/n621 ,\u2_Display/n623 }),
    .b({\u2_Display/n620 ,\u2_Display/n622 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add24/c3 ),
    .f({\u2_Display/n629 [5],\u2_Display/n629 [3]}),
    .fco(\u2_Display/add24/c7 ),
    .fx({\u2_Display/n629 [6],\u2_Display/n629 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u7_al_u4521  (
    .a({\u2_Display/n617 ,\u2_Display/n619 }),
    .b({\u2_Display/n616 ,\u2_Display/n618 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add24/c7 ),
    .f({\u2_Display/n629 [9],\u2_Display/n629 [7]}),
    .fco(\u2_Display/add24/c11 ),
    .fx({\u2_Display/n629 [10],\u2_Display/n629 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/ucin_al_u4519  (
    .a({\u2_Display/n625 ,1'b1}),
    .b({\u2_Display/n624 ,\u2_Display/n626 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n629 [1],open_n59703}),
    .fco(\u2_Display/add24/c3 ),
    .fx({\u2_Display/n629 [2],\u2_Display/n629 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u11_al_u4531  (
    .a({\u2_Display/n648 ,\u2_Display/n650 }),
    .b({\u2_Display/n647 ,\u2_Display/n649 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add25/c11 ),
    .f({\u2_Display/n664 [13],\u2_Display/n664 [11]}),
    .fco(\u2_Display/add25/c15 ),
    .fx({\u2_Display/n664 [14],\u2_Display/n664 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u15_al_u4532  (
    .a({\u2_Display/n644 ,\u2_Display/n646 }),
    .b({\u2_Display/n643 ,\u2_Display/n645 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add25/c15 ),
    .f({\u2_Display/n664 [17],\u2_Display/n664 [15]}),
    .fco(\u2_Display/add25/c19 ),
    .fx({\u2_Display/n664 [18],\u2_Display/n664 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u19_al_u4533  (
    .a({\u2_Display/n640 ,\u2_Display/n642 }),
    .b({\u2_Display/n639 ,\u2_Display/n641 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add25/c19 ),
    .f({\u2_Display/n664 [21],\u2_Display/n664 [19]}),
    .fco(\u2_Display/add25/c23 ),
    .fx({\u2_Display/n664 [22],\u2_Display/n664 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u23_al_u4534  (
    .a({\u2_Display/n636 ,\u2_Display/n638 }),
    .b({\u2_Display/n635 ,\u2_Display/n637 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add25/c23 ),
    .f({\u2_Display/n664 [25],\u2_Display/n664 [23]}),
    .fco(\u2_Display/add25/c27 ),
    .fx({\u2_Display/n664 [26],\u2_Display/n664 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u27_al_u4535  (
    .a({\u2_Display/n632 ,\u2_Display/n634 }),
    .b({\u2_Display/n631 ,\u2_Display/n633 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add25/c27 ),
    .f({\u2_Display/n664 [29],\u2_Display/n664 [27]}),
    .fco(\u2_Display/add25/c31 ),
    .fx({\u2_Display/n664 [30],\u2_Display/n664 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u31_al_u4536  (
    .a({open_n59796,\u2_Display/n630 }),
    .c(2'b00),
    .d({open_n59801,1'b1}),
    .fci(\u2_Display/add25/c31 ),
    .f({open_n59818,\u2_Display/n664 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u3_al_u4529  (
    .a({\u2_Display/n656 ,\u2_Display/n658 }),
    .b({\u2_Display/n655 ,\u2_Display/n657 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add25/c3 ),
    .f({\u2_Display/n664 [5],\u2_Display/n664 [3]}),
    .fco(\u2_Display/add25/c7 ),
    .fx({\u2_Display/n664 [6],\u2_Display/n664 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u7_al_u4530  (
    .a({\u2_Display/n652 ,\u2_Display/n654 }),
    .b({\u2_Display/n651 ,\u2_Display/n653 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add25/c7 ),
    .f({\u2_Display/n664 [9],\u2_Display/n664 [7]}),
    .fco(\u2_Display/add25/c11 ),
    .fx({\u2_Display/n664 [10],\u2_Display/n664 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/ucin_al_u4528  (
    .a({\u2_Display/n660 ,1'b1}),
    .b({\u2_Display/n659 ,\u2_Display/n661 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n664 [1],open_n59877}),
    .fco(\u2_Display/add25/c3 ),
    .fx({\u2_Display/n664 [2],\u2_Display/n664 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u11_al_u4540  (
    .a({\u2_Display/n683 ,\u2_Display/n685 }),
    .b({\u2_Display/n682 ,\u2_Display/n684 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add26/c11 ),
    .f({\u2_Display/n699 [13],\u2_Display/n699 [11]}),
    .fco(\u2_Display/add26/c15 ),
    .fx({\u2_Display/n699 [14],\u2_Display/n699 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u15_al_u4541  (
    .a({\u2_Display/n679 ,\u2_Display/n681 }),
    .b({\u2_Display/n678 ,\u2_Display/n680 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add26/c15 ),
    .f({\u2_Display/n699 [17],\u2_Display/n699 [15]}),
    .fco(\u2_Display/add26/c19 ),
    .fx({\u2_Display/n699 [18],\u2_Display/n699 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u19_al_u4542  (
    .a({\u2_Display/n675 ,\u2_Display/n677 }),
    .b({\u2_Display/n674 ,\u2_Display/n676 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add26/c19 ),
    .f({\u2_Display/n699 [21],\u2_Display/n699 [19]}),
    .fco(\u2_Display/add26/c23 ),
    .fx({\u2_Display/n699 [22],\u2_Display/n699 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u23_al_u4543  (
    .a({\u2_Display/n671 ,\u2_Display/n673 }),
    .b({\u2_Display/n670 ,\u2_Display/n672 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add26/c23 ),
    .f({\u2_Display/n699 [25],\u2_Display/n699 [23]}),
    .fco(\u2_Display/add26/c27 ),
    .fx({\u2_Display/n699 [26],\u2_Display/n699 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u27_al_u4544  (
    .a({\u2_Display/n667 ,\u2_Display/n669 }),
    .b({\u2_Display/n666 ,\u2_Display/n668 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add26/c27 ),
    .f({\u2_Display/n699 [29],\u2_Display/n699 [27]}),
    .fco(\u2_Display/add26/c31 ),
    .fx({\u2_Display/n699 [30],\u2_Display/n699 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u31_al_u4545  (
    .a({open_n59970,\u2_Display/n665 }),
    .c(2'b00),
    .d({open_n59975,1'b1}),
    .fci(\u2_Display/add26/c31 ),
    .f({open_n59992,\u2_Display/n699 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u3_al_u4538  (
    .a({\u2_Display/n691 ,\u2_Display/n693 }),
    .b({\u2_Display/n690 ,\u2_Display/n692 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add26/c3 ),
    .f({\u2_Display/n699 [5],\u2_Display/n699 [3]}),
    .fco(\u2_Display/add26/c7 ),
    .fx({\u2_Display/n699 [6],\u2_Display/n699 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u7_al_u4539  (
    .a({\u2_Display/n687 ,\u2_Display/n689 }),
    .b({\u2_Display/n686 ,\u2_Display/n688 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add26/c7 ),
    .f({\u2_Display/n699 [9],\u2_Display/n699 [7]}),
    .fco(\u2_Display/add26/c11 ),
    .fx({\u2_Display/n699 [10],\u2_Display/n699 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/ucin_al_u4537  (
    .a({\u2_Display/n695 ,1'b1}),
    .b({\u2_Display/n694 ,\u2_Display/n696 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n699 [1],open_n60051}),
    .fco(\u2_Display/add26/c3 ),
    .fx({\u2_Display/n699 [2],\u2_Display/n699 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u11_al_u4549  (
    .a({\u2_Display/n718 ,\u2_Display/n720 }),
    .b({\u2_Display/n717 ,\u2_Display/n719 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add27/c11 ),
    .f({\u2_Display/n734 [13],\u2_Display/n734 [11]}),
    .fco(\u2_Display/add27/c15 ),
    .fx({\u2_Display/n734 [14],\u2_Display/n734 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u15_al_u4550  (
    .a({\u2_Display/n714 ,\u2_Display/n716 }),
    .b({\u2_Display/n713 ,\u2_Display/n715 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add27/c15 ),
    .f({\u2_Display/n734 [17],\u2_Display/n734 [15]}),
    .fco(\u2_Display/add27/c19 ),
    .fx({\u2_Display/n734 [18],\u2_Display/n734 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u19_al_u4551  (
    .a({\u2_Display/n710 ,\u2_Display/n712 }),
    .b({\u2_Display/n709 ,\u2_Display/n711 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add27/c19 ),
    .f({\u2_Display/n734 [21],\u2_Display/n734 [19]}),
    .fco(\u2_Display/add27/c23 ),
    .fx({\u2_Display/n734 [22],\u2_Display/n734 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u23_al_u4552  (
    .a({\u2_Display/n706 ,\u2_Display/n708 }),
    .b({\u2_Display/n705 ,\u2_Display/n707 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add27/c23 ),
    .f({\u2_Display/n734 [25],\u2_Display/n734 [23]}),
    .fco(\u2_Display/add27/c27 ),
    .fx({\u2_Display/n734 [26],\u2_Display/n734 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u27_al_u4553  (
    .a({\u2_Display/n702 ,\u2_Display/n704 }),
    .b({\u2_Display/n701 ,\u2_Display/n703 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add27/c27 ),
    .f({\u2_Display/n734 [29],\u2_Display/n734 [27]}),
    .fco(\u2_Display/add27/c31 ),
    .fx({\u2_Display/n734 [30],\u2_Display/n734 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u31_al_u4554  (
    .a({open_n60144,\u2_Display/n700 }),
    .c(2'b00),
    .d({open_n60149,1'b1}),
    .fci(\u2_Display/add27/c31 ),
    .f({open_n60166,\u2_Display/n734 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u3_al_u4547  (
    .a({\u2_Display/n726 ,\u2_Display/n728 }),
    .b({\u2_Display/n725 ,\u2_Display/n727 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add27/c3 ),
    .f({\u2_Display/n734 [5],\u2_Display/n734 [3]}),
    .fco(\u2_Display/add27/c7 ),
    .fx({\u2_Display/n734 [6],\u2_Display/n734 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u7_al_u4548  (
    .a({\u2_Display/n722 ,\u2_Display/n724 }),
    .b({\u2_Display/n721 ,\u2_Display/n723 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add27/c7 ),
    .f({\u2_Display/n734 [9],\u2_Display/n734 [7]}),
    .fco(\u2_Display/add27/c11 ),
    .fx({\u2_Display/n734 [10],\u2_Display/n734 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/ucin_al_u4546  (
    .a({\u2_Display/n730 ,1'b1}),
    .b({\u2_Display/n729 ,\u2_Display/n731 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n734 [1],open_n60225}),
    .fco(\u2_Display/add27/c3 ),
    .fx({\u2_Display/n734 [2],\u2_Display/n734 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u11_al_u4558  (
    .a({\u2_Display/n753 ,\u2_Display/n755 }),
    .b({\u2_Display/n752 ,\u2_Display/n754 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add28/c11 ),
    .f({\u2_Display/n769 [13],\u2_Display/n769 [11]}),
    .fco(\u2_Display/add28/c15 ),
    .fx({\u2_Display/n769 [14],\u2_Display/n769 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u15_al_u4559  (
    .a({\u2_Display/n749 ,\u2_Display/n751 }),
    .b({\u2_Display/n748 ,\u2_Display/n750 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b01),
    .fci(\u2_Display/add28/c15 ),
    .f({\u2_Display/n769 [17],\u2_Display/n769 [15]}),
    .fco(\u2_Display/add28/c19 ),
    .fx({\u2_Display/n769 [18],\u2_Display/n769 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u19_al_u4560  (
    .a({\u2_Display/n745 ,\u2_Display/n747 }),
    .b({\u2_Display/n744 ,\u2_Display/n746 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add28/c19 ),
    .f({\u2_Display/n769 [21],\u2_Display/n769 [19]}),
    .fco(\u2_Display/add28/c23 ),
    .fx({\u2_Display/n769 [22],\u2_Display/n769 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u23_al_u4561  (
    .a({\u2_Display/n741 ,\u2_Display/n743 }),
    .b({\u2_Display/n740 ,\u2_Display/n742 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add28/c23 ),
    .f({\u2_Display/n769 [25],\u2_Display/n769 [23]}),
    .fco(\u2_Display/add28/c27 ),
    .fx({\u2_Display/n769 [26],\u2_Display/n769 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u27_al_u4562  (
    .a({\u2_Display/n737 ,\u2_Display/n739 }),
    .b({\u2_Display/n736 ,\u2_Display/n738 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add28/c27 ),
    .f({\u2_Display/n769 [29],\u2_Display/n769 [27]}),
    .fco(\u2_Display/add28/c31 ),
    .fx({\u2_Display/n769 [30],\u2_Display/n769 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u31_al_u4563  (
    .a({open_n60318,\u2_Display/n735 }),
    .c(2'b00),
    .d({open_n60323,1'b1}),
    .fci(\u2_Display/add28/c31 ),
    .f({open_n60340,\u2_Display/n769 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u3_al_u4556  (
    .a({\u2_Display/n761 ,\u2_Display/n763 }),
    .b({\u2_Display/n760 ,\u2_Display/n762 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add28/c3 ),
    .f({\u2_Display/n769 [5],\u2_Display/n769 [3]}),
    .fco(\u2_Display/add28/c7 ),
    .fx({\u2_Display/n769 [6],\u2_Display/n769 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u7_al_u4557  (
    .a({\u2_Display/n757 ,\u2_Display/n759 }),
    .b({\u2_Display/n756 ,\u2_Display/n758 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add28/c7 ),
    .f({\u2_Display/n769 [9],\u2_Display/n769 [7]}),
    .fco(\u2_Display/add28/c11 ),
    .fx({\u2_Display/n769 [10],\u2_Display/n769 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/ucin_al_u4555  (
    .a({\u2_Display/n765 ,1'b1}),
    .b({\u2_Display/n764 ,\u2_Display/n766 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n769 [1],open_n60399}),
    .fco(\u2_Display/add28/c3 ),
    .fx({\u2_Display/n769 [2],\u2_Display/n769 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u11_al_u4567  (
    .a({\u2_Display/n788 ,\u2_Display/n790 }),
    .b({\u2_Display/n787 ,\u2_Display/n789 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add29/c11 ),
    .f({\u2_Display/n804 [13],\u2_Display/n804 [11]}),
    .fco(\u2_Display/add29/c15 ),
    .fx({\u2_Display/n804 [14],\u2_Display/n804 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u15_al_u4568  (
    .a({\u2_Display/n784 ,\u2_Display/n786 }),
    .b({\u2_Display/n783 ,\u2_Display/n785 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add29/c15 ),
    .f({\u2_Display/n804 [17],\u2_Display/n804 [15]}),
    .fco(\u2_Display/add29/c19 ),
    .fx({\u2_Display/n804 [18],\u2_Display/n804 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u19_al_u4569  (
    .a({\u2_Display/n780 ,\u2_Display/n782 }),
    .b({\u2_Display/n779 ,\u2_Display/n781 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add29/c19 ),
    .f({\u2_Display/n804 [21],\u2_Display/n804 [19]}),
    .fco(\u2_Display/add29/c23 ),
    .fx({\u2_Display/n804 [22],\u2_Display/n804 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u23_al_u4570  (
    .a({\u2_Display/n776 ,\u2_Display/n778 }),
    .b({\u2_Display/n775 ,\u2_Display/n777 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add29/c23 ),
    .f({\u2_Display/n804 [25],\u2_Display/n804 [23]}),
    .fco(\u2_Display/add29/c27 ),
    .fx({\u2_Display/n804 [26],\u2_Display/n804 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u27_al_u4571  (
    .a({\u2_Display/n772 ,\u2_Display/n774 }),
    .b({\u2_Display/n771 ,\u2_Display/n773 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add29/c27 ),
    .f({\u2_Display/n804 [29],\u2_Display/n804 [27]}),
    .fco(\u2_Display/add29/c31 ),
    .fx({\u2_Display/n804 [30],\u2_Display/n804 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u31_al_u4572  (
    .a({open_n60492,\u2_Display/n770 }),
    .c(2'b00),
    .d({open_n60497,1'b1}),
    .fci(\u2_Display/add29/c31 ),
    .f({open_n60514,\u2_Display/n804 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u3_al_u4565  (
    .a({\u2_Display/n796 ,\u2_Display/n798 }),
    .b({\u2_Display/n795 ,\u2_Display/n797 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add29/c3 ),
    .f({\u2_Display/n804 [5],\u2_Display/n804 [3]}),
    .fco(\u2_Display/add29/c7 ),
    .fx({\u2_Display/n804 [6],\u2_Display/n804 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u7_al_u4566  (
    .a({\u2_Display/n792 ,\u2_Display/n794 }),
    .b({\u2_Display/n791 ,\u2_Display/n793 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add29/c7 ),
    .f({\u2_Display/n804 [9],\u2_Display/n804 [7]}),
    .fco(\u2_Display/add29/c11 ),
    .fx({\u2_Display/n804 [10],\u2_Display/n804 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/ucin_al_u4564  (
    .a({\u2_Display/n800 ,1'b1}),
    .b({\u2_Display/n799 ,\u2_Display/n801 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n804 [1],open_n60573}),
    .fco(\u2_Display/add29/c3 ),
    .fx({\u2_Display/n804 [2],\u2_Display/n804 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add2_2/u0|u2_Display/add2_2/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add2_2/u0|u2_Display/add2_2/ucin  (
    .a(2'b10),
    .b({\u2_Display/i [8],open_n60576}),
    .f({\u2_Display/n43 [0],open_n60596}),
    .fco(\u2_Display/add2_2/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add2_2/u0|u2_Display/add2_2/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add2_2/u2|u2_Display/add2_2/u1  (
    .a(2'b10),
    .b(\u2_Display/i [10:9]),
    .fci(\u2_Display/add2_2/c1 ),
    .f(\u2_Display/n43 [2:1]),
    .fco(\u2_Display/add2_2/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add2_2/u0|u2_Display/add2_2/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add2_2/ucout_al_u5058  (
    .fci(\u2_Display/add2_2/c3 ),
    .f({open_n60645,\u2_Display/add2_2_co }));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u11_al_u4576  (
    .a({\u2_Display/n823 ,\u2_Display/n825 }),
    .b({\u2_Display/n822 ,\u2_Display/n824 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add30/c11 ),
    .f({\u2_Display/n839 [13],\u2_Display/n839 [11]}),
    .fco(\u2_Display/add30/c15 ),
    .fx({\u2_Display/n839 [14],\u2_Display/n839 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u15_al_u4577  (
    .a({\u2_Display/n819 ,\u2_Display/n821 }),
    .b({\u2_Display/n818 ,\u2_Display/n820 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add30/c15 ),
    .f({\u2_Display/n839 [17],\u2_Display/n839 [15]}),
    .fco(\u2_Display/add30/c19 ),
    .fx({\u2_Display/n839 [18],\u2_Display/n839 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u19_al_u4578  (
    .a({\u2_Display/n815 ,\u2_Display/n817 }),
    .b({\u2_Display/n814 ,\u2_Display/n816 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add30/c19 ),
    .f({\u2_Display/n839 [21],\u2_Display/n839 [19]}),
    .fco(\u2_Display/add30/c23 ),
    .fx({\u2_Display/n839 [22],\u2_Display/n839 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u23_al_u4579  (
    .a({\u2_Display/n811 ,\u2_Display/n813 }),
    .b({\u2_Display/n810 ,\u2_Display/n812 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add30/c23 ),
    .f({\u2_Display/n839 [25],\u2_Display/n839 [23]}),
    .fco(\u2_Display/add30/c27 ),
    .fx({\u2_Display/n839 [26],\u2_Display/n839 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u27_al_u4580  (
    .a({\u2_Display/n807 ,\u2_Display/n809 }),
    .b({\u2_Display/n806 ,\u2_Display/n808 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add30/c27 ),
    .f({\u2_Display/n839 [29],\u2_Display/n839 [27]}),
    .fco(\u2_Display/add30/c31 ),
    .fx({\u2_Display/n839 [30],\u2_Display/n839 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u31_al_u4581  (
    .a({open_n60741,\u2_Display/n805 }),
    .c(2'b00),
    .d({open_n60746,1'b1}),
    .fci(\u2_Display/add30/c31 ),
    .f({open_n60763,\u2_Display/n839 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u3_al_u4574  (
    .a({\u2_Display/n831 ,\u2_Display/n833 }),
    .b({\u2_Display/n830 ,\u2_Display/n832 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add30/c3 ),
    .f({\u2_Display/n839 [5],\u2_Display/n839 [3]}),
    .fco(\u2_Display/add30/c7 ),
    .fx({\u2_Display/n839 [6],\u2_Display/n839 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u7_al_u4575  (
    .a({\u2_Display/n827 ,\u2_Display/n829 }),
    .b({\u2_Display/n826 ,\u2_Display/n828 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add30/c7 ),
    .f({\u2_Display/n839 [9],\u2_Display/n839 [7]}),
    .fco(\u2_Display/add30/c11 ),
    .fx({\u2_Display/n839 [10],\u2_Display/n839 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/ucin_al_u4573  (
    .a({\u2_Display/n835 ,1'b1}),
    .b({\u2_Display/n834 ,\u2_Display/n836 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n839 [1],open_n60822}),
    .fco(\u2_Display/add30/c3 ),
    .fx({\u2_Display/n839 [2],\u2_Display/n839 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u11_al_u4585  (
    .a({\u2_Display/n858 ,\u2_Display/n860 }),
    .b({\u2_Display/n857 ,\u2_Display/n859 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add31/c11 ),
    .f({\u2_Display/n874 [13],\u2_Display/n874 [11]}),
    .fco(\u2_Display/add31/c15 ),
    .fx({\u2_Display/n874 [14],\u2_Display/n874 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u15_al_u4586  (
    .a({\u2_Display/n854 ,\u2_Display/n856 }),
    .b({\u2_Display/n853 ,\u2_Display/n855 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add31/c15 ),
    .f({\u2_Display/n874 [17],\u2_Display/n874 [15]}),
    .fco(\u2_Display/add31/c19 ),
    .fx({\u2_Display/n874 [18],\u2_Display/n874 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u19_al_u4587  (
    .a({\u2_Display/n850 ,\u2_Display/n852 }),
    .b({\u2_Display/n849 ,\u2_Display/n851 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add31/c19 ),
    .f({\u2_Display/n874 [21],\u2_Display/n874 [19]}),
    .fco(\u2_Display/add31/c23 ),
    .fx({\u2_Display/n874 [22],\u2_Display/n874 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u23_al_u4588  (
    .a({\u2_Display/n846 ,\u2_Display/n848 }),
    .b({\u2_Display/n845 ,\u2_Display/n847 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add31/c23 ),
    .f({\u2_Display/n874 [25],\u2_Display/n874 [23]}),
    .fco(\u2_Display/add31/c27 ),
    .fx({\u2_Display/n874 [26],\u2_Display/n874 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u27_al_u4589  (
    .a({\u2_Display/n842 ,\u2_Display/n844 }),
    .b({\u2_Display/n841 ,\u2_Display/n843 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add31/c27 ),
    .f({\u2_Display/n874 [29],\u2_Display/n874 [27]}),
    .fco(\u2_Display/add31/c31 ),
    .fx({\u2_Display/n874 [30],\u2_Display/n874 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u31_al_u4590  (
    .a({open_n60915,\u2_Display/n840 }),
    .c(2'b00),
    .d({open_n60920,1'b1}),
    .fci(\u2_Display/add31/c31 ),
    .f({open_n60937,\u2_Display/n874 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u3_al_u4583  (
    .a({\u2_Display/n866 ,\u2_Display/n868 }),
    .b({\u2_Display/n865 ,\u2_Display/n867 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add31/c3 ),
    .f({\u2_Display/n874 [5],\u2_Display/n874 [3]}),
    .fco(\u2_Display/add31/c7 ),
    .fx({\u2_Display/n874 [6],\u2_Display/n874 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u7_al_u4584  (
    .a({\u2_Display/n862 ,\u2_Display/n864 }),
    .b({\u2_Display/n861 ,\u2_Display/n863 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add31/c7 ),
    .f({\u2_Display/n874 [9],\u2_Display/n874 [7]}),
    .fco(\u2_Display/add31/c11 ),
    .fx({\u2_Display/n874 [10],\u2_Display/n874 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/ucin_al_u4582  (
    .a({\u2_Display/n870 ,1'b1}),
    .b({\u2_Display/n869 ,\u2_Display/n871 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n874 [1],open_n60996}),
    .fco(\u2_Display/add31/c3 ),
    .fx({\u2_Display/n874 [2],\u2_Display/n874 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u11_al_u4594  (
    .a({\u2_Display/n893 ,\u2_Display/n895 }),
    .b({\u2_Display/n892 ,\u2_Display/n894 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b01),
    .fci(\u2_Display/add32/c11 ),
    .f({\u2_Display/n909 [13],\u2_Display/n909 [11]}),
    .fco(\u2_Display/add32/c15 ),
    .fx({\u2_Display/n909 [14],\u2_Display/n909 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u15_al_u4595  (
    .a({\u2_Display/n889 ,\u2_Display/n891 }),
    .b({\u2_Display/n888 ,\u2_Display/n890 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add32/c15 ),
    .f({\u2_Display/n909 [17],\u2_Display/n909 [15]}),
    .fco(\u2_Display/add32/c19 ),
    .fx({\u2_Display/n909 [18],\u2_Display/n909 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u19_al_u4596  (
    .a({\u2_Display/n885 ,\u2_Display/n887 }),
    .b({\u2_Display/n884 ,\u2_Display/n886 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add32/c19 ),
    .f({\u2_Display/n909 [21],\u2_Display/n909 [19]}),
    .fco(\u2_Display/add32/c23 ),
    .fx({\u2_Display/n909 [22],\u2_Display/n909 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u23_al_u4597  (
    .a({\u2_Display/n881 ,\u2_Display/n883 }),
    .b({\u2_Display/n880 ,\u2_Display/n882 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add32/c23 ),
    .f({\u2_Display/n909 [25],\u2_Display/n909 [23]}),
    .fco(\u2_Display/add32/c27 ),
    .fx({\u2_Display/n909 [26],\u2_Display/n909 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u27_al_u4598  (
    .a({\u2_Display/n877 ,\u2_Display/n879 }),
    .b({\u2_Display/n876 ,\u2_Display/n878 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add32/c27 ),
    .f({\u2_Display/n909 [29],\u2_Display/n909 [27]}),
    .fco(\u2_Display/add32/c31 ),
    .fx({\u2_Display/n909 [30],\u2_Display/n909 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u31_al_u4599  (
    .a({open_n61089,\u2_Display/n875 }),
    .c(2'b00),
    .d({open_n61094,1'b1}),
    .fci(\u2_Display/add32/c31 ),
    .f({open_n61111,\u2_Display/n909 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u3_al_u4592  (
    .a({\u2_Display/n901 ,\u2_Display/n903 }),
    .b({\u2_Display/n900 ,\u2_Display/n902 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add32/c3 ),
    .f({\u2_Display/n909 [5],\u2_Display/n909 [3]}),
    .fco(\u2_Display/add32/c7 ),
    .fx({\u2_Display/n909 [6],\u2_Display/n909 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u7_al_u4593  (
    .a({\u2_Display/n897 ,\u2_Display/n899 }),
    .b({\u2_Display/n896 ,\u2_Display/n898 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add32/c7 ),
    .f({\u2_Display/n909 [9],\u2_Display/n909 [7]}),
    .fco(\u2_Display/add32/c11 ),
    .fx({\u2_Display/n909 [10],\u2_Display/n909 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/ucin_al_u4591  (
    .a({\u2_Display/n905 ,1'b1}),
    .b({\u2_Display/n904 ,\u2_Display/n906 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n909 [1],open_n61170}),
    .fco(\u2_Display/add32/c3 ),
    .fx({\u2_Display/n909 [2],\u2_Display/n909 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u11_al_u4603  (
    .a({\u2_Display/n928 ,\u2_Display/n930 }),
    .b({\u2_Display/n927 ,\u2_Display/n929 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add33/c11 ),
    .f({\u2_Display/n944 [13],\u2_Display/n944 [11]}),
    .fco(\u2_Display/add33/c15 ),
    .fx({\u2_Display/n944 [14],\u2_Display/n944 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u15_al_u4604  (
    .a({\u2_Display/n924 ,\u2_Display/n926 }),
    .b({\u2_Display/n923 ,\u2_Display/n925 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add33/c15 ),
    .f({\u2_Display/n944 [17],\u2_Display/n944 [15]}),
    .fco(\u2_Display/add33/c19 ),
    .fx({\u2_Display/n944 [18],\u2_Display/n944 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u19_al_u4605  (
    .a({\u2_Display/n920 ,\u2_Display/n922 }),
    .b({\u2_Display/n919 ,\u2_Display/n921 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add33/c19 ),
    .f({\u2_Display/n944 [21],\u2_Display/n944 [19]}),
    .fco(\u2_Display/add33/c23 ),
    .fx({\u2_Display/n944 [22],\u2_Display/n944 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u23_al_u4606  (
    .a({\u2_Display/n916 ,\u2_Display/n918 }),
    .b({\u2_Display/n915 ,\u2_Display/n917 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add33/c23 ),
    .f({\u2_Display/n944 [25],\u2_Display/n944 [23]}),
    .fco(\u2_Display/add33/c27 ),
    .fx({\u2_Display/n944 [26],\u2_Display/n944 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u27_al_u4607  (
    .a({\u2_Display/n912 ,\u2_Display/n914 }),
    .b({\u2_Display/n911 ,\u2_Display/n913 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add33/c27 ),
    .f({\u2_Display/n944 [29],\u2_Display/n944 [27]}),
    .fco(\u2_Display/add33/c31 ),
    .fx({\u2_Display/n944 [30],\u2_Display/n944 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u31_al_u4608  (
    .a({open_n61263,\u2_Display/n910 }),
    .c(2'b00),
    .d({open_n61268,1'b1}),
    .fci(\u2_Display/add33/c31 ),
    .f({open_n61285,\u2_Display/n944 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u3_al_u4601  (
    .a({\u2_Display/n936 ,\u2_Display/n938 }),
    .b({\u2_Display/n935 ,\u2_Display/n937 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add33/c3 ),
    .f({\u2_Display/n944 [5],\u2_Display/n944 [3]}),
    .fco(\u2_Display/add33/c7 ),
    .fx({\u2_Display/n944 [6],\u2_Display/n944 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u7_al_u4602  (
    .a({\u2_Display/n932 ,\u2_Display/n934 }),
    .b({\u2_Display/n931 ,\u2_Display/n933 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add33/c7 ),
    .f({\u2_Display/n944 [9],\u2_Display/n944 [7]}),
    .fco(\u2_Display/add33/c11 ),
    .fx({\u2_Display/n944 [10],\u2_Display/n944 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/ucin_al_u4600  (
    .a({\u2_Display/n940 ,1'b1}),
    .b({\u2_Display/n939 ,\u2_Display/n941 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n944 [1],open_n61344}),
    .fco(\u2_Display/add33/c3 ),
    .fx({\u2_Display/n944 [2],\u2_Display/n944 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u11_al_u4612  (
    .a({\u2_Display/n963 ,\u2_Display/n965 }),
    .b({\u2_Display/n962 ,\u2_Display/n964 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add34/c11 ),
    .f({\u2_Display/n979 [13],\u2_Display/n979 [11]}),
    .fco(\u2_Display/add34/c15 ),
    .fx({\u2_Display/n979 [14],\u2_Display/n979 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u15_al_u4613  (
    .a({\u2_Display/n959 ,\u2_Display/n961 }),
    .b({\u2_Display/n958 ,\u2_Display/n960 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add34/c15 ),
    .f({\u2_Display/n979 [17],\u2_Display/n979 [15]}),
    .fco(\u2_Display/add34/c19 ),
    .fx({\u2_Display/n979 [18],\u2_Display/n979 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u19_al_u4614  (
    .a({\u2_Display/n955 ,\u2_Display/n957 }),
    .b({\u2_Display/n954 ,\u2_Display/n956 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add34/c19 ),
    .f({\u2_Display/n979 [21],\u2_Display/n979 [19]}),
    .fco(\u2_Display/add34/c23 ),
    .fx({\u2_Display/n979 [22],\u2_Display/n979 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u23_al_u4615  (
    .a({\u2_Display/n951 ,\u2_Display/n953 }),
    .b({\u2_Display/n950 ,\u2_Display/n952 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add34/c23 ),
    .f({\u2_Display/n979 [25],\u2_Display/n979 [23]}),
    .fco(\u2_Display/add34/c27 ),
    .fx({\u2_Display/n979 [26],\u2_Display/n979 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u27_al_u4616  (
    .a({\u2_Display/n947 ,\u2_Display/n949 }),
    .b({\u2_Display/n946 ,\u2_Display/n948 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add34/c27 ),
    .f({\u2_Display/n979 [29],\u2_Display/n979 [27]}),
    .fco(\u2_Display/add34/c31 ),
    .fx({\u2_Display/n979 [30],\u2_Display/n979 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u31_al_u4617  (
    .a({open_n61437,\u2_Display/n945 }),
    .c(2'b00),
    .d({open_n61442,1'b1}),
    .fci(\u2_Display/add34/c31 ),
    .f({open_n61459,\u2_Display/n979 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u3_al_u4610  (
    .a({\u2_Display/n971 ,\u2_Display/n973 }),
    .b({\u2_Display/n970 ,\u2_Display/n972 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add34/c3 ),
    .f({\u2_Display/n979 [5],\u2_Display/n979 [3]}),
    .fco(\u2_Display/add34/c7 ),
    .fx({\u2_Display/n979 [6],\u2_Display/n979 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u7_al_u4611  (
    .a({\u2_Display/n967 ,\u2_Display/n969 }),
    .b({\u2_Display/n966 ,\u2_Display/n968 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add34/c7 ),
    .f({\u2_Display/n979 [9],\u2_Display/n979 [7]}),
    .fco(\u2_Display/add34/c11 ),
    .fx({\u2_Display/n979 [10],\u2_Display/n979 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/ucin_al_u4609  (
    .a({\u2_Display/n975 ,1'b1}),
    .b({\u2_Display/n974 ,\u2_Display/n976 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n979 [1],open_n61518}),
    .fco(\u2_Display/add34/c3 ),
    .fx({\u2_Display/n979 [2],\u2_Display/n979 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u11_al_u4621  (
    .a({\u2_Display/n998 ,\u2_Display/n1000 }),
    .b({\u2_Display/n997 ,\u2_Display/n999 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add35/c11 ),
    .f({\u2_Display/n1014 [13],\u2_Display/n1014 [11]}),
    .fco(\u2_Display/add35/c15 ),
    .fx({\u2_Display/n1014 [14],\u2_Display/n1014 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u15_al_u4622  (
    .a({\u2_Display/n994 ,\u2_Display/n996 }),
    .b({\u2_Display/n993 ,\u2_Display/n995 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add35/c15 ),
    .f({\u2_Display/n1014 [17],\u2_Display/n1014 [15]}),
    .fco(\u2_Display/add35/c19 ),
    .fx({\u2_Display/n1014 [18],\u2_Display/n1014 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u19_al_u4623  (
    .a({\u2_Display/n990 ,\u2_Display/n992 }),
    .b({\u2_Display/n989 ,\u2_Display/n991 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add35/c19 ),
    .f({\u2_Display/n1014 [21],\u2_Display/n1014 [19]}),
    .fco(\u2_Display/add35/c23 ),
    .fx({\u2_Display/n1014 [22],\u2_Display/n1014 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u23_al_u4624  (
    .a({\u2_Display/n986 ,\u2_Display/n988 }),
    .b({\u2_Display/n985 ,\u2_Display/n987 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add35/c23 ),
    .f({\u2_Display/n1014 [25],\u2_Display/n1014 [23]}),
    .fco(\u2_Display/add35/c27 ),
    .fx({\u2_Display/n1014 [26],\u2_Display/n1014 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u27_al_u4625  (
    .a({\u2_Display/n982 ,\u2_Display/n984 }),
    .b({\u2_Display/n981 ,\u2_Display/n983 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add35/c27 ),
    .f({\u2_Display/n1014 [29],\u2_Display/n1014 [27]}),
    .fco(\u2_Display/add35/c31 ),
    .fx({\u2_Display/n1014 [30],\u2_Display/n1014 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u31_al_u4626  (
    .a({open_n61611,\u2_Display/n980 }),
    .c(2'b00),
    .d({open_n61616,1'b1}),
    .fci(\u2_Display/add35/c31 ),
    .f({open_n61633,\u2_Display/n1014 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u3_al_u4619  (
    .a({\u2_Display/n1006 ,\u2_Display/n1008 }),
    .b({\u2_Display/n1005 ,\u2_Display/n1007 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add35/c3 ),
    .f({\u2_Display/n1014 [5],\u2_Display/n1014 [3]}),
    .fco(\u2_Display/add35/c7 ),
    .fx({\u2_Display/n1014 [6],\u2_Display/n1014 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u7_al_u4620  (
    .a({\u2_Display/n1002 ,\u2_Display/n1004 }),
    .b({\u2_Display/n1001 ,\u2_Display/n1003 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add35/c7 ),
    .f({\u2_Display/n1014 [9],\u2_Display/n1014 [7]}),
    .fco(\u2_Display/add35/c11 ),
    .fx({\u2_Display/n1014 [10],\u2_Display/n1014 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/ucin_al_u4618  (
    .a({\u2_Display/n1010 ,1'b1}),
    .b({\u2_Display/n1009 ,\u2_Display/n1011 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1014 [1],open_n61692}),
    .fco(\u2_Display/add35/c3 ),
    .fx({\u2_Display/n1014 [2],\u2_Display/n1014 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u11_al_u4630  (
    .a({\u2_Display/n1033 ,\u2_Display/n1035 }),
    .b({\u2_Display/n1032 ,\u2_Display/n1034 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add36/c11 ),
    .f({\u2_Display/n1049 [13],\u2_Display/n1049 [11]}),
    .fco(\u2_Display/add36/c15 ),
    .fx({\u2_Display/n1049 [14],\u2_Display/n1049 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u15_al_u4631  (
    .a({\u2_Display/n1029 ,\u2_Display/n1031 }),
    .b({\u2_Display/n1028 ,\u2_Display/n1030 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add36/c15 ),
    .f({\u2_Display/n1049 [17],\u2_Display/n1049 [15]}),
    .fco(\u2_Display/add36/c19 ),
    .fx({\u2_Display/n1049 [18],\u2_Display/n1049 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u19_al_u4632  (
    .a({\u2_Display/n1025 ,\u2_Display/n1027 }),
    .b({\u2_Display/n1024 ,\u2_Display/n1026 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add36/c19 ),
    .f({\u2_Display/n1049 [21],\u2_Display/n1049 [19]}),
    .fco(\u2_Display/add36/c23 ),
    .fx({\u2_Display/n1049 [22],\u2_Display/n1049 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u23_al_u4633  (
    .a({\u2_Display/n1021 ,\u2_Display/n1023 }),
    .b({\u2_Display/n1020 ,\u2_Display/n1022 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add36/c23 ),
    .f({\u2_Display/n1049 [25],\u2_Display/n1049 [23]}),
    .fco(\u2_Display/add36/c27 ),
    .fx({\u2_Display/n1049 [26],\u2_Display/n1049 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u27_al_u4634  (
    .a({\u2_Display/n1017 ,\u2_Display/n1019 }),
    .b({\u2_Display/n1016 ,\u2_Display/n1018 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add36/c27 ),
    .f({\u2_Display/n1049 [29],\u2_Display/n1049 [27]}),
    .fco(\u2_Display/add36/c31 ),
    .fx({\u2_Display/n1049 [30],\u2_Display/n1049 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u31_al_u4635  (
    .a({open_n61785,\u2_Display/n1015 }),
    .c(2'b00),
    .d({open_n61790,1'b1}),
    .fci(\u2_Display/add36/c31 ),
    .f({open_n61807,\u2_Display/n1049 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u3_al_u4628  (
    .a({\u2_Display/n1041 ,\u2_Display/n1043 }),
    .b({\u2_Display/n1040 ,\u2_Display/n1042 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add36/c3 ),
    .f({\u2_Display/n1049 [5],\u2_Display/n1049 [3]}),
    .fco(\u2_Display/add36/c7 ),
    .fx({\u2_Display/n1049 [6],\u2_Display/n1049 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u7_al_u4629  (
    .a({\u2_Display/n1037 ,\u2_Display/n1039 }),
    .b({\u2_Display/n1036 ,\u2_Display/n1038 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b01),
    .fci(\u2_Display/add36/c7 ),
    .f({\u2_Display/n1049 [9],\u2_Display/n1049 [7]}),
    .fco(\u2_Display/add36/c11 ),
    .fx({\u2_Display/n1049 [10],\u2_Display/n1049 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/ucin_al_u4627  (
    .a({\u2_Display/n1045 ,1'b1}),
    .b({\u2_Display/n1044 ,\u2_Display/n1046 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1049 [1],open_n61866}),
    .fco(\u2_Display/add36/c3 ),
    .fx({\u2_Display/n1049 [2],\u2_Display/n1049 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u11_al_u4639  (
    .a({\u2_Display/n1068 ,\u2_Display/n1070 }),
    .b({\u2_Display/n1067 ,\u2_Display/n1069 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add37/c11 ),
    .f({\u2_Display/n1084 [13],\u2_Display/n1084 [11]}),
    .fco(\u2_Display/add37/c15 ),
    .fx({\u2_Display/n1084 [14],\u2_Display/n1084 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u15_al_u4640  (
    .a({\u2_Display/n1064 ,\u2_Display/n1066 }),
    .b({\u2_Display/n1063 ,\u2_Display/n1065 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add37/c15 ),
    .f({\u2_Display/n1084 [17],\u2_Display/n1084 [15]}),
    .fco(\u2_Display/add37/c19 ),
    .fx({\u2_Display/n1084 [18],\u2_Display/n1084 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u19_al_u4641  (
    .a({\u2_Display/n1060 ,\u2_Display/n1062 }),
    .b({\u2_Display/n1059 ,\u2_Display/n1061 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add37/c19 ),
    .f({\u2_Display/n1084 [21],\u2_Display/n1084 [19]}),
    .fco(\u2_Display/add37/c23 ),
    .fx({\u2_Display/n1084 [22],\u2_Display/n1084 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u23_al_u4642  (
    .a({\u2_Display/n1056 ,\u2_Display/n1058 }),
    .b({\u2_Display/n1055 ,\u2_Display/n1057 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add37/c23 ),
    .f({\u2_Display/n1084 [25],\u2_Display/n1084 [23]}),
    .fco(\u2_Display/add37/c27 ),
    .fx({\u2_Display/n1084 [26],\u2_Display/n1084 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u27_al_u4643  (
    .a({\u2_Display/n1052 ,\u2_Display/n1054 }),
    .b({\u2_Display/n1051 ,\u2_Display/n1053 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add37/c27 ),
    .f({\u2_Display/n1084 [29],\u2_Display/n1084 [27]}),
    .fco(\u2_Display/add37/c31 ),
    .fx({\u2_Display/n1084 [30],\u2_Display/n1084 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u31_al_u4644  (
    .a({open_n61959,\u2_Display/n1050 }),
    .c(2'b00),
    .d({open_n61964,1'b1}),
    .fci(\u2_Display/add37/c31 ),
    .f({open_n61981,\u2_Display/n1084 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u3_al_u4637  (
    .a({\u2_Display/n1076 ,\u2_Display/n1078 }),
    .b({\u2_Display/n1075 ,\u2_Display/n1077 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add37/c3 ),
    .f({\u2_Display/n1084 [5],\u2_Display/n1084 [3]}),
    .fco(\u2_Display/add37/c7 ),
    .fx({\u2_Display/n1084 [6],\u2_Display/n1084 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u7_al_u4638  (
    .a({\u2_Display/n1072 ,\u2_Display/n1074 }),
    .b({\u2_Display/n1071 ,\u2_Display/n1073 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add37/c7 ),
    .f({\u2_Display/n1084 [9],\u2_Display/n1084 [7]}),
    .fco(\u2_Display/add37/c11 ),
    .fx({\u2_Display/n1084 [10],\u2_Display/n1084 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/ucin_al_u4636  (
    .a({\u2_Display/n1080 ,1'b1}),
    .b({\u2_Display/n1079 ,\u2_Display/n1081 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1084 [1],open_n62040}),
    .fco(\u2_Display/add37/c3 ),
    .fx({\u2_Display/n1084 [2],\u2_Display/n1084 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u11_al_u4648  (
    .a({\u2_Display/n1103 ,\u2_Display/n1105 }),
    .b({\u2_Display/n1102 ,\u2_Display/n1104 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add38/c11 ),
    .f({\u2_Display/n1119 [13],\u2_Display/n1119 [11]}),
    .fco(\u2_Display/add38/c15 ),
    .fx({\u2_Display/n1119 [14],\u2_Display/n1119 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u15_al_u4649  (
    .a({\u2_Display/n1099 ,\u2_Display/n1101 }),
    .b({\u2_Display/n1098 ,\u2_Display/n1100 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add38/c15 ),
    .f({\u2_Display/n1119 [17],\u2_Display/n1119 [15]}),
    .fco(\u2_Display/add38/c19 ),
    .fx({\u2_Display/n1119 [18],\u2_Display/n1119 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u19_al_u4650  (
    .a({\u2_Display/n1095 ,\u2_Display/n1097 }),
    .b({\u2_Display/n1094 ,\u2_Display/n1096 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add38/c19 ),
    .f({\u2_Display/n1119 [21],\u2_Display/n1119 [19]}),
    .fco(\u2_Display/add38/c23 ),
    .fx({\u2_Display/n1119 [22],\u2_Display/n1119 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u23_al_u4651  (
    .a({\u2_Display/n1091 ,\u2_Display/n1093 }),
    .b({\u2_Display/n1090 ,\u2_Display/n1092 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add38/c23 ),
    .f({\u2_Display/n1119 [25],\u2_Display/n1119 [23]}),
    .fco(\u2_Display/add38/c27 ),
    .fx({\u2_Display/n1119 [26],\u2_Display/n1119 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u27_al_u4652  (
    .a({\u2_Display/n1087 ,\u2_Display/n1089 }),
    .b({\u2_Display/n1086 ,\u2_Display/n1088 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add38/c27 ),
    .f({\u2_Display/n1119 [29],\u2_Display/n1119 [27]}),
    .fco(\u2_Display/add38/c31 ),
    .fx({\u2_Display/n1119 [30],\u2_Display/n1119 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u31_al_u4653  (
    .a({open_n62133,\u2_Display/n1085 }),
    .c(2'b00),
    .d({open_n62138,1'b1}),
    .fci(\u2_Display/add38/c31 ),
    .f({open_n62155,\u2_Display/n1119 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u3_al_u4646  (
    .a({\u2_Display/n1111 ,\u2_Display/n1113 }),
    .b({\u2_Display/n1110 ,\u2_Display/n1112 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add38/c3 ),
    .f({\u2_Display/n1119 [5],\u2_Display/n1119 [3]}),
    .fco(\u2_Display/add38/c7 ),
    .fx({\u2_Display/n1119 [6],\u2_Display/n1119 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u7_al_u4647  (
    .a({\u2_Display/n1107 ,\u2_Display/n1109 }),
    .b({\u2_Display/n1106 ,\u2_Display/n1108 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add38/c7 ),
    .f({\u2_Display/n1119 [9],\u2_Display/n1119 [7]}),
    .fco(\u2_Display/add38/c11 ),
    .fx({\u2_Display/n1119 [10],\u2_Display/n1119 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/ucin_al_u4645  (
    .a({\u2_Display/n1115 ,1'b1}),
    .b({\u2_Display/n1114 ,\u2_Display/n1116 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1119 [1],open_n62214}),
    .fco(\u2_Display/add38/c3 ),
    .fx({\u2_Display/n1119 [2],\u2_Display/n1119 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u11_al_u4657  (
    .a({\u2_Display/n1138 ,\u2_Display/n1140 }),
    .b({\u2_Display/n1137 ,\u2_Display/n1139 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add39/c11 ),
    .f({\u2_Display/n1154 [13],\u2_Display/n1154 [11]}),
    .fco(\u2_Display/add39/c15 ),
    .fx({\u2_Display/n1154 [14],\u2_Display/n1154 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u15_al_u4658  (
    .a({\u2_Display/n1134 ,\u2_Display/n1136 }),
    .b({\u2_Display/n1133 ,\u2_Display/n1135 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add39/c15 ),
    .f({\u2_Display/n1154 [17],\u2_Display/n1154 [15]}),
    .fco(\u2_Display/add39/c19 ),
    .fx({\u2_Display/n1154 [18],\u2_Display/n1154 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u19_al_u4659  (
    .a({\u2_Display/n1130 ,\u2_Display/n1132 }),
    .b({\u2_Display/n1129 ,\u2_Display/n1131 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add39/c19 ),
    .f({\u2_Display/n1154 [21],\u2_Display/n1154 [19]}),
    .fco(\u2_Display/add39/c23 ),
    .fx({\u2_Display/n1154 [22],\u2_Display/n1154 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u23_al_u4660  (
    .a({\u2_Display/n1126 ,\u2_Display/n1128 }),
    .b({\u2_Display/n1125 ,\u2_Display/n1127 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add39/c23 ),
    .f({\u2_Display/n1154 [25],\u2_Display/n1154 [23]}),
    .fco(\u2_Display/add39/c27 ),
    .fx({\u2_Display/n1154 [26],\u2_Display/n1154 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u27_al_u4661  (
    .a({\u2_Display/n1122 ,\u2_Display/n1124 }),
    .b({\u2_Display/n1121 ,\u2_Display/n1123 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add39/c27 ),
    .f({\u2_Display/n1154 [29],\u2_Display/n1154 [27]}),
    .fco(\u2_Display/add39/c31 ),
    .fx({\u2_Display/n1154 [30],\u2_Display/n1154 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u31_al_u4662  (
    .a({open_n62307,\u2_Display/n1120 }),
    .c(2'b00),
    .d({open_n62312,1'b1}),
    .fci(\u2_Display/add39/c31 ),
    .f({open_n62329,\u2_Display/n1154 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u3_al_u4655  (
    .a({\u2_Display/n1146 ,\u2_Display/n1148 }),
    .b({\u2_Display/n1145 ,\u2_Display/n1147 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add39/c3 ),
    .f({\u2_Display/n1154 [5],\u2_Display/n1154 [3]}),
    .fco(\u2_Display/add39/c7 ),
    .fx({\u2_Display/n1154 [6],\u2_Display/n1154 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u7_al_u4656  (
    .a({\u2_Display/n1142 ,\u2_Display/n1144 }),
    .b({\u2_Display/n1141 ,\u2_Display/n1143 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add39/c7 ),
    .f({\u2_Display/n1154 [9],\u2_Display/n1154 [7]}),
    .fco(\u2_Display/add39/c11 ),
    .fx({\u2_Display/n1154 [10],\u2_Display/n1154 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/ucin_al_u4654  (
    .a({\u2_Display/n1150 ,1'b1}),
    .b({\u2_Display/n1149 ,\u2_Display/n1151 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1154 [1],open_n62388}),
    .fco(\u2_Display/add39/c3 ),
    .fx({\u2_Display/n1154 [2],\u2_Display/n1154 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add40/ucin_al_u5052"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add40/u3_al_u5053  (
    .a({\u2_Display/n1181 ,\u2_Display/n1183 }),
    .b({\u2_Display/n1180 ,\u2_Display/n1182 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b01),
    .fci(\u2_Display/add40/c3 ),
    .f({\u2_Display/n1189 [5],\u2_Display/n1189 [3]}),
    .fco(\u2_Display/add40/c7 ),
    .fx({\u2_Display/n1189 [6],\u2_Display/n1189 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add40/ucin_al_u5052"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add40/u7_al_u5054  (
    .a({\u2_Display/n1177 ,\u2_Display/n1179 }),
    .b({open_n62409,\u2_Display/n1178 }),
    .c(2'b00),
    .d(2'b00),
    .e({open_n62412,1'b0}),
    .fci(\u2_Display/add40/c7 ),
    .f({\u2_Display/n1189 [9],\u2_Display/n1189 [7]}),
    .fx({open_n62428,\u2_Display/n1189 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add40/ucin_al_u5052"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add40/ucin_al_u5052  (
    .a({\u2_Display/n1185 ,1'b1}),
    .b({\u2_Display/n1184 ,\u2_Display/n1186 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1189 [1],open_n62448}),
    .fco(\u2_Display/add40/c3 ),
    .fx({\u2_Display/n1189 [2],\u2_Display/n1189 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add4_2/u0|u2_Display/add4_2/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add4_2/u0|u2_Display/add4_2/ucin  (
    .a(2'b10),
    .b({\u2_Display/i [7],open_n62451}),
    .f({\u2_Display/n94 [0],open_n62471}),
    .fco(\u2_Display/add4_2/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add4_2/u0|u2_Display/add4_2/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add4_2/u2|u2_Display/add4_2/u1  (
    .a(2'b10),
    .b(\u2_Display/i [9:8]),
    .fci(\u2_Display/add4_2/c1 ),
    .f(\u2_Display/n94 [2:1]),
    .fco(\u2_Display/add4_2/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add4_2/u0|u2_Display/add4_2/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add4_2/ucout|u2_Display/add4_2/u3  (
    .a({open_n62498,1'b0}),
    .b({open_n62499,\u2_Display/i [10]}),
    .fci(\u2_Display/add4_2/c3 ),
    .f({\u2_Display/add4_2_co ,\u2_Display/n94 [3]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u11_al_u4666  (
    .a({\u2_Display/counta [13],\u2_Display/counta [11]}),
    .b({\u2_Display/counta [14],\u2_Display/counta [12]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add51/c11 ),
    .f({\u2_Display/n1542 [13],\u2_Display/n1542 [11]}),
    .fco(\u2_Display/add51/c15 ),
    .fx({\u2_Display/n1542 [14],\u2_Display/n1542 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u15_al_u4667  (
    .a({\u2_Display/counta [17],\u2_Display/counta [15]}),
    .b({\u2_Display/counta [18],\u2_Display/counta [16]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add51/c15 ),
    .f({\u2_Display/n1542 [17],\u2_Display/n1542 [15]}),
    .fco(\u2_Display/add51/c19 ),
    .fx({\u2_Display/n1542 [18],\u2_Display/n1542 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u19_al_u4668  (
    .a({\u2_Display/counta [21],\u2_Display/counta [19]}),
    .b({\u2_Display/counta [22],\u2_Display/counta [20]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add51/c19 ),
    .f({\u2_Display/n1542 [21],\u2_Display/n1542 [19]}),
    .fco(\u2_Display/add51/c23 ),
    .fx({\u2_Display/n1542 [22],\u2_Display/n1542 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u23_al_u4669  (
    .a({\u2_Display/counta [25],\u2_Display/counta [23]}),
    .b({\u2_Display/counta [26],\u2_Display/counta [24]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add51/c23 ),
    .f({\u2_Display/n1542 [25],\u2_Display/n1542 [23]}),
    .fco(\u2_Display/add51/c27 ),
    .fx({\u2_Display/n1542 [26],\u2_Display/n1542 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u27_al_u4670  (
    .a({\u2_Display/counta [29],\u2_Display/counta [27]}),
    .b({\u2_Display/counta [30],\u2_Display/counta [28]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add51/c27 ),
    .f({\u2_Display/n1542 [29],\u2_Display/n1542 [27]}),
    .fco(\u2_Display/add51/c31 ),
    .fx({\u2_Display/n1542 [30],\u2_Display/n1542 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u31_al_u4671  (
    .a({open_n62613,\u2_Display/counta [31]}),
    .c(2'b00),
    .d({open_n62618,1'b0}),
    .fci(\u2_Display/add51/c31 ),
    .f({open_n62635,\u2_Display/n1542 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u3_al_u4664  (
    .a({\u2_Display/counta [5],\u2_Display/counta [3]}),
    .b({\u2_Display/counta [6],\u2_Display/counta [4]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add51/c3 ),
    .f({\u2_Display/n1542 [5],\u2_Display/n1542 [3]}),
    .fco(\u2_Display/add51/c7 ),
    .fx({\u2_Display/n1542 [6],\u2_Display/n1542 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u7_al_u4665  (
    .a({\u2_Display/counta [9],\u2_Display/counta [7]}),
    .b({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add51/c7 ),
    .f({\u2_Display/n1542 [9],\u2_Display/n1542 [7]}),
    .fco(\u2_Display/add51/c11 ),
    .fx({\u2_Display/n1542 [10],\u2_Display/n1542 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/ucin_al_u4663  (
    .a({\u2_Display/counta [1],1'b1}),
    .b({\u2_Display/counta [2],\u2_Display/counta [0]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1542 [1],open_n62694}),
    .fco(\u2_Display/add51/c3 ),
    .fx({\u2_Display/n1542 [2],\u2_Display/n1542 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u11_al_u4675  (
    .a({\u2_Display/n1561 ,\u2_Display/n1563 }),
    .b({\u2_Display/n1560 ,\u2_Display/n1562 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add52/c11 ),
    .f({\u2_Display/n1577 [13],\u2_Display/n1577 [11]}),
    .fco(\u2_Display/add52/c15 ),
    .fx({\u2_Display/n1577 [14],\u2_Display/n1577 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u15_al_u4676  (
    .a({\u2_Display/n1557 ,\u2_Display/n1559 }),
    .b({\u2_Display/n1556 ,\u2_Display/n1558 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add52/c15 ),
    .f({\u2_Display/n1577 [17],\u2_Display/n1577 [15]}),
    .fco(\u2_Display/add52/c19 ),
    .fx({\u2_Display/n1577 [18],\u2_Display/n1577 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u19_al_u4677  (
    .a({\u2_Display/n1553 ,\u2_Display/n1555 }),
    .b({\u2_Display/n1552 ,\u2_Display/n1554 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add52/c19 ),
    .f({\u2_Display/n1577 [21],\u2_Display/n1577 [19]}),
    .fco(\u2_Display/add52/c23 ),
    .fx({\u2_Display/n1577 [22],\u2_Display/n1577 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u23_al_u4678  (
    .a({\u2_Display/n1549 ,\u2_Display/n1551 }),
    .b({\u2_Display/n1548 ,\u2_Display/n1550 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add52/c23 ),
    .f({\u2_Display/n1577 [25],\u2_Display/n1577 [23]}),
    .fco(\u2_Display/add52/c27 ),
    .fx({\u2_Display/n1577 [26],\u2_Display/n1577 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u27_al_u4679  (
    .a({\u2_Display/n1545 ,\u2_Display/n1547 }),
    .b({\u2_Display/n1544 ,\u2_Display/n1546 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add52/c27 ),
    .f({\u2_Display/n1577 [29],\u2_Display/n1577 [27]}),
    .fco(\u2_Display/add52/c31 ),
    .fx({\u2_Display/n1577 [30],\u2_Display/n1577 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u31_al_u4680  (
    .a({open_n62787,\u2_Display/n1543 }),
    .c(2'b00),
    .d({open_n62792,1'b1}),
    .fci(\u2_Display/add52/c31 ),
    .f({open_n62809,\u2_Display/n1577 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u3_al_u4673  (
    .a({\u2_Display/n1569 ,\u2_Display/n1571 }),
    .b({\u2_Display/n1568 ,\u2_Display/n1570 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add52/c3 ),
    .f({\u2_Display/n1577 [5],\u2_Display/n1577 [3]}),
    .fco(\u2_Display/add52/c7 ),
    .fx({\u2_Display/n1577 [6],\u2_Display/n1577 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u7_al_u4674  (
    .a({\u2_Display/n1565 ,\u2_Display/n1567 }),
    .b({\u2_Display/n1564 ,\u2_Display/n1566 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add52/c7 ),
    .f({\u2_Display/n1577 [9],\u2_Display/n1577 [7]}),
    .fco(\u2_Display/add52/c11 ),
    .fx({\u2_Display/n1577 [10],\u2_Display/n1577 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/ucin_al_u4672  (
    .a({\u2_Display/n1573 ,1'b1}),
    .b({\u2_Display/n1572 ,\u2_Display/n1574 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1577 [1],open_n62868}),
    .fco(\u2_Display/add52/c3 ),
    .fx({\u2_Display/n1577 [2],\u2_Display/n1577 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u11_al_u4684  (
    .a({\u2_Display/n1596 ,\u2_Display/n1598 }),
    .b({\u2_Display/n1595 ,\u2_Display/n1597 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add53/c11 ),
    .f({\u2_Display/n1612 [13],\u2_Display/n1612 [11]}),
    .fco(\u2_Display/add53/c15 ),
    .fx({\u2_Display/n1612 [14],\u2_Display/n1612 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u15_al_u4685  (
    .a({\u2_Display/n1592 ,\u2_Display/n1594 }),
    .b({\u2_Display/n1591 ,\u2_Display/n1593 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add53/c15 ),
    .f({\u2_Display/n1612 [17],\u2_Display/n1612 [15]}),
    .fco(\u2_Display/add53/c19 ),
    .fx({\u2_Display/n1612 [18],\u2_Display/n1612 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u19_al_u4686  (
    .a({\u2_Display/n1588 ,\u2_Display/n1590 }),
    .b({\u2_Display/n1587 ,\u2_Display/n1589 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add53/c19 ),
    .f({\u2_Display/n1612 [21],\u2_Display/n1612 [19]}),
    .fco(\u2_Display/add53/c23 ),
    .fx({\u2_Display/n1612 [22],\u2_Display/n1612 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u23_al_u4687  (
    .a({\u2_Display/n1584 ,\u2_Display/n1586 }),
    .b({\u2_Display/n1583 ,\u2_Display/n1585 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add53/c23 ),
    .f({\u2_Display/n1612 [25],\u2_Display/n1612 [23]}),
    .fco(\u2_Display/add53/c27 ),
    .fx({\u2_Display/n1612 [26],\u2_Display/n1612 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u27_al_u4688  (
    .a({\u2_Display/n1580 ,\u2_Display/n1582 }),
    .b({\u2_Display/n1579 ,\u2_Display/n1581 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add53/c27 ),
    .f({\u2_Display/n1612 [29],\u2_Display/n1612 [27]}),
    .fco(\u2_Display/add53/c31 ),
    .fx({\u2_Display/n1612 [30],\u2_Display/n1612 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u31_al_u4689  (
    .a({open_n62961,\u2_Display/n1578 }),
    .c(2'b00),
    .d({open_n62966,1'b1}),
    .fci(\u2_Display/add53/c31 ),
    .f({open_n62983,\u2_Display/n1612 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u3_al_u4682  (
    .a({\u2_Display/n1604 ,\u2_Display/n1606 }),
    .b({\u2_Display/n1603 ,\u2_Display/n1605 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add53/c3 ),
    .f({\u2_Display/n1612 [5],\u2_Display/n1612 [3]}),
    .fco(\u2_Display/add53/c7 ),
    .fx({\u2_Display/n1612 [6],\u2_Display/n1612 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u7_al_u4683  (
    .a({\u2_Display/n1600 ,\u2_Display/n1602 }),
    .b({\u2_Display/n1599 ,\u2_Display/n1601 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add53/c7 ),
    .f({\u2_Display/n1612 [9],\u2_Display/n1612 [7]}),
    .fco(\u2_Display/add53/c11 ),
    .fx({\u2_Display/n1612 [10],\u2_Display/n1612 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/ucin_al_u4681  (
    .a({\u2_Display/n1608 ,1'b1}),
    .b({\u2_Display/n1607 ,\u2_Display/n1609 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1612 [1],open_n63042}),
    .fco(\u2_Display/add53/c3 ),
    .fx({\u2_Display/n1612 [2],\u2_Display/n1612 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u11_al_u4693  (
    .a({\u2_Display/n1631 ,\u2_Display/n1633 }),
    .b({\u2_Display/n1630 ,\u2_Display/n1632 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add54/c11 ),
    .f({\u2_Display/n1647 [13],\u2_Display/n1647 [11]}),
    .fco(\u2_Display/add54/c15 ),
    .fx({\u2_Display/n1647 [14],\u2_Display/n1647 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u15_al_u4694  (
    .a({\u2_Display/n1627 ,\u2_Display/n1629 }),
    .b({\u2_Display/n1626 ,\u2_Display/n1628 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add54/c15 ),
    .f({\u2_Display/n1647 [17],\u2_Display/n1647 [15]}),
    .fco(\u2_Display/add54/c19 ),
    .fx({\u2_Display/n1647 [18],\u2_Display/n1647 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u19_al_u4695  (
    .a({\u2_Display/n1623 ,\u2_Display/n1625 }),
    .b({\u2_Display/n1622 ,\u2_Display/n1624 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add54/c19 ),
    .f({\u2_Display/n1647 [21],\u2_Display/n1647 [19]}),
    .fco(\u2_Display/add54/c23 ),
    .fx({\u2_Display/n1647 [22],\u2_Display/n1647 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u23_al_u4696  (
    .a({\u2_Display/n1619 ,\u2_Display/n1621 }),
    .b({\u2_Display/n1618 ,\u2_Display/n1620 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add54/c23 ),
    .f({\u2_Display/n1647 [25],\u2_Display/n1647 [23]}),
    .fco(\u2_Display/add54/c27 ),
    .fx({\u2_Display/n1647 [26],\u2_Display/n1647 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u27_al_u4697  (
    .a({\u2_Display/n1615 ,\u2_Display/n1617 }),
    .b({\u2_Display/n1614 ,\u2_Display/n1616 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add54/c27 ),
    .f({\u2_Display/n1647 [29],\u2_Display/n1647 [27]}),
    .fco(\u2_Display/add54/c31 ),
    .fx({\u2_Display/n1647 [30],\u2_Display/n1647 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u31_al_u4698  (
    .a({open_n63135,\u2_Display/n1613 }),
    .c(2'b00),
    .d({open_n63140,1'b1}),
    .fci(\u2_Display/add54/c31 ),
    .f({open_n63157,\u2_Display/n1647 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u3_al_u4691  (
    .a({\u2_Display/n1639 ,\u2_Display/n1641 }),
    .b({\u2_Display/n1638 ,\u2_Display/n1640 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add54/c3 ),
    .f({\u2_Display/n1647 [5],\u2_Display/n1647 [3]}),
    .fco(\u2_Display/add54/c7 ),
    .fx({\u2_Display/n1647 [6],\u2_Display/n1647 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u7_al_u4692  (
    .a({\u2_Display/n1635 ,\u2_Display/n1637 }),
    .b({\u2_Display/n1634 ,\u2_Display/n1636 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add54/c7 ),
    .f({\u2_Display/n1647 [9],\u2_Display/n1647 [7]}),
    .fco(\u2_Display/add54/c11 ),
    .fx({\u2_Display/n1647 [10],\u2_Display/n1647 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/ucin_al_u4690  (
    .a({\u2_Display/n1643 ,1'b1}),
    .b({\u2_Display/n1642 ,\u2_Display/n1644 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1647 [1],open_n63216}),
    .fco(\u2_Display/add54/c3 ),
    .fx({\u2_Display/n1647 [2],\u2_Display/n1647 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u11_al_u4702  (
    .a({\u2_Display/n1666 ,\u2_Display/n1668 }),
    .b({\u2_Display/n1665 ,\u2_Display/n1667 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add55/c11 ),
    .f({\u2_Display/n1682 [13],\u2_Display/n1682 [11]}),
    .fco(\u2_Display/add55/c15 ),
    .fx({\u2_Display/n1682 [14],\u2_Display/n1682 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u15_al_u4703  (
    .a({\u2_Display/n1662 ,\u2_Display/n1664 }),
    .b({\u2_Display/n1661 ,\u2_Display/n1663 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add55/c15 ),
    .f({\u2_Display/n1682 [17],\u2_Display/n1682 [15]}),
    .fco(\u2_Display/add55/c19 ),
    .fx({\u2_Display/n1682 [18],\u2_Display/n1682 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u19_al_u4704  (
    .a({\u2_Display/n1658 ,\u2_Display/n1660 }),
    .b({\u2_Display/n1657 ,\u2_Display/n1659 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add55/c19 ),
    .f({\u2_Display/n1682 [21],\u2_Display/n1682 [19]}),
    .fco(\u2_Display/add55/c23 ),
    .fx({\u2_Display/n1682 [22],\u2_Display/n1682 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u23_al_u4705  (
    .a({\u2_Display/n1654 ,\u2_Display/n1656 }),
    .b({\u2_Display/n1653 ,\u2_Display/n1655 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add55/c23 ),
    .f({\u2_Display/n1682 [25],\u2_Display/n1682 [23]}),
    .fco(\u2_Display/add55/c27 ),
    .fx({\u2_Display/n1682 [26],\u2_Display/n1682 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u27_al_u4706  (
    .a({\u2_Display/n1650 ,\u2_Display/n1652 }),
    .b({\u2_Display/n1649 ,\u2_Display/n1651 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add55/c27 ),
    .f({\u2_Display/n1682 [29],\u2_Display/n1682 [27]}),
    .fco(\u2_Display/add55/c31 ),
    .fx({\u2_Display/n1682 [30],\u2_Display/n1682 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u31_al_u4707  (
    .a({open_n63309,\u2_Display/n1648 }),
    .c(2'b00),
    .d({open_n63314,1'b1}),
    .fci(\u2_Display/add55/c31 ),
    .f({open_n63331,\u2_Display/n1682 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u3_al_u4700  (
    .a({\u2_Display/n1674 ,\u2_Display/n1676 }),
    .b({\u2_Display/n1673 ,\u2_Display/n1675 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add55/c3 ),
    .f({\u2_Display/n1682 [5],\u2_Display/n1682 [3]}),
    .fco(\u2_Display/add55/c7 ),
    .fx({\u2_Display/n1682 [6],\u2_Display/n1682 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u7_al_u4701  (
    .a({\u2_Display/n1670 ,\u2_Display/n1672 }),
    .b({\u2_Display/n1669 ,\u2_Display/n1671 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add55/c7 ),
    .f({\u2_Display/n1682 [9],\u2_Display/n1682 [7]}),
    .fco(\u2_Display/add55/c11 ),
    .fx({\u2_Display/n1682 [10],\u2_Display/n1682 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/ucin_al_u4699  (
    .a({\u2_Display/n1678 ,1'b1}),
    .b({\u2_Display/n1677 ,\u2_Display/n1679 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1682 [1],open_n63390}),
    .fco(\u2_Display/add55/c3 ),
    .fx({\u2_Display/n1682 [2],\u2_Display/n1682 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u11_al_u4711  (
    .a({\u2_Display/n1701 ,\u2_Display/n1703 }),
    .b({\u2_Display/n1700 ,\u2_Display/n1702 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add56/c11 ),
    .f({\u2_Display/n1717 [13],\u2_Display/n1717 [11]}),
    .fco(\u2_Display/add56/c15 ),
    .fx({\u2_Display/n1717 [14],\u2_Display/n1717 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u15_al_u4712  (
    .a({\u2_Display/n1697 ,\u2_Display/n1699 }),
    .b({\u2_Display/n1696 ,\u2_Display/n1698 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add56/c15 ),
    .f({\u2_Display/n1717 [17],\u2_Display/n1717 [15]}),
    .fco(\u2_Display/add56/c19 ),
    .fx({\u2_Display/n1717 [18],\u2_Display/n1717 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u19_al_u4713  (
    .a({\u2_Display/n1693 ,\u2_Display/n1695 }),
    .b({\u2_Display/n1692 ,\u2_Display/n1694 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add56/c19 ),
    .f({\u2_Display/n1717 [21],\u2_Display/n1717 [19]}),
    .fco(\u2_Display/add56/c23 ),
    .fx({\u2_Display/n1717 [22],\u2_Display/n1717 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u23_al_u4714  (
    .a({\u2_Display/n1689 ,\u2_Display/n1691 }),
    .b({\u2_Display/n1688 ,\u2_Display/n1690 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add56/c23 ),
    .f({\u2_Display/n1717 [25],\u2_Display/n1717 [23]}),
    .fco(\u2_Display/add56/c27 ),
    .fx({\u2_Display/n1717 [26],\u2_Display/n1717 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u27_al_u4715  (
    .a({\u2_Display/n1685 ,\u2_Display/n1687 }),
    .b({\u2_Display/n1684 ,\u2_Display/n1686 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add56/c27 ),
    .f({\u2_Display/n1717 [29],\u2_Display/n1717 [27]}),
    .fco(\u2_Display/add56/c31 ),
    .fx({\u2_Display/n1717 [30],\u2_Display/n1717 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u31_al_u4716  (
    .a({open_n63483,\u2_Display/n1683 }),
    .c(2'b00),
    .d({open_n63488,1'b1}),
    .fci(\u2_Display/add56/c31 ),
    .f({open_n63505,\u2_Display/n1717 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u3_al_u4709  (
    .a({\u2_Display/n1709 ,\u2_Display/n1711 }),
    .b({\u2_Display/n1708 ,\u2_Display/n1710 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add56/c3 ),
    .f({\u2_Display/n1717 [5],\u2_Display/n1717 [3]}),
    .fco(\u2_Display/add56/c7 ),
    .fx({\u2_Display/n1717 [6],\u2_Display/n1717 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u7_al_u4710  (
    .a({\u2_Display/n1705 ,\u2_Display/n1707 }),
    .b({\u2_Display/n1704 ,\u2_Display/n1706 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add56/c7 ),
    .f({\u2_Display/n1717 [9],\u2_Display/n1717 [7]}),
    .fco(\u2_Display/add56/c11 ),
    .fx({\u2_Display/n1717 [10],\u2_Display/n1717 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/ucin_al_u4708  (
    .a({\u2_Display/n1713 ,1'b1}),
    .b({\u2_Display/n1712 ,\u2_Display/n1714 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1717 [1],open_n63564}),
    .fco(\u2_Display/add56/c3 ),
    .fx({\u2_Display/n1717 [2],\u2_Display/n1717 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u11_al_u4720  (
    .a({\u2_Display/n1736 ,\u2_Display/n1738 }),
    .b({\u2_Display/n1735 ,\u2_Display/n1737 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add57/c11 ),
    .f({\u2_Display/n1752 [13],\u2_Display/n1752 [11]}),
    .fco(\u2_Display/add57/c15 ),
    .fx({\u2_Display/n1752 [14],\u2_Display/n1752 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u15_al_u4721  (
    .a({\u2_Display/n1732 ,\u2_Display/n1734 }),
    .b({\u2_Display/n1731 ,\u2_Display/n1733 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add57/c15 ),
    .f({\u2_Display/n1752 [17],\u2_Display/n1752 [15]}),
    .fco(\u2_Display/add57/c19 ),
    .fx({\u2_Display/n1752 [18],\u2_Display/n1752 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u19_al_u4722  (
    .a({\u2_Display/n1728 ,\u2_Display/n1730 }),
    .b({\u2_Display/n1727 ,\u2_Display/n1729 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add57/c19 ),
    .f({\u2_Display/n1752 [21],\u2_Display/n1752 [19]}),
    .fco(\u2_Display/add57/c23 ),
    .fx({\u2_Display/n1752 [22],\u2_Display/n1752 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u23_al_u4723  (
    .a({\u2_Display/n1724 ,\u2_Display/n1726 }),
    .b({\u2_Display/n1723 ,\u2_Display/n1725 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add57/c23 ),
    .f({\u2_Display/n1752 [25],\u2_Display/n1752 [23]}),
    .fco(\u2_Display/add57/c27 ),
    .fx({\u2_Display/n1752 [26],\u2_Display/n1752 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u27_al_u4724  (
    .a({\u2_Display/n1720 ,\u2_Display/n1722 }),
    .b({\u2_Display/n1719 ,\u2_Display/n1721 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add57/c27 ),
    .f({\u2_Display/n1752 [29],\u2_Display/n1752 [27]}),
    .fco(\u2_Display/add57/c31 ),
    .fx({\u2_Display/n1752 [30],\u2_Display/n1752 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u31_al_u4725  (
    .a({open_n63657,\u2_Display/n1718 }),
    .c(2'b00),
    .d({open_n63662,1'b1}),
    .fci(\u2_Display/add57/c31 ),
    .f({open_n63679,\u2_Display/n1752 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u3_al_u4718  (
    .a({\u2_Display/n1744 ,\u2_Display/n1746 }),
    .b({\u2_Display/n1743 ,\u2_Display/n1745 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add57/c3 ),
    .f({\u2_Display/n1752 [5],\u2_Display/n1752 [3]}),
    .fco(\u2_Display/add57/c7 ),
    .fx({\u2_Display/n1752 [6],\u2_Display/n1752 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u7_al_u4719  (
    .a({\u2_Display/n1740 ,\u2_Display/n1742 }),
    .b({\u2_Display/n1739 ,\u2_Display/n1741 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add57/c7 ),
    .f({\u2_Display/n1752 [9],\u2_Display/n1752 [7]}),
    .fco(\u2_Display/add57/c11 ),
    .fx({\u2_Display/n1752 [10],\u2_Display/n1752 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/ucin_al_u4717  (
    .a({\u2_Display/n1748 ,1'b1}),
    .b({\u2_Display/n1747 ,\u2_Display/n1749 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1752 [1],open_n63738}),
    .fco(\u2_Display/add57/c3 ),
    .fx({\u2_Display/n1752 [2],\u2_Display/n1752 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u11_al_u4729  (
    .a({\u2_Display/n1771 ,\u2_Display/n1773 }),
    .b({\u2_Display/n1770 ,\u2_Display/n1772 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add58/c11 ),
    .f({\u2_Display/n1787 [13],\u2_Display/n1787 [11]}),
    .fco(\u2_Display/add58/c15 ),
    .fx({\u2_Display/n1787 [14],\u2_Display/n1787 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u15_al_u4730  (
    .a({\u2_Display/n1767 ,\u2_Display/n1769 }),
    .b({\u2_Display/n1766 ,\u2_Display/n1768 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add58/c15 ),
    .f({\u2_Display/n1787 [17],\u2_Display/n1787 [15]}),
    .fco(\u2_Display/add58/c19 ),
    .fx({\u2_Display/n1787 [18],\u2_Display/n1787 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u19_al_u4731  (
    .a({\u2_Display/n1763 ,\u2_Display/n1765 }),
    .b({\u2_Display/n1762 ,\u2_Display/n1764 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add58/c19 ),
    .f({\u2_Display/n1787 [21],\u2_Display/n1787 [19]}),
    .fco(\u2_Display/add58/c23 ),
    .fx({\u2_Display/n1787 [22],\u2_Display/n1787 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u23_al_u4732  (
    .a({\u2_Display/n1759 ,\u2_Display/n1761 }),
    .b({\u2_Display/n1758 ,\u2_Display/n1760 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add58/c23 ),
    .f({\u2_Display/n1787 [25],\u2_Display/n1787 [23]}),
    .fco(\u2_Display/add58/c27 ),
    .fx({\u2_Display/n1787 [26],\u2_Display/n1787 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u27_al_u4733  (
    .a({\u2_Display/n1755 ,\u2_Display/n1757 }),
    .b({\u2_Display/n1754 ,\u2_Display/n1756 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add58/c27 ),
    .f({\u2_Display/n1787 [29],\u2_Display/n1787 [27]}),
    .fco(\u2_Display/add58/c31 ),
    .fx({\u2_Display/n1787 [30],\u2_Display/n1787 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u31_al_u4734  (
    .a({open_n63831,\u2_Display/n1753 }),
    .c(2'b00),
    .d({open_n63836,1'b1}),
    .fci(\u2_Display/add58/c31 ),
    .f({open_n63853,\u2_Display/n1787 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u3_al_u4727  (
    .a({\u2_Display/n1779 ,\u2_Display/n1781 }),
    .b({\u2_Display/n1778 ,\u2_Display/n1780 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add58/c3 ),
    .f({\u2_Display/n1787 [5],\u2_Display/n1787 [3]}),
    .fco(\u2_Display/add58/c7 ),
    .fx({\u2_Display/n1787 [6],\u2_Display/n1787 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u7_al_u4728  (
    .a({\u2_Display/n1775 ,\u2_Display/n1777 }),
    .b({\u2_Display/n1774 ,\u2_Display/n1776 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add58/c7 ),
    .f({\u2_Display/n1787 [9],\u2_Display/n1787 [7]}),
    .fco(\u2_Display/add58/c11 ),
    .fx({\u2_Display/n1787 [10],\u2_Display/n1787 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/ucin_al_u4726  (
    .a({\u2_Display/n1783 ,1'b1}),
    .b({\u2_Display/n1782 ,\u2_Display/n1784 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1787 [1],open_n63912}),
    .fco(\u2_Display/add58/c3 ),
    .fx({\u2_Display/n1787 [2],\u2_Display/n1787 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u11_al_u4738  (
    .a({\u2_Display/n1806 ,\u2_Display/n1808 }),
    .b({\u2_Display/n1805 ,\u2_Display/n1807 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add59/c11 ),
    .f({\u2_Display/n1822 [13],\u2_Display/n1822 [11]}),
    .fco(\u2_Display/add59/c15 ),
    .fx({\u2_Display/n1822 [14],\u2_Display/n1822 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u15_al_u4739  (
    .a({\u2_Display/n1802 ,\u2_Display/n1804 }),
    .b({\u2_Display/n1801 ,\u2_Display/n1803 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add59/c15 ),
    .f({\u2_Display/n1822 [17],\u2_Display/n1822 [15]}),
    .fco(\u2_Display/add59/c19 ),
    .fx({\u2_Display/n1822 [18],\u2_Display/n1822 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u19_al_u4740  (
    .a({\u2_Display/n1798 ,\u2_Display/n1800 }),
    .b({\u2_Display/n1797 ,\u2_Display/n1799 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add59/c19 ),
    .f({\u2_Display/n1822 [21],\u2_Display/n1822 [19]}),
    .fco(\u2_Display/add59/c23 ),
    .fx({\u2_Display/n1822 [22],\u2_Display/n1822 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u23_al_u4741  (
    .a({\u2_Display/n1794 ,\u2_Display/n1796 }),
    .b({\u2_Display/n1793 ,\u2_Display/n1795 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add59/c23 ),
    .f({\u2_Display/n1822 [25],\u2_Display/n1822 [23]}),
    .fco(\u2_Display/add59/c27 ),
    .fx({\u2_Display/n1822 [26],\u2_Display/n1822 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u27_al_u4742  (
    .a({\u2_Display/n1790 ,\u2_Display/n1792 }),
    .b({\u2_Display/n1789 ,\u2_Display/n1791 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add59/c27 ),
    .f({\u2_Display/n1822 [29],\u2_Display/n1822 [27]}),
    .fco(\u2_Display/add59/c31 ),
    .fx({\u2_Display/n1822 [30],\u2_Display/n1822 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u31_al_u4743  (
    .a({open_n64005,\u2_Display/n1788 }),
    .c(2'b00),
    .d({open_n64010,1'b1}),
    .fci(\u2_Display/add59/c31 ),
    .f({open_n64027,\u2_Display/n1822 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u3_al_u4736  (
    .a({\u2_Display/n1814 ,\u2_Display/n1816 }),
    .b({\u2_Display/n1813 ,\u2_Display/n1815 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add59/c3 ),
    .f({\u2_Display/n1822 [5],\u2_Display/n1822 [3]}),
    .fco(\u2_Display/add59/c7 ),
    .fx({\u2_Display/n1822 [6],\u2_Display/n1822 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u7_al_u4737  (
    .a({\u2_Display/n1810 ,\u2_Display/n1812 }),
    .b({\u2_Display/n1809 ,\u2_Display/n1811 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add59/c7 ),
    .f({\u2_Display/n1822 [9],\u2_Display/n1822 [7]}),
    .fco(\u2_Display/add59/c11 ),
    .fx({\u2_Display/n1822 [10],\u2_Display/n1822 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/ucin_al_u4735  (
    .a({\u2_Display/n1818 ,1'b1}),
    .b({\u2_Display/n1817 ,\u2_Display/n1819 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1822 [1],open_n64086}),
    .fco(\u2_Display/add59/c3 ),
    .fx({\u2_Display/n1822 [2],\u2_Display/n1822 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u11_al_u4747  (
    .a({\u2_Display/n1841 ,\u2_Display/n1843 }),
    .b({\u2_Display/n1840 ,\u2_Display/n1842 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add60/c11 ),
    .f({\u2_Display/n1857 [13],\u2_Display/n1857 [11]}),
    .fco(\u2_Display/add60/c15 ),
    .fx({\u2_Display/n1857 [14],\u2_Display/n1857 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u15_al_u4748  (
    .a({\u2_Display/n1837 ,\u2_Display/n1839 }),
    .b({\u2_Display/n1836 ,\u2_Display/n1838 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add60/c15 ),
    .f({\u2_Display/n1857 [17],\u2_Display/n1857 [15]}),
    .fco(\u2_Display/add60/c19 ),
    .fx({\u2_Display/n1857 [18],\u2_Display/n1857 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u19_al_u4749  (
    .a({\u2_Display/n1833 ,\u2_Display/n1835 }),
    .b({\u2_Display/n1832 ,\u2_Display/n1834 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add60/c19 ),
    .f({\u2_Display/n1857 [21],\u2_Display/n1857 [19]}),
    .fco(\u2_Display/add60/c23 ),
    .fx({\u2_Display/n1857 [22],\u2_Display/n1857 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u23_al_u4750  (
    .a({\u2_Display/n1829 ,\u2_Display/n1831 }),
    .b({\u2_Display/n1828 ,\u2_Display/n1830 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add60/c23 ),
    .f({\u2_Display/n1857 [25],\u2_Display/n1857 [23]}),
    .fco(\u2_Display/add60/c27 ),
    .fx({\u2_Display/n1857 [26],\u2_Display/n1857 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u27_al_u4751  (
    .a({\u2_Display/n1825 ,\u2_Display/n1827 }),
    .b({\u2_Display/n1824 ,\u2_Display/n1826 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add60/c27 ),
    .f({\u2_Display/n1857 [29],\u2_Display/n1857 [27]}),
    .fco(\u2_Display/add60/c31 ),
    .fx({\u2_Display/n1857 [30],\u2_Display/n1857 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u31_al_u4752  (
    .a({open_n64179,\u2_Display/n1823 }),
    .c(2'b00),
    .d({open_n64184,1'b1}),
    .fci(\u2_Display/add60/c31 ),
    .f({open_n64201,\u2_Display/n1857 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u3_al_u4745  (
    .a({\u2_Display/n1849 ,\u2_Display/n1851 }),
    .b({\u2_Display/n1848 ,\u2_Display/n1850 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add60/c3 ),
    .f({\u2_Display/n1857 [5],\u2_Display/n1857 [3]}),
    .fco(\u2_Display/add60/c7 ),
    .fx({\u2_Display/n1857 [6],\u2_Display/n1857 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u7_al_u4746  (
    .a({\u2_Display/n1845 ,\u2_Display/n1847 }),
    .b({\u2_Display/n1844 ,\u2_Display/n1846 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add60/c7 ),
    .f({\u2_Display/n1857 [9],\u2_Display/n1857 [7]}),
    .fco(\u2_Display/add60/c11 ),
    .fx({\u2_Display/n1857 [10],\u2_Display/n1857 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/ucin_al_u4744  (
    .a({\u2_Display/n1853 ,1'b1}),
    .b({\u2_Display/n1852 ,\u2_Display/n1854 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1857 [1],open_n64260}),
    .fco(\u2_Display/add60/c3 ),
    .fx({\u2_Display/n1857 [2],\u2_Display/n1857 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u11_al_u4756  (
    .a({\u2_Display/n1876 ,\u2_Display/n1878 }),
    .b({\u2_Display/n1875 ,\u2_Display/n1877 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add61/c11 ),
    .f({\u2_Display/n1892 [13],\u2_Display/n1892 [11]}),
    .fco(\u2_Display/add61/c15 ),
    .fx({\u2_Display/n1892 [14],\u2_Display/n1892 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u15_al_u4757  (
    .a({\u2_Display/n1872 ,\u2_Display/n1874 }),
    .b({\u2_Display/n1871 ,\u2_Display/n1873 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add61/c15 ),
    .f({\u2_Display/n1892 [17],\u2_Display/n1892 [15]}),
    .fco(\u2_Display/add61/c19 ),
    .fx({\u2_Display/n1892 [18],\u2_Display/n1892 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u19_al_u4758  (
    .a({\u2_Display/n1868 ,\u2_Display/n1870 }),
    .b({\u2_Display/n1867 ,\u2_Display/n1869 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add61/c19 ),
    .f({\u2_Display/n1892 [21],\u2_Display/n1892 [19]}),
    .fco(\u2_Display/add61/c23 ),
    .fx({\u2_Display/n1892 [22],\u2_Display/n1892 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u23_al_u4759  (
    .a({\u2_Display/n1864 ,\u2_Display/n1866 }),
    .b({\u2_Display/n1863 ,\u2_Display/n1865 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add61/c23 ),
    .f({\u2_Display/n1892 [25],\u2_Display/n1892 [23]}),
    .fco(\u2_Display/add61/c27 ),
    .fx({\u2_Display/n1892 [26],\u2_Display/n1892 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u27_al_u4760  (
    .a({\u2_Display/n1860 ,\u2_Display/n1862 }),
    .b({\u2_Display/n1859 ,\u2_Display/n1861 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add61/c27 ),
    .f({\u2_Display/n1892 [29],\u2_Display/n1892 [27]}),
    .fco(\u2_Display/add61/c31 ),
    .fx({\u2_Display/n1892 [30],\u2_Display/n1892 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u31_al_u4761  (
    .a({open_n64353,\u2_Display/n1858 }),
    .c(2'b00),
    .d({open_n64358,1'b1}),
    .fci(\u2_Display/add61/c31 ),
    .f({open_n64375,\u2_Display/n1892 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u3_al_u4754  (
    .a({\u2_Display/n1884 ,\u2_Display/n1886 }),
    .b({\u2_Display/n1883 ,\u2_Display/n1885 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add61/c3 ),
    .f({\u2_Display/n1892 [5],\u2_Display/n1892 [3]}),
    .fco(\u2_Display/add61/c7 ),
    .fx({\u2_Display/n1892 [6],\u2_Display/n1892 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u7_al_u4755  (
    .a({\u2_Display/n1880 ,\u2_Display/n1882 }),
    .b({\u2_Display/n1879 ,\u2_Display/n1881 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add61/c7 ),
    .f({\u2_Display/n1892 [9],\u2_Display/n1892 [7]}),
    .fco(\u2_Display/add61/c11 ),
    .fx({\u2_Display/n1892 [10],\u2_Display/n1892 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/ucin_al_u4753  (
    .a({\u2_Display/n1888 ,1'b1}),
    .b({\u2_Display/n1887 ,\u2_Display/n1889 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1892 [1],open_n64434}),
    .fco(\u2_Display/add61/c3 ),
    .fx({\u2_Display/n1892 [2],\u2_Display/n1892 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u11_al_u4765  (
    .a({\u2_Display/n1911 ,\u2_Display/n1913 }),
    .b({\u2_Display/n1910 ,\u2_Display/n1912 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add62/c11 ),
    .f({\u2_Display/n1927 [13],\u2_Display/n1927 [11]}),
    .fco(\u2_Display/add62/c15 ),
    .fx({\u2_Display/n1927 [14],\u2_Display/n1927 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u15_al_u4766  (
    .a({\u2_Display/n1907 ,\u2_Display/n1909 }),
    .b({\u2_Display/n1906 ,\u2_Display/n1908 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add62/c15 ),
    .f({\u2_Display/n1927 [17],\u2_Display/n1927 [15]}),
    .fco(\u2_Display/add62/c19 ),
    .fx({\u2_Display/n1927 [18],\u2_Display/n1927 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u19_al_u4767  (
    .a({\u2_Display/n1903 ,\u2_Display/n1905 }),
    .b({\u2_Display/n1902 ,\u2_Display/n1904 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add62/c19 ),
    .f({\u2_Display/n1927 [21],\u2_Display/n1927 [19]}),
    .fco(\u2_Display/add62/c23 ),
    .fx({\u2_Display/n1927 [22],\u2_Display/n1927 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u23_al_u4768  (
    .a({\u2_Display/n1899 ,\u2_Display/n1901 }),
    .b({\u2_Display/n1898 ,\u2_Display/n1900 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add62/c23 ),
    .f({\u2_Display/n1927 [25],\u2_Display/n1927 [23]}),
    .fco(\u2_Display/add62/c27 ),
    .fx({\u2_Display/n1927 [26],\u2_Display/n1927 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u27_al_u4769  (
    .a({\u2_Display/n1895 ,\u2_Display/n1897 }),
    .b({\u2_Display/n1894 ,\u2_Display/n1896 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add62/c27 ),
    .f({\u2_Display/n1927 [29],\u2_Display/n1927 [27]}),
    .fco(\u2_Display/add62/c31 ),
    .fx({\u2_Display/n1927 [30],\u2_Display/n1927 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u31_al_u4770  (
    .a({open_n64527,\u2_Display/n1893 }),
    .c(2'b00),
    .d({open_n64532,1'b1}),
    .fci(\u2_Display/add62/c31 ),
    .f({open_n64549,\u2_Display/n1927 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u3_al_u4763  (
    .a({\u2_Display/n1919 ,\u2_Display/n1921 }),
    .b({\u2_Display/n1918 ,\u2_Display/n1920 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add62/c3 ),
    .f({\u2_Display/n1927 [5],\u2_Display/n1927 [3]}),
    .fco(\u2_Display/add62/c7 ),
    .fx({\u2_Display/n1927 [6],\u2_Display/n1927 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u7_al_u4764  (
    .a({\u2_Display/n1915 ,\u2_Display/n1917 }),
    .b({\u2_Display/n1914 ,\u2_Display/n1916 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add62/c7 ),
    .f({\u2_Display/n1927 [9],\u2_Display/n1927 [7]}),
    .fco(\u2_Display/add62/c11 ),
    .fx({\u2_Display/n1927 [10],\u2_Display/n1927 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/ucin_al_u4762  (
    .a({\u2_Display/n1923 ,1'b1}),
    .b({\u2_Display/n1922 ,\u2_Display/n1924 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1927 [1],open_n64608}),
    .fco(\u2_Display/add62/c3 ),
    .fx({\u2_Display/n1927 [2],\u2_Display/n1927 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u11_al_u4774  (
    .a({\u2_Display/n1946 ,\u2_Display/n1948 }),
    .b({\u2_Display/n1945 ,\u2_Display/n1947 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add63/c11 ),
    .f({\u2_Display/n1962 [13],\u2_Display/n1962 [11]}),
    .fco(\u2_Display/add63/c15 ),
    .fx({\u2_Display/n1962 [14],\u2_Display/n1962 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u15_al_u4775  (
    .a({\u2_Display/n1942 ,\u2_Display/n1944 }),
    .b({\u2_Display/n1941 ,\u2_Display/n1943 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add63/c15 ),
    .f({\u2_Display/n1962 [17],\u2_Display/n1962 [15]}),
    .fco(\u2_Display/add63/c19 ),
    .fx({\u2_Display/n1962 [18],\u2_Display/n1962 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u19_al_u4776  (
    .a({\u2_Display/n1938 ,\u2_Display/n1940 }),
    .b({\u2_Display/n1937 ,\u2_Display/n1939 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add63/c19 ),
    .f({\u2_Display/n1962 [21],\u2_Display/n1962 [19]}),
    .fco(\u2_Display/add63/c23 ),
    .fx({\u2_Display/n1962 [22],\u2_Display/n1962 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u23_al_u4777  (
    .a({\u2_Display/n1934 ,\u2_Display/n1936 }),
    .b({\u2_Display/n1933 ,\u2_Display/n1935 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add63/c23 ),
    .f({\u2_Display/n1962 [25],\u2_Display/n1962 [23]}),
    .fco(\u2_Display/add63/c27 ),
    .fx({\u2_Display/n1962 [26],\u2_Display/n1962 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u27_al_u4778  (
    .a({\u2_Display/n1930 ,\u2_Display/n1932 }),
    .b({\u2_Display/n1929 ,\u2_Display/n1931 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add63/c27 ),
    .f({\u2_Display/n1962 [29],\u2_Display/n1962 [27]}),
    .fco(\u2_Display/add63/c31 ),
    .fx({\u2_Display/n1962 [30],\u2_Display/n1962 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u31_al_u4779  (
    .a({open_n64701,\u2_Display/n1928 }),
    .c(2'b00),
    .d({open_n64706,1'b1}),
    .fci(\u2_Display/add63/c31 ),
    .f({open_n64723,\u2_Display/n1962 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u3_al_u4772  (
    .a({\u2_Display/n1954 ,\u2_Display/n1956 }),
    .b({\u2_Display/n1953 ,\u2_Display/n1955 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add63/c3 ),
    .f({\u2_Display/n1962 [5],\u2_Display/n1962 [3]}),
    .fco(\u2_Display/add63/c7 ),
    .fx({\u2_Display/n1962 [6],\u2_Display/n1962 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u7_al_u4773  (
    .a({\u2_Display/n1950 ,\u2_Display/n1952 }),
    .b({\u2_Display/n1949 ,\u2_Display/n1951 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add63/c7 ),
    .f({\u2_Display/n1962 [9],\u2_Display/n1962 [7]}),
    .fco(\u2_Display/add63/c11 ),
    .fx({\u2_Display/n1962 [10],\u2_Display/n1962 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/ucin_al_u4771  (
    .a({\u2_Display/n1958 ,1'b1}),
    .b({\u2_Display/n1957 ,\u2_Display/n1959 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1962 [1],open_n64782}),
    .fco(\u2_Display/add63/c3 ),
    .fx({\u2_Display/n1962 [2],\u2_Display/n1962 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u11_al_u4783  (
    .a({\u2_Display/n1981 ,\u2_Display/n1983 }),
    .b({\u2_Display/n1980 ,\u2_Display/n1982 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add64/c11 ),
    .f({\u2_Display/n1997 [13],\u2_Display/n1997 [11]}),
    .fco(\u2_Display/add64/c15 ),
    .fx({\u2_Display/n1997 [14],\u2_Display/n1997 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u15_al_u4784  (
    .a({\u2_Display/n1977 ,\u2_Display/n1979 }),
    .b({\u2_Display/n1976 ,\u2_Display/n1978 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add64/c15 ),
    .f({\u2_Display/n1997 [17],\u2_Display/n1997 [15]}),
    .fco(\u2_Display/add64/c19 ),
    .fx({\u2_Display/n1997 [18],\u2_Display/n1997 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u19_al_u4785  (
    .a({\u2_Display/n1973 ,\u2_Display/n1975 }),
    .b({\u2_Display/n1972 ,\u2_Display/n1974 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add64/c19 ),
    .f({\u2_Display/n1997 [21],\u2_Display/n1997 [19]}),
    .fco(\u2_Display/add64/c23 ),
    .fx({\u2_Display/n1997 [22],\u2_Display/n1997 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u23_al_u4786  (
    .a({\u2_Display/n1969 ,\u2_Display/n1971 }),
    .b({\u2_Display/n1968 ,\u2_Display/n1970 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add64/c23 ),
    .f({\u2_Display/n1997 [25],\u2_Display/n1997 [23]}),
    .fco(\u2_Display/add64/c27 ),
    .fx({\u2_Display/n1997 [26],\u2_Display/n1997 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u27_al_u4787  (
    .a({\u2_Display/n1965 ,\u2_Display/n1967 }),
    .b({\u2_Display/n1964 ,\u2_Display/n1966 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add64/c27 ),
    .f({\u2_Display/n1997 [29],\u2_Display/n1997 [27]}),
    .fco(\u2_Display/add64/c31 ),
    .fx({\u2_Display/n1997 [30],\u2_Display/n1997 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u31_al_u4788  (
    .a({open_n64875,\u2_Display/n1963 }),
    .c(2'b00),
    .d({open_n64880,1'b1}),
    .fci(\u2_Display/add64/c31 ),
    .f({open_n64897,\u2_Display/n1997 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u3_al_u4781  (
    .a({\u2_Display/n1989 ,\u2_Display/n1991 }),
    .b({\u2_Display/n1988 ,\u2_Display/n1990 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add64/c3 ),
    .f({\u2_Display/n1997 [5],\u2_Display/n1997 [3]}),
    .fco(\u2_Display/add64/c7 ),
    .fx({\u2_Display/n1997 [6],\u2_Display/n1997 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u7_al_u4782  (
    .a({\u2_Display/n1985 ,\u2_Display/n1987 }),
    .b({\u2_Display/n1984 ,\u2_Display/n1986 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add64/c7 ),
    .f({\u2_Display/n1997 [9],\u2_Display/n1997 [7]}),
    .fco(\u2_Display/add64/c11 ),
    .fx({\u2_Display/n1997 [10],\u2_Display/n1997 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/ucin_al_u4780  (
    .a({\u2_Display/n1993 ,1'b1}),
    .b({\u2_Display/n1992 ,\u2_Display/n1994 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1997 [1],open_n64956}),
    .fco(\u2_Display/add64/c3 ),
    .fx({\u2_Display/n1997 [2],\u2_Display/n1997 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u11_al_u4792  (
    .a({\u2_Display/n2016 ,\u2_Display/n2018 }),
    .b({\u2_Display/n2015 ,\u2_Display/n2017 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add65/c11 ),
    .f({\u2_Display/n2032 [13],\u2_Display/n2032 [11]}),
    .fco(\u2_Display/add65/c15 ),
    .fx({\u2_Display/n2032 [14],\u2_Display/n2032 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u15_al_u4793  (
    .a({\u2_Display/n2012 ,\u2_Display/n2014 }),
    .b({\u2_Display/n2011 ,\u2_Display/n2013 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add65/c15 ),
    .f({\u2_Display/n2032 [17],\u2_Display/n2032 [15]}),
    .fco(\u2_Display/add65/c19 ),
    .fx({\u2_Display/n2032 [18],\u2_Display/n2032 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u19_al_u4794  (
    .a({\u2_Display/n2008 ,\u2_Display/n2010 }),
    .b({\u2_Display/n2007 ,\u2_Display/n2009 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add65/c19 ),
    .f({\u2_Display/n2032 [21],\u2_Display/n2032 [19]}),
    .fco(\u2_Display/add65/c23 ),
    .fx({\u2_Display/n2032 [22],\u2_Display/n2032 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u23_al_u4795  (
    .a({\u2_Display/n2004 ,\u2_Display/n2006 }),
    .b({\u2_Display/n2003 ,\u2_Display/n2005 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add65/c23 ),
    .f({\u2_Display/n2032 [25],\u2_Display/n2032 [23]}),
    .fco(\u2_Display/add65/c27 ),
    .fx({\u2_Display/n2032 [26],\u2_Display/n2032 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u27_al_u4796  (
    .a({\u2_Display/n2000 ,\u2_Display/n2002 }),
    .b({\u2_Display/n1999 ,\u2_Display/n2001 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add65/c27 ),
    .f({\u2_Display/n2032 [29],\u2_Display/n2032 [27]}),
    .fco(\u2_Display/add65/c31 ),
    .fx({\u2_Display/n2032 [30],\u2_Display/n2032 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u31_al_u4797  (
    .a({open_n65049,\u2_Display/n1998 }),
    .c(2'b00),
    .d({open_n65054,1'b1}),
    .fci(\u2_Display/add65/c31 ),
    .f({open_n65071,\u2_Display/n2032 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u3_al_u4790  (
    .a({\u2_Display/n2024 ,\u2_Display/n2026 }),
    .b({\u2_Display/n2023 ,\u2_Display/n2025 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add65/c3 ),
    .f({\u2_Display/n2032 [5],\u2_Display/n2032 [3]}),
    .fco(\u2_Display/add65/c7 ),
    .fx({\u2_Display/n2032 [6],\u2_Display/n2032 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u7_al_u4791  (
    .a({\u2_Display/n2020 ,\u2_Display/n2022 }),
    .b({\u2_Display/n2019 ,\u2_Display/n2021 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add65/c7 ),
    .f({\u2_Display/n2032 [9],\u2_Display/n2032 [7]}),
    .fco(\u2_Display/add65/c11 ),
    .fx({\u2_Display/n2032 [10],\u2_Display/n2032 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/ucin_al_u4789  (
    .a({\u2_Display/n2028 ,1'b1}),
    .b({\u2_Display/n2027 ,\u2_Display/n2029 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2032 [1],open_n65130}),
    .fco(\u2_Display/add65/c3 ),
    .fx({\u2_Display/n2032 [2],\u2_Display/n2032 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u11_al_u4801  (
    .a({\u2_Display/n2051 ,\u2_Display/n2053 }),
    .b({\u2_Display/n2050 ,\u2_Display/n2052 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add66/c11 ),
    .f({\u2_Display/n2067 [13],\u2_Display/n2067 [11]}),
    .fco(\u2_Display/add66/c15 ),
    .fx({\u2_Display/n2067 [14],\u2_Display/n2067 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u15_al_u4802  (
    .a({\u2_Display/n2047 ,\u2_Display/n2049 }),
    .b({\u2_Display/n2046 ,\u2_Display/n2048 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add66/c15 ),
    .f({\u2_Display/n2067 [17],\u2_Display/n2067 [15]}),
    .fco(\u2_Display/add66/c19 ),
    .fx({\u2_Display/n2067 [18],\u2_Display/n2067 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u19_al_u4803  (
    .a({\u2_Display/n2043 ,\u2_Display/n2045 }),
    .b({\u2_Display/n2042 ,\u2_Display/n2044 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add66/c19 ),
    .f({\u2_Display/n2067 [21],\u2_Display/n2067 [19]}),
    .fco(\u2_Display/add66/c23 ),
    .fx({\u2_Display/n2067 [22],\u2_Display/n2067 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u23_al_u4804  (
    .a({\u2_Display/n2039 ,\u2_Display/n2041 }),
    .b({\u2_Display/n2038 ,\u2_Display/n2040 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add66/c23 ),
    .f({\u2_Display/n2067 [25],\u2_Display/n2067 [23]}),
    .fco(\u2_Display/add66/c27 ),
    .fx({\u2_Display/n2067 [26],\u2_Display/n2067 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u27_al_u4805  (
    .a({\u2_Display/n2035 ,\u2_Display/n2037 }),
    .b({\u2_Display/n2034 ,\u2_Display/n2036 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add66/c27 ),
    .f({\u2_Display/n2067 [29],\u2_Display/n2067 [27]}),
    .fco(\u2_Display/add66/c31 ),
    .fx({\u2_Display/n2067 [30],\u2_Display/n2067 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u31_al_u4806  (
    .a({open_n65223,\u2_Display/n2033 }),
    .c(2'b00),
    .d({open_n65228,1'b1}),
    .fci(\u2_Display/add66/c31 ),
    .f({open_n65245,\u2_Display/n2067 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u3_al_u4799  (
    .a({\u2_Display/n2059 ,\u2_Display/n2061 }),
    .b({\u2_Display/n2058 ,\u2_Display/n2060 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add66/c3 ),
    .f({\u2_Display/n2067 [5],\u2_Display/n2067 [3]}),
    .fco(\u2_Display/add66/c7 ),
    .fx({\u2_Display/n2067 [6],\u2_Display/n2067 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u7_al_u4800  (
    .a({\u2_Display/n2055 ,\u2_Display/n2057 }),
    .b({\u2_Display/n2054 ,\u2_Display/n2056 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add66/c7 ),
    .f({\u2_Display/n2067 [9],\u2_Display/n2067 [7]}),
    .fco(\u2_Display/add66/c11 ),
    .fx({\u2_Display/n2067 [10],\u2_Display/n2067 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/ucin_al_u4798  (
    .a({\u2_Display/n2063 ,1'b1}),
    .b({\u2_Display/n2062 ,\u2_Display/n2064 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2067 [1],open_n65304}),
    .fco(\u2_Display/add66/c3 ),
    .fx({\u2_Display/n2067 [2],\u2_Display/n2067 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u11_al_u4810  (
    .a({\u2_Display/n2086 ,\u2_Display/n2088 }),
    .b({\u2_Display/n2085 ,\u2_Display/n2087 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add67/c11 ),
    .f({\u2_Display/n2102 [13],\u2_Display/n2102 [11]}),
    .fco(\u2_Display/add67/c15 ),
    .fx({\u2_Display/n2102 [14],\u2_Display/n2102 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u15_al_u4811  (
    .a({\u2_Display/n2082 ,\u2_Display/n2084 }),
    .b({\u2_Display/n2081 ,\u2_Display/n2083 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add67/c15 ),
    .f({\u2_Display/n2102 [17],\u2_Display/n2102 [15]}),
    .fco(\u2_Display/add67/c19 ),
    .fx({\u2_Display/n2102 [18],\u2_Display/n2102 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u19_al_u4812  (
    .a({\u2_Display/n2078 ,\u2_Display/n2080 }),
    .b({\u2_Display/n2077 ,\u2_Display/n2079 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add67/c19 ),
    .f({\u2_Display/n2102 [21],\u2_Display/n2102 [19]}),
    .fco(\u2_Display/add67/c23 ),
    .fx({\u2_Display/n2102 [22],\u2_Display/n2102 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u23_al_u4813  (
    .a({\u2_Display/n2074 ,\u2_Display/n2076 }),
    .b({\u2_Display/n2073 ,\u2_Display/n2075 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add67/c23 ),
    .f({\u2_Display/n2102 [25],\u2_Display/n2102 [23]}),
    .fco(\u2_Display/add67/c27 ),
    .fx({\u2_Display/n2102 [26],\u2_Display/n2102 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u27_al_u4814  (
    .a({\u2_Display/n2070 ,\u2_Display/n2072 }),
    .b({\u2_Display/n2069 ,\u2_Display/n2071 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add67/c27 ),
    .f({\u2_Display/n2102 [29],\u2_Display/n2102 [27]}),
    .fco(\u2_Display/add67/c31 ),
    .fx({\u2_Display/n2102 [30],\u2_Display/n2102 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u31_al_u4815  (
    .a({open_n65397,\u2_Display/n2068 }),
    .c(2'b00),
    .d({open_n65402,1'b1}),
    .fci(\u2_Display/add67/c31 ),
    .f({open_n65419,\u2_Display/n2102 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u3_al_u4808  (
    .a({\u2_Display/n2094 ,\u2_Display/n2096 }),
    .b({\u2_Display/n2093 ,\u2_Display/n2095 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add67/c3 ),
    .f({\u2_Display/n2102 [5],\u2_Display/n2102 [3]}),
    .fco(\u2_Display/add67/c7 ),
    .fx({\u2_Display/n2102 [6],\u2_Display/n2102 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u7_al_u4809  (
    .a({\u2_Display/n2090 ,\u2_Display/n2092 }),
    .b({\u2_Display/n2089 ,\u2_Display/n2091 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add67/c7 ),
    .f({\u2_Display/n2102 [9],\u2_Display/n2102 [7]}),
    .fco(\u2_Display/add67/c11 ),
    .fx({\u2_Display/n2102 [10],\u2_Display/n2102 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/ucin_al_u4807  (
    .a({\u2_Display/n2098 ,1'b1}),
    .b({\u2_Display/n2097 ,\u2_Display/n2099 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2102 [1],open_n65478}),
    .fco(\u2_Display/add67/c3 ),
    .fx({\u2_Display/n2102 [2],\u2_Display/n2102 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u11_al_u4819  (
    .a({\u2_Display/n2121 ,\u2_Display/n2123 }),
    .b({\u2_Display/n2120 ,\u2_Display/n2122 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add68/c11 ),
    .f({\u2_Display/n2137 [13],\u2_Display/n2137 [11]}),
    .fco(\u2_Display/add68/c15 ),
    .fx({\u2_Display/n2137 [14],\u2_Display/n2137 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u15_al_u4820  (
    .a({\u2_Display/n2117 ,\u2_Display/n2119 }),
    .b({\u2_Display/n2116 ,\u2_Display/n2118 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add68/c15 ),
    .f({\u2_Display/n2137 [17],\u2_Display/n2137 [15]}),
    .fco(\u2_Display/add68/c19 ),
    .fx({\u2_Display/n2137 [18],\u2_Display/n2137 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u19_al_u4821  (
    .a({\u2_Display/n2113 ,\u2_Display/n2115 }),
    .b({\u2_Display/n2112 ,\u2_Display/n2114 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add68/c19 ),
    .f({\u2_Display/n2137 [21],\u2_Display/n2137 [19]}),
    .fco(\u2_Display/add68/c23 ),
    .fx({\u2_Display/n2137 [22],\u2_Display/n2137 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u23_al_u4822  (
    .a({\u2_Display/n2109 ,\u2_Display/n2111 }),
    .b({\u2_Display/n2108 ,\u2_Display/n2110 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add68/c23 ),
    .f({\u2_Display/n2137 [25],\u2_Display/n2137 [23]}),
    .fco(\u2_Display/add68/c27 ),
    .fx({\u2_Display/n2137 [26],\u2_Display/n2137 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u27_al_u4823  (
    .a({\u2_Display/n2105 ,\u2_Display/n2107 }),
    .b({\u2_Display/n2104 ,\u2_Display/n2106 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add68/c27 ),
    .f({\u2_Display/n2137 [29],\u2_Display/n2137 [27]}),
    .fco(\u2_Display/add68/c31 ),
    .fx({\u2_Display/n2137 [30],\u2_Display/n2137 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u31_al_u4824  (
    .a({open_n65571,\u2_Display/n2103 }),
    .c(2'b00),
    .d({open_n65576,1'b1}),
    .fci(\u2_Display/add68/c31 ),
    .f({open_n65593,\u2_Display/n2137 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u3_al_u4817  (
    .a({\u2_Display/n2129 ,\u2_Display/n2131 }),
    .b({\u2_Display/n2128 ,\u2_Display/n2130 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add68/c3 ),
    .f({\u2_Display/n2137 [5],\u2_Display/n2137 [3]}),
    .fco(\u2_Display/add68/c7 ),
    .fx({\u2_Display/n2137 [6],\u2_Display/n2137 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u7_al_u4818  (
    .a({\u2_Display/n2125 ,\u2_Display/n2127 }),
    .b({\u2_Display/n2124 ,\u2_Display/n2126 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add68/c7 ),
    .f({\u2_Display/n2137 [9],\u2_Display/n2137 [7]}),
    .fco(\u2_Display/add68/c11 ),
    .fx({\u2_Display/n2137 [10],\u2_Display/n2137 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/ucin_al_u4816  (
    .a({\u2_Display/n2133 ,1'b1}),
    .b({\u2_Display/n2132 ,\u2_Display/n2134 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2137 [1],open_n65652}),
    .fco(\u2_Display/add68/c3 ),
    .fx({\u2_Display/n2137 [2],\u2_Display/n2137 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u11_al_u4828  (
    .a({\u2_Display/n2156 ,\u2_Display/n2158 }),
    .b({\u2_Display/n2155 ,\u2_Display/n2157 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add69/c11 ),
    .f({\u2_Display/n2172 [13],\u2_Display/n2172 [11]}),
    .fco(\u2_Display/add69/c15 ),
    .fx({\u2_Display/n2172 [14],\u2_Display/n2172 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u15_al_u4829  (
    .a({\u2_Display/n2152 ,\u2_Display/n2154 }),
    .b({\u2_Display/n2151 ,\u2_Display/n2153 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add69/c15 ),
    .f({\u2_Display/n2172 [17],\u2_Display/n2172 [15]}),
    .fco(\u2_Display/add69/c19 ),
    .fx({\u2_Display/n2172 [18],\u2_Display/n2172 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u19_al_u4830  (
    .a({\u2_Display/n2148 ,\u2_Display/n2150 }),
    .b({\u2_Display/n2147 ,\u2_Display/n2149 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add69/c19 ),
    .f({\u2_Display/n2172 [21],\u2_Display/n2172 [19]}),
    .fco(\u2_Display/add69/c23 ),
    .fx({\u2_Display/n2172 [22],\u2_Display/n2172 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u23_al_u4831  (
    .a({\u2_Display/n2144 ,\u2_Display/n2146 }),
    .b({\u2_Display/n2143 ,\u2_Display/n2145 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add69/c23 ),
    .f({\u2_Display/n2172 [25],\u2_Display/n2172 [23]}),
    .fco(\u2_Display/add69/c27 ),
    .fx({\u2_Display/n2172 [26],\u2_Display/n2172 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u27_al_u4832  (
    .a({\u2_Display/n2140 ,\u2_Display/n2142 }),
    .b({\u2_Display/n2139 ,\u2_Display/n2141 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add69/c27 ),
    .f({\u2_Display/n2172 [29],\u2_Display/n2172 [27]}),
    .fco(\u2_Display/add69/c31 ),
    .fx({\u2_Display/n2172 [30],\u2_Display/n2172 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u31_al_u4833  (
    .a({open_n65745,\u2_Display/n2138 }),
    .c(2'b00),
    .d({open_n65750,1'b1}),
    .fci(\u2_Display/add69/c31 ),
    .f({open_n65767,\u2_Display/n2172 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u3_al_u4826  (
    .a({\u2_Display/n2164 ,\u2_Display/n2166 }),
    .b({\u2_Display/n2163 ,\u2_Display/n2165 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add69/c3 ),
    .f({\u2_Display/n2172 [5],\u2_Display/n2172 [3]}),
    .fco(\u2_Display/add69/c7 ),
    .fx({\u2_Display/n2172 [6],\u2_Display/n2172 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u7_al_u4827  (
    .a({\u2_Display/n2160 ,\u2_Display/n2162 }),
    .b({\u2_Display/n2159 ,\u2_Display/n2161 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add69/c7 ),
    .f({\u2_Display/n2172 [9],\u2_Display/n2172 [7]}),
    .fco(\u2_Display/add69/c11 ),
    .fx({\u2_Display/n2172 [10],\u2_Display/n2172 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/ucin_al_u4825  (
    .a({\u2_Display/n2168 ,1'b1}),
    .b({\u2_Display/n2167 ,\u2_Display/n2169 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2172 [1],open_n65826}),
    .fco(\u2_Display/add69/c3 ),
    .fx({\u2_Display/n2172 [2],\u2_Display/n2172 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add6_2/u0|u2_Display/add6_2/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add6_2/u0|u2_Display/add6_2/ucin  (
    .a(2'b10),
    .b({\u2_Display/j [7],open_n65829}),
    .f({\u2_Display/n135 [0],open_n65849}),
    .fco(\u2_Display/add6_2/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add6_2/u0|u2_Display/add6_2/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add6_2/u2|u2_Display/add6_2/u1  (
    .a(2'b10),
    .b(\u2_Display/j [9:8]),
    .fci(\u2_Display/add6_2/c1 ),
    .f(\u2_Display/n135 [2:1]),
    .fco(\u2_Display/add6_2/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add6_2/u0|u2_Display/add6_2/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add6_2/ucout_al_u5059  (
    .fci(\u2_Display/add6_2/c3 ),
    .f({open_n65898,\u2_Display/add6_2_co }));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u11_al_u4837  (
    .a({\u2_Display/n2191 ,\u2_Display/n2193 }),
    .b({\u2_Display/n2190 ,\u2_Display/n2192 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add70/c11 ),
    .f({\u2_Display/n2207 [13],\u2_Display/n2207 [11]}),
    .fco(\u2_Display/add70/c15 ),
    .fx({\u2_Display/n2207 [14],\u2_Display/n2207 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u15_al_u4838  (
    .a({\u2_Display/n2187 ,\u2_Display/n2189 }),
    .b({\u2_Display/n2186 ,\u2_Display/n2188 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add70/c15 ),
    .f({\u2_Display/n2207 [17],\u2_Display/n2207 [15]}),
    .fco(\u2_Display/add70/c19 ),
    .fx({\u2_Display/n2207 [18],\u2_Display/n2207 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u19_al_u4839  (
    .a({\u2_Display/n2183 ,\u2_Display/n2185 }),
    .b({\u2_Display/n2182 ,\u2_Display/n2184 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add70/c19 ),
    .f({\u2_Display/n2207 [21],\u2_Display/n2207 [19]}),
    .fco(\u2_Display/add70/c23 ),
    .fx({\u2_Display/n2207 [22],\u2_Display/n2207 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u23_al_u4840  (
    .a({\u2_Display/n2179 ,\u2_Display/n2181 }),
    .b({\u2_Display/n2178 ,\u2_Display/n2180 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add70/c23 ),
    .f({\u2_Display/n2207 [25],\u2_Display/n2207 [23]}),
    .fco(\u2_Display/add70/c27 ),
    .fx({\u2_Display/n2207 [26],\u2_Display/n2207 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u27_al_u4841  (
    .a({\u2_Display/n2175 ,\u2_Display/n2177 }),
    .b({\u2_Display/n2174 ,\u2_Display/n2176 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add70/c27 ),
    .f({\u2_Display/n2207 [29],\u2_Display/n2207 [27]}),
    .fco(\u2_Display/add70/c31 ),
    .fx({\u2_Display/n2207 [30],\u2_Display/n2207 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u31_al_u4842  (
    .a({open_n65994,\u2_Display/n2173 }),
    .c(2'b00),
    .d({open_n65999,1'b1}),
    .fci(\u2_Display/add70/c31 ),
    .f({open_n66016,\u2_Display/n2207 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u3_al_u4835  (
    .a({\u2_Display/n2199 ,\u2_Display/n2201 }),
    .b({\u2_Display/n2198 ,\u2_Display/n2200 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add70/c3 ),
    .f({\u2_Display/n2207 [5],\u2_Display/n2207 [3]}),
    .fco(\u2_Display/add70/c7 ),
    .fx({\u2_Display/n2207 [6],\u2_Display/n2207 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u7_al_u4836  (
    .a({\u2_Display/n2195 ,\u2_Display/n2197 }),
    .b({\u2_Display/n2194 ,\u2_Display/n2196 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add70/c7 ),
    .f({\u2_Display/n2207 [9],\u2_Display/n2207 [7]}),
    .fco(\u2_Display/add70/c11 ),
    .fx({\u2_Display/n2207 [10],\u2_Display/n2207 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/ucin_al_u4834  (
    .a({\u2_Display/n2203 ,1'b1}),
    .b({\u2_Display/n2202 ,\u2_Display/n2204 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2207 [1],open_n66075}),
    .fco(\u2_Display/add70/c3 ),
    .fx({\u2_Display/n2207 [2],\u2_Display/n2207 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u11_al_u4846  (
    .a({\u2_Display/n2226 ,\u2_Display/n2228 }),
    .b({\u2_Display/n2225 ,\u2_Display/n2227 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add71/c11 ),
    .f({\u2_Display/n2242 [13],\u2_Display/n2242 [11]}),
    .fco(\u2_Display/add71/c15 ),
    .fx({\u2_Display/n2242 [14],\u2_Display/n2242 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u15_al_u4847  (
    .a({\u2_Display/n2222 ,\u2_Display/n2224 }),
    .b({\u2_Display/n2221 ,\u2_Display/n2223 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add71/c15 ),
    .f({\u2_Display/n2242 [17],\u2_Display/n2242 [15]}),
    .fco(\u2_Display/add71/c19 ),
    .fx({\u2_Display/n2242 [18],\u2_Display/n2242 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u19_al_u4848  (
    .a({\u2_Display/n2218 ,\u2_Display/n2220 }),
    .b({\u2_Display/n2217 ,\u2_Display/n2219 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add71/c19 ),
    .f({\u2_Display/n2242 [21],\u2_Display/n2242 [19]}),
    .fco(\u2_Display/add71/c23 ),
    .fx({\u2_Display/n2242 [22],\u2_Display/n2242 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u23_al_u4849  (
    .a({\u2_Display/n2214 ,\u2_Display/n2216 }),
    .b({\u2_Display/n2213 ,\u2_Display/n2215 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add71/c23 ),
    .f({\u2_Display/n2242 [25],\u2_Display/n2242 [23]}),
    .fco(\u2_Display/add71/c27 ),
    .fx({\u2_Display/n2242 [26],\u2_Display/n2242 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u27_al_u4850  (
    .a({\u2_Display/n2210 ,\u2_Display/n2212 }),
    .b({\u2_Display/n2209 ,\u2_Display/n2211 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add71/c27 ),
    .f({\u2_Display/n2242 [29],\u2_Display/n2242 [27]}),
    .fco(\u2_Display/add71/c31 ),
    .fx({\u2_Display/n2242 [30],\u2_Display/n2242 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u31_al_u4851  (
    .a({open_n66168,\u2_Display/n2208 }),
    .c(2'b00),
    .d({open_n66173,1'b1}),
    .fci(\u2_Display/add71/c31 ),
    .f({open_n66190,\u2_Display/n2242 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u3_al_u4844  (
    .a({\u2_Display/n2234 ,\u2_Display/n2236 }),
    .b({\u2_Display/n2233 ,\u2_Display/n2235 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add71/c3 ),
    .f({\u2_Display/n2242 [5],\u2_Display/n2242 [3]}),
    .fco(\u2_Display/add71/c7 ),
    .fx({\u2_Display/n2242 [6],\u2_Display/n2242 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u7_al_u4845  (
    .a({\u2_Display/n2230 ,\u2_Display/n2232 }),
    .b({\u2_Display/n2229 ,\u2_Display/n2231 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add71/c7 ),
    .f({\u2_Display/n2242 [9],\u2_Display/n2242 [7]}),
    .fco(\u2_Display/add71/c11 ),
    .fx({\u2_Display/n2242 [10],\u2_Display/n2242 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/ucin_al_u4843  (
    .a({\u2_Display/n2238 ,1'b1}),
    .b({\u2_Display/n2237 ,\u2_Display/n2239 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2242 [1],open_n66249}),
    .fco(\u2_Display/add71/c3 ),
    .fx({\u2_Display/n2242 [2],\u2_Display/n2242 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u11_al_u4855  (
    .a({\u2_Display/n2261 ,\u2_Display/n2263 }),
    .b({\u2_Display/n2260 ,\u2_Display/n2262 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add72/c11 ),
    .f({\u2_Display/n2277 [13],\u2_Display/n2277 [11]}),
    .fco(\u2_Display/add72/c15 ),
    .fx({\u2_Display/n2277 [14],\u2_Display/n2277 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u15_al_u4856  (
    .a({\u2_Display/n2257 ,\u2_Display/n2259 }),
    .b({\u2_Display/n2256 ,\u2_Display/n2258 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add72/c15 ),
    .f({\u2_Display/n2277 [17],\u2_Display/n2277 [15]}),
    .fco(\u2_Display/add72/c19 ),
    .fx({\u2_Display/n2277 [18],\u2_Display/n2277 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u19_al_u4857  (
    .a({\u2_Display/n2253 ,\u2_Display/n2255 }),
    .b({\u2_Display/n2252 ,\u2_Display/n2254 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add72/c19 ),
    .f({\u2_Display/n2277 [21],\u2_Display/n2277 [19]}),
    .fco(\u2_Display/add72/c23 ),
    .fx({\u2_Display/n2277 [22],\u2_Display/n2277 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u23_al_u4858  (
    .a({\u2_Display/n2249 ,\u2_Display/n2251 }),
    .b({\u2_Display/n2248 ,\u2_Display/n2250 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add72/c23 ),
    .f({\u2_Display/n2277 [25],\u2_Display/n2277 [23]}),
    .fco(\u2_Display/add72/c27 ),
    .fx({\u2_Display/n2277 [26],\u2_Display/n2277 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u27_al_u4859  (
    .a({\u2_Display/n2245 ,\u2_Display/n2247 }),
    .b({\u2_Display/n2244 ,\u2_Display/n2246 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add72/c27 ),
    .f({\u2_Display/n2277 [29],\u2_Display/n2277 [27]}),
    .fco(\u2_Display/add72/c31 ),
    .fx({\u2_Display/n2277 [30],\u2_Display/n2277 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u31_al_u4860  (
    .a({open_n66342,\u2_Display/n2243 }),
    .c(2'b00),
    .d({open_n66347,1'b1}),
    .fci(\u2_Display/add72/c31 ),
    .f({open_n66364,\u2_Display/n2277 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u3_al_u4853  (
    .a({\u2_Display/n2269 ,\u2_Display/n2271 }),
    .b({\u2_Display/n2268 ,\u2_Display/n2270 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add72/c3 ),
    .f({\u2_Display/n2277 [5],\u2_Display/n2277 [3]}),
    .fco(\u2_Display/add72/c7 ),
    .fx({\u2_Display/n2277 [6],\u2_Display/n2277 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u7_al_u4854  (
    .a({\u2_Display/n2265 ,\u2_Display/n2267 }),
    .b({\u2_Display/n2264 ,\u2_Display/n2266 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add72/c7 ),
    .f({\u2_Display/n2277 [9],\u2_Display/n2277 [7]}),
    .fco(\u2_Display/add72/c11 ),
    .fx({\u2_Display/n2277 [10],\u2_Display/n2277 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/ucin_al_u4852  (
    .a({\u2_Display/n2273 ,1'b1}),
    .b({\u2_Display/n2272 ,\u2_Display/n2274 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2277 [1],open_n66423}),
    .fco(\u2_Display/add72/c3 ),
    .fx({\u2_Display/n2277 [2],\u2_Display/n2277 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add73/ucin_al_u5055"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add73/u3_al_u5056  (
    .a({\u2_Display/n2304 ,\u2_Display/n2306 }),
    .b({\u2_Display/n2303 ,\u2_Display/n2305 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add73/c3 ),
    .f({\u2_Display/n2312 [5],\u2_Display/n2312 [3]}),
    .fco(\u2_Display/add73/c7 ),
    .fx({\u2_Display/n2312 [6],\u2_Display/n2312 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add73/ucin_al_u5055"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add73/u7_al_u5057  (
    .a({\u2_Display/n2300 ,\u2_Display/n2302 }),
    .b({open_n66444,\u2_Display/n2301 }),
    .c(2'b00),
    .d(2'b00),
    .e({open_n66447,1'b0}),
    .fci(\u2_Display/add73/c7 ),
    .f({\u2_Display/n2312 [9],\u2_Display/n2312 [7]}),
    .fx({open_n66463,\u2_Display/n2312 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add73/ucin_al_u5055"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add73/ucin_al_u5055  (
    .a({\u2_Display/n2308 ,1'b1}),
    .b({\u2_Display/n2307 ,\u2_Display/n2309 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .f({\u2_Display/n2312 [1],open_n66483}),
    .fco(\u2_Display/add73/c3 ),
    .fx({\u2_Display/n2312 [2],\u2_Display/n2312 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u11_al_u4864  (
    .a({\u2_Display/counta [13],\u2_Display/counta [11]}),
    .b({\u2_Display/counta [14],\u2_Display/counta [12]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add84/c11 ),
    .f({\u2_Display/n2665 [13],\u2_Display/n2665 [11]}),
    .fco(\u2_Display/add84/c15 ),
    .fx({\u2_Display/n2665 [14],\u2_Display/n2665 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u15_al_u4865  (
    .a({\u2_Display/counta [17],\u2_Display/counta [15]}),
    .b({\u2_Display/counta [18],\u2_Display/counta [16]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add84/c15 ),
    .f({\u2_Display/n2665 [17],\u2_Display/n2665 [15]}),
    .fco(\u2_Display/add84/c19 ),
    .fx({\u2_Display/n2665 [18],\u2_Display/n2665 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u19_al_u4866  (
    .a({\u2_Display/counta [21],\u2_Display/counta [19]}),
    .b({\u2_Display/counta [22],\u2_Display/counta [20]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add84/c19 ),
    .f({\u2_Display/n2665 [21],\u2_Display/n2665 [19]}),
    .fco(\u2_Display/add84/c23 ),
    .fx({\u2_Display/n2665 [22],\u2_Display/n2665 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u23_al_u4867  (
    .a({\u2_Display/counta [25],\u2_Display/counta [23]}),
    .b({\u2_Display/counta [26],\u2_Display/counta [24]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add84/c23 ),
    .f({\u2_Display/n2665 [25],\u2_Display/n2665 [23]}),
    .fco(\u2_Display/add84/c27 ),
    .fx({\u2_Display/n2665 [26],\u2_Display/n2665 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u27_al_u4868  (
    .a({\u2_Display/counta [29],\u2_Display/counta [27]}),
    .b({\u2_Display/counta [30],\u2_Display/counta [28]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add84/c27 ),
    .f({\u2_Display/n2665 [29],\u2_Display/n2665 [27]}),
    .fco(\u2_Display/add84/c31 ),
    .fx({\u2_Display/n2665 [30],\u2_Display/n2665 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u31_al_u4869  (
    .a({open_n66576,\u2_Display/counta [31]}),
    .c(2'b00),
    .d({open_n66581,1'b0}),
    .fci(\u2_Display/add84/c31 ),
    .f({open_n66598,\u2_Display/n2665 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u3_al_u4862  (
    .a({\u2_Display/counta [5],\u2_Display/counta [3]}),
    .b({\u2_Display/counta [6],\u2_Display/counta [4]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add84/c3 ),
    .f({\u2_Display/n2665 [5],\u2_Display/n2665 [3]}),
    .fco(\u2_Display/add84/c7 ),
    .fx({\u2_Display/n2665 [6],\u2_Display/n2665 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u7_al_u4863  (
    .a({\u2_Display/counta [9],\u2_Display/counta [7]}),
    .b({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add84/c7 ),
    .f({\u2_Display/n2665 [9],\u2_Display/n2665 [7]}),
    .fco(\u2_Display/add84/c11 ),
    .fx({\u2_Display/n2665 [10],\u2_Display/n2665 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/ucin_al_u4861  (
    .a({\u2_Display/counta [1],1'b1}),
    .b({\u2_Display/counta [2],\u2_Display/counta [0]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2665 [1],open_n66657}),
    .fco(\u2_Display/add84/c3 ),
    .fx({\u2_Display/n2665 [2],\u2_Display/n2665 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u11_al_u4873  (
    .a({\u2_Display/n2684 ,\u2_Display/n2686 }),
    .b({\u2_Display/n2683 ,\u2_Display/n2685 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add85/c11 ),
    .f({\u2_Display/n2700 [13],\u2_Display/n2700 [11]}),
    .fco(\u2_Display/add85/c15 ),
    .fx({\u2_Display/n2700 [14],\u2_Display/n2700 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u15_al_u4874  (
    .a({\u2_Display/n2680 ,\u2_Display/n2682 }),
    .b({\u2_Display/n2679 ,\u2_Display/n2681 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add85/c15 ),
    .f({\u2_Display/n2700 [17],\u2_Display/n2700 [15]}),
    .fco(\u2_Display/add85/c19 ),
    .fx({\u2_Display/n2700 [18],\u2_Display/n2700 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u19_al_u4875  (
    .a({\u2_Display/n2676 ,\u2_Display/n2678 }),
    .b({\u2_Display/n2675 ,\u2_Display/n2677 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add85/c19 ),
    .f({\u2_Display/n2700 [21],\u2_Display/n2700 [19]}),
    .fco(\u2_Display/add85/c23 ),
    .fx({\u2_Display/n2700 [22],\u2_Display/n2700 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u23_al_u4876  (
    .a({\u2_Display/n2672 ,\u2_Display/n2674 }),
    .b({\u2_Display/n2671 ,\u2_Display/n2673 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add85/c23 ),
    .f({\u2_Display/n2700 [25],\u2_Display/n2700 [23]}),
    .fco(\u2_Display/add85/c27 ),
    .fx({\u2_Display/n2700 [26],\u2_Display/n2700 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u27_al_u4877  (
    .a({\u2_Display/n2668 ,\u2_Display/n2670 }),
    .b({\u2_Display/n2667 ,\u2_Display/n2669 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add85/c27 ),
    .f({\u2_Display/n2700 [29],\u2_Display/n2700 [27]}),
    .fco(\u2_Display/add85/c31 ),
    .fx({\u2_Display/n2700 [30],\u2_Display/n2700 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u31_al_u4878  (
    .a({open_n66750,\u2_Display/n2666 }),
    .c(2'b00),
    .d({open_n66755,1'b1}),
    .fci(\u2_Display/add85/c31 ),
    .f({open_n66772,\u2_Display/n2700 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u3_al_u4871  (
    .a({\u2_Display/n2692 ,\u2_Display/n2694 }),
    .b({\u2_Display/n2691 ,\u2_Display/n2693 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add85/c3 ),
    .f({\u2_Display/n2700 [5],\u2_Display/n2700 [3]}),
    .fco(\u2_Display/add85/c7 ),
    .fx({\u2_Display/n2700 [6],\u2_Display/n2700 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u7_al_u4872  (
    .a({\u2_Display/n2688 ,\u2_Display/n2690 }),
    .b({\u2_Display/n2687 ,\u2_Display/n2689 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add85/c7 ),
    .f({\u2_Display/n2700 [9],\u2_Display/n2700 [7]}),
    .fco(\u2_Display/add85/c11 ),
    .fx({\u2_Display/n2700 [10],\u2_Display/n2700 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/ucin_al_u4870  (
    .a({\u2_Display/n2696 ,1'b1}),
    .b({\u2_Display/n2695 ,\u2_Display/n2697 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2700 [1],open_n66831}),
    .fco(\u2_Display/add85/c3 ),
    .fx({\u2_Display/n2700 [2],\u2_Display/n2700 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u11_al_u4882  (
    .a({\u2_Display/n2719 ,\u2_Display/n2721 }),
    .b({\u2_Display/n2718 ,\u2_Display/n2720 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add86/c11 ),
    .f({\u2_Display/n2735 [13],\u2_Display/n2735 [11]}),
    .fco(\u2_Display/add86/c15 ),
    .fx({\u2_Display/n2735 [14],\u2_Display/n2735 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u15_al_u4883  (
    .a({\u2_Display/n2715 ,\u2_Display/n2717 }),
    .b({\u2_Display/n2714 ,\u2_Display/n2716 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add86/c15 ),
    .f({\u2_Display/n2735 [17],\u2_Display/n2735 [15]}),
    .fco(\u2_Display/add86/c19 ),
    .fx({\u2_Display/n2735 [18],\u2_Display/n2735 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u19_al_u4884  (
    .a({\u2_Display/n2711 ,\u2_Display/n2713 }),
    .b({\u2_Display/n2710 ,\u2_Display/n2712 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add86/c19 ),
    .f({\u2_Display/n2735 [21],\u2_Display/n2735 [19]}),
    .fco(\u2_Display/add86/c23 ),
    .fx({\u2_Display/n2735 [22],\u2_Display/n2735 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u23_al_u4885  (
    .a({\u2_Display/n2707 ,\u2_Display/n2709 }),
    .b({\u2_Display/n2706 ,\u2_Display/n2708 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b00),
    .fci(\u2_Display/add86/c23 ),
    .f({\u2_Display/n2735 [25],\u2_Display/n2735 [23]}),
    .fco(\u2_Display/add86/c27 ),
    .fx({\u2_Display/n2735 [26],\u2_Display/n2735 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u27_al_u4886  (
    .a({\u2_Display/n2703 ,\u2_Display/n2705 }),
    .b({\u2_Display/n2702 ,\u2_Display/n2704 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add86/c27 ),
    .f({\u2_Display/n2735 [29],\u2_Display/n2735 [27]}),
    .fco(\u2_Display/add86/c31 ),
    .fx({\u2_Display/n2735 [30],\u2_Display/n2735 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u31_al_u4887  (
    .a({open_n66924,\u2_Display/n2701 }),
    .c(2'b00),
    .d({open_n66929,1'b1}),
    .fci(\u2_Display/add86/c31 ),
    .f({open_n66946,\u2_Display/n2735 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u3_al_u4880  (
    .a({\u2_Display/n2727 ,\u2_Display/n2729 }),
    .b({\u2_Display/n2726 ,\u2_Display/n2728 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add86/c3 ),
    .f({\u2_Display/n2735 [5],\u2_Display/n2735 [3]}),
    .fco(\u2_Display/add86/c7 ),
    .fx({\u2_Display/n2735 [6],\u2_Display/n2735 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u7_al_u4881  (
    .a({\u2_Display/n2723 ,\u2_Display/n2725 }),
    .b({\u2_Display/n2722 ,\u2_Display/n2724 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add86/c7 ),
    .f({\u2_Display/n2735 [9],\u2_Display/n2735 [7]}),
    .fco(\u2_Display/add86/c11 ),
    .fx({\u2_Display/n2735 [10],\u2_Display/n2735 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/ucin_al_u4879  (
    .a({\u2_Display/n2731 ,1'b1}),
    .b({\u2_Display/n2730 ,\u2_Display/n2732 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2735 [1],open_n67005}),
    .fco(\u2_Display/add86/c3 ),
    .fx({\u2_Display/n2735 [2],\u2_Display/n2735 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u11_al_u4891  (
    .a({\u2_Display/n2754 ,\u2_Display/n2756 }),
    .b({\u2_Display/n2753 ,\u2_Display/n2755 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add87/c11 ),
    .f({\u2_Display/n2770 [13],\u2_Display/n2770 [11]}),
    .fco(\u2_Display/add87/c15 ),
    .fx({\u2_Display/n2770 [14],\u2_Display/n2770 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u15_al_u4892  (
    .a({\u2_Display/n2750 ,\u2_Display/n2752 }),
    .b({\u2_Display/n2749 ,\u2_Display/n2751 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add87/c15 ),
    .f({\u2_Display/n2770 [17],\u2_Display/n2770 [15]}),
    .fco(\u2_Display/add87/c19 ),
    .fx({\u2_Display/n2770 [18],\u2_Display/n2770 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u19_al_u4893  (
    .a({\u2_Display/n2746 ,\u2_Display/n2748 }),
    .b({\u2_Display/n2745 ,\u2_Display/n2747 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add87/c19 ),
    .f({\u2_Display/n2770 [21],\u2_Display/n2770 [19]}),
    .fco(\u2_Display/add87/c23 ),
    .fx({\u2_Display/n2770 [22],\u2_Display/n2770 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u23_al_u4894  (
    .a({\u2_Display/n2742 ,\u2_Display/n2744 }),
    .b({\u2_Display/n2741 ,\u2_Display/n2743 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add87/c23 ),
    .f({\u2_Display/n2770 [25],\u2_Display/n2770 [23]}),
    .fco(\u2_Display/add87/c27 ),
    .fx({\u2_Display/n2770 [26],\u2_Display/n2770 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u27_al_u4895  (
    .a({\u2_Display/n2738 ,\u2_Display/n2740 }),
    .b({\u2_Display/n2737 ,\u2_Display/n2739 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add87/c27 ),
    .f({\u2_Display/n2770 [29],\u2_Display/n2770 [27]}),
    .fco(\u2_Display/add87/c31 ),
    .fx({\u2_Display/n2770 [30],\u2_Display/n2770 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u31_al_u4896  (
    .a({open_n67098,\u2_Display/n2736 }),
    .c(2'b00),
    .d({open_n67103,1'b1}),
    .fci(\u2_Display/add87/c31 ),
    .f({open_n67120,\u2_Display/n2770 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u3_al_u4889  (
    .a({\u2_Display/n2762 ,\u2_Display/n2764 }),
    .b({\u2_Display/n2761 ,\u2_Display/n2763 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add87/c3 ),
    .f({\u2_Display/n2770 [5],\u2_Display/n2770 [3]}),
    .fco(\u2_Display/add87/c7 ),
    .fx({\u2_Display/n2770 [6],\u2_Display/n2770 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u7_al_u4890  (
    .a({\u2_Display/n2758 ,\u2_Display/n2760 }),
    .b({\u2_Display/n2757 ,\u2_Display/n2759 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add87/c7 ),
    .f({\u2_Display/n2770 [9],\u2_Display/n2770 [7]}),
    .fco(\u2_Display/add87/c11 ),
    .fx({\u2_Display/n2770 [10],\u2_Display/n2770 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/ucin_al_u4888  (
    .a({\u2_Display/n2766 ,1'b1}),
    .b({\u2_Display/n2765 ,\u2_Display/n2767 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2770 [1],open_n67179}),
    .fco(\u2_Display/add87/c3 ),
    .fx({\u2_Display/n2770 [2],\u2_Display/n2770 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u11_al_u4900  (
    .a({\u2_Display/n2789 ,\u2_Display/n2791 }),
    .b({\u2_Display/n2788 ,\u2_Display/n2790 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add88/c11 ),
    .f({\u2_Display/n2805 [13],\u2_Display/n2805 [11]}),
    .fco(\u2_Display/add88/c15 ),
    .fx({\u2_Display/n2805 [14],\u2_Display/n2805 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u15_al_u4901  (
    .a({\u2_Display/n2785 ,\u2_Display/n2787 }),
    .b({\u2_Display/n2784 ,\u2_Display/n2786 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add88/c15 ),
    .f({\u2_Display/n2805 [17],\u2_Display/n2805 [15]}),
    .fco(\u2_Display/add88/c19 ),
    .fx({\u2_Display/n2805 [18],\u2_Display/n2805 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u19_al_u4902  (
    .a({\u2_Display/n2781 ,\u2_Display/n2783 }),
    .b({\u2_Display/n2780 ,\u2_Display/n2782 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add88/c19 ),
    .f({\u2_Display/n2805 [21],\u2_Display/n2805 [19]}),
    .fco(\u2_Display/add88/c23 ),
    .fx({\u2_Display/n2805 [22],\u2_Display/n2805 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u23_al_u4903  (
    .a({\u2_Display/n2777 ,\u2_Display/n2779 }),
    .b({\u2_Display/n2776 ,\u2_Display/n2778 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add88/c23 ),
    .f({\u2_Display/n2805 [25],\u2_Display/n2805 [23]}),
    .fco(\u2_Display/add88/c27 ),
    .fx({\u2_Display/n2805 [26],\u2_Display/n2805 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u27_al_u4904  (
    .a({\u2_Display/n2773 ,\u2_Display/n2775 }),
    .b({\u2_Display/n2772 ,\u2_Display/n2774 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add88/c27 ),
    .f({\u2_Display/n2805 [29],\u2_Display/n2805 [27]}),
    .fco(\u2_Display/add88/c31 ),
    .fx({\u2_Display/n2805 [30],\u2_Display/n2805 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u31_al_u4905  (
    .a({open_n67272,\u2_Display/n2771 }),
    .c(2'b00),
    .d({open_n67277,1'b1}),
    .fci(\u2_Display/add88/c31 ),
    .f({open_n67294,\u2_Display/n2805 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u3_al_u4898  (
    .a({\u2_Display/n2797 ,\u2_Display/n2799 }),
    .b({\u2_Display/n2796 ,\u2_Display/n2798 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add88/c3 ),
    .f({\u2_Display/n2805 [5],\u2_Display/n2805 [3]}),
    .fco(\u2_Display/add88/c7 ),
    .fx({\u2_Display/n2805 [6],\u2_Display/n2805 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u7_al_u4899  (
    .a({\u2_Display/n2793 ,\u2_Display/n2795 }),
    .b({\u2_Display/n2792 ,\u2_Display/n2794 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add88/c7 ),
    .f({\u2_Display/n2805 [9],\u2_Display/n2805 [7]}),
    .fco(\u2_Display/add88/c11 ),
    .fx({\u2_Display/n2805 [10],\u2_Display/n2805 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/ucin_al_u4897  (
    .a({\u2_Display/n2801 ,1'b1}),
    .b({\u2_Display/n2800 ,\u2_Display/n2802 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2805 [1],open_n67353}),
    .fco(\u2_Display/add88/c3 ),
    .fx({\u2_Display/n2805 [2],\u2_Display/n2805 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u11_al_u4909  (
    .a({\u2_Display/n2824 ,\u2_Display/n2826 }),
    .b({\u2_Display/n2823 ,\u2_Display/n2825 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add89/c11 ),
    .f({\u2_Display/n2840 [13],\u2_Display/n2840 [11]}),
    .fco(\u2_Display/add89/c15 ),
    .fx({\u2_Display/n2840 [14],\u2_Display/n2840 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u15_al_u4910  (
    .a({\u2_Display/n2820 ,\u2_Display/n2822 }),
    .b({\u2_Display/n2819 ,\u2_Display/n2821 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add89/c15 ),
    .f({\u2_Display/n2840 [17],\u2_Display/n2840 [15]}),
    .fco(\u2_Display/add89/c19 ),
    .fx({\u2_Display/n2840 [18],\u2_Display/n2840 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u19_al_u4911  (
    .a({\u2_Display/n2816 ,\u2_Display/n2818 }),
    .b({\u2_Display/n2815 ,\u2_Display/n2817 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add89/c19 ),
    .f({\u2_Display/n2840 [21],\u2_Display/n2840 [19]}),
    .fco(\u2_Display/add89/c23 ),
    .fx({\u2_Display/n2840 [22],\u2_Display/n2840 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u23_al_u4912  (
    .a({\u2_Display/n2812 ,\u2_Display/n2814 }),
    .b({\u2_Display/n2811 ,\u2_Display/n2813 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add89/c23 ),
    .f({\u2_Display/n2840 [25],\u2_Display/n2840 [23]}),
    .fco(\u2_Display/add89/c27 ),
    .fx({\u2_Display/n2840 [26],\u2_Display/n2840 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u27_al_u4913  (
    .a({\u2_Display/n2808 ,\u2_Display/n2810 }),
    .b({\u2_Display/n2807 ,\u2_Display/n2809 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add89/c27 ),
    .f({\u2_Display/n2840 [29],\u2_Display/n2840 [27]}),
    .fco(\u2_Display/add89/c31 ),
    .fx({\u2_Display/n2840 [30],\u2_Display/n2840 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u31_al_u4914  (
    .a({open_n67446,\u2_Display/n2806 }),
    .c(2'b00),
    .d({open_n67451,1'b1}),
    .fci(\u2_Display/add89/c31 ),
    .f({open_n67468,\u2_Display/n2840 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u3_al_u4907  (
    .a({\u2_Display/n2832 ,\u2_Display/n2834 }),
    .b({\u2_Display/n2831 ,\u2_Display/n2833 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add89/c3 ),
    .f({\u2_Display/n2840 [5],\u2_Display/n2840 [3]}),
    .fco(\u2_Display/add89/c7 ),
    .fx({\u2_Display/n2840 [6],\u2_Display/n2840 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u7_al_u4908  (
    .a({\u2_Display/n2828 ,\u2_Display/n2830 }),
    .b({\u2_Display/n2827 ,\u2_Display/n2829 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add89/c7 ),
    .f({\u2_Display/n2840 [9],\u2_Display/n2840 [7]}),
    .fco(\u2_Display/add89/c11 ),
    .fx({\u2_Display/n2840 [10],\u2_Display/n2840 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/ucin_al_u4906  (
    .a({\u2_Display/n2836 ,1'b1}),
    .b({\u2_Display/n2835 ,\u2_Display/n2837 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2840 [1],open_n67527}),
    .fco(\u2_Display/add89/c3 ),
    .fx({\u2_Display/n2840 [2],\u2_Display/n2840 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u11_al_u4918  (
    .a({\u2_Display/n2859 ,\u2_Display/n2861 }),
    .b({\u2_Display/n2858 ,\u2_Display/n2860 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add90/c11 ),
    .f({\u2_Display/n2875 [13],\u2_Display/n2875 [11]}),
    .fco(\u2_Display/add90/c15 ),
    .fx({\u2_Display/n2875 [14],\u2_Display/n2875 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u15_al_u4919  (
    .a({\u2_Display/n2855 ,\u2_Display/n2857 }),
    .b({\u2_Display/n2854 ,\u2_Display/n2856 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add90/c15 ),
    .f({\u2_Display/n2875 [17],\u2_Display/n2875 [15]}),
    .fco(\u2_Display/add90/c19 ),
    .fx({\u2_Display/n2875 [18],\u2_Display/n2875 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u19_al_u4920  (
    .a({\u2_Display/n2851 ,\u2_Display/n2853 }),
    .b({\u2_Display/n2850 ,\u2_Display/n2852 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b00),
    .fci(\u2_Display/add90/c19 ),
    .f({\u2_Display/n2875 [21],\u2_Display/n2875 [19]}),
    .fco(\u2_Display/add90/c23 ),
    .fx({\u2_Display/n2875 [22],\u2_Display/n2875 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u23_al_u4921  (
    .a({\u2_Display/n2847 ,\u2_Display/n2849 }),
    .b({\u2_Display/n2846 ,\u2_Display/n2848 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add90/c23 ),
    .f({\u2_Display/n2875 [25],\u2_Display/n2875 [23]}),
    .fco(\u2_Display/add90/c27 ),
    .fx({\u2_Display/n2875 [26],\u2_Display/n2875 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u27_al_u4922  (
    .a({\u2_Display/n2843 ,\u2_Display/n2845 }),
    .b({\u2_Display/n2842 ,\u2_Display/n2844 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add90/c27 ),
    .f({\u2_Display/n2875 [29],\u2_Display/n2875 [27]}),
    .fco(\u2_Display/add90/c31 ),
    .fx({\u2_Display/n2875 [30],\u2_Display/n2875 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u31_al_u4923  (
    .a({open_n67620,\u2_Display/n2841 }),
    .c(2'b00),
    .d({open_n67625,1'b1}),
    .fci(\u2_Display/add90/c31 ),
    .f({open_n67642,\u2_Display/n2875 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u3_al_u4916  (
    .a({\u2_Display/n2867 ,\u2_Display/n2869 }),
    .b({\u2_Display/n2866 ,\u2_Display/n2868 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add90/c3 ),
    .f({\u2_Display/n2875 [5],\u2_Display/n2875 [3]}),
    .fco(\u2_Display/add90/c7 ),
    .fx({\u2_Display/n2875 [6],\u2_Display/n2875 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u7_al_u4917  (
    .a({\u2_Display/n2863 ,\u2_Display/n2865 }),
    .b({\u2_Display/n2862 ,\u2_Display/n2864 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add90/c7 ),
    .f({\u2_Display/n2875 [9],\u2_Display/n2875 [7]}),
    .fco(\u2_Display/add90/c11 ),
    .fx({\u2_Display/n2875 [10],\u2_Display/n2875 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/ucin_al_u4915  (
    .a({\u2_Display/n2871 ,1'b1}),
    .b({\u2_Display/n2870 ,\u2_Display/n2872 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2875 [1],open_n67701}),
    .fco(\u2_Display/add90/c3 ),
    .fx({\u2_Display/n2875 [2],\u2_Display/n2875 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u11_al_u4927  (
    .a({\u2_Display/n2894 ,\u2_Display/n2896 }),
    .b({\u2_Display/n2893 ,\u2_Display/n2895 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add91/c11 ),
    .f({\u2_Display/n2910 [13],\u2_Display/n2910 [11]}),
    .fco(\u2_Display/add91/c15 ),
    .fx({\u2_Display/n2910 [14],\u2_Display/n2910 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u15_al_u4928  (
    .a({\u2_Display/n2890 ,\u2_Display/n2892 }),
    .b({\u2_Display/n2889 ,\u2_Display/n2891 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add91/c15 ),
    .f({\u2_Display/n2910 [17],\u2_Display/n2910 [15]}),
    .fco(\u2_Display/add91/c19 ),
    .fx({\u2_Display/n2910 [18],\u2_Display/n2910 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u19_al_u4929  (
    .a({\u2_Display/n2886 ,\u2_Display/n2888 }),
    .b({\u2_Display/n2885 ,\u2_Display/n2887 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add91/c19 ),
    .f({\u2_Display/n2910 [21],\u2_Display/n2910 [19]}),
    .fco(\u2_Display/add91/c23 ),
    .fx({\u2_Display/n2910 [22],\u2_Display/n2910 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u23_al_u4930  (
    .a({\u2_Display/n2882 ,\u2_Display/n2884 }),
    .b({\u2_Display/n2881 ,\u2_Display/n2883 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add91/c23 ),
    .f({\u2_Display/n2910 [25],\u2_Display/n2910 [23]}),
    .fco(\u2_Display/add91/c27 ),
    .fx({\u2_Display/n2910 [26],\u2_Display/n2910 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u27_al_u4931  (
    .a({\u2_Display/n2878 ,\u2_Display/n2880 }),
    .b({\u2_Display/n2877 ,\u2_Display/n2879 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add91/c27 ),
    .f({\u2_Display/n2910 [29],\u2_Display/n2910 [27]}),
    .fco(\u2_Display/add91/c31 ),
    .fx({\u2_Display/n2910 [30],\u2_Display/n2910 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u31_al_u4932  (
    .a({open_n67794,\u2_Display/n2876 }),
    .c(2'b00),
    .d({open_n67799,1'b1}),
    .fci(\u2_Display/add91/c31 ),
    .f({open_n67816,\u2_Display/n2910 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u3_al_u4925  (
    .a({\u2_Display/n2902 ,\u2_Display/n2904 }),
    .b({\u2_Display/n2901 ,\u2_Display/n2903 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add91/c3 ),
    .f({\u2_Display/n2910 [5],\u2_Display/n2910 [3]}),
    .fco(\u2_Display/add91/c7 ),
    .fx({\u2_Display/n2910 [6],\u2_Display/n2910 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u7_al_u4926  (
    .a({\u2_Display/n2898 ,\u2_Display/n2900 }),
    .b({\u2_Display/n2897 ,\u2_Display/n2899 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add91/c7 ),
    .f({\u2_Display/n2910 [9],\u2_Display/n2910 [7]}),
    .fco(\u2_Display/add91/c11 ),
    .fx({\u2_Display/n2910 [10],\u2_Display/n2910 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/ucin_al_u4924  (
    .a({\u2_Display/n2906 ,1'b1}),
    .b({\u2_Display/n2905 ,\u2_Display/n2907 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2910 [1],open_n67875}),
    .fco(\u2_Display/add91/c3 ),
    .fx({\u2_Display/n2910 [2],\u2_Display/n2910 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u11_al_u4936  (
    .a({\u2_Display/n2929 ,\u2_Display/n2931 }),
    .b({\u2_Display/n2928 ,\u2_Display/n2930 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add92/c11 ),
    .f({\u2_Display/n2945 [13],\u2_Display/n2945 [11]}),
    .fco(\u2_Display/add92/c15 ),
    .fx({\u2_Display/n2945 [14],\u2_Display/n2945 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u15_al_u4937  (
    .a({\u2_Display/n2925 ,\u2_Display/n2927 }),
    .b({\u2_Display/n2924 ,\u2_Display/n2926 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add92/c15 ),
    .f({\u2_Display/n2945 [17],\u2_Display/n2945 [15]}),
    .fco(\u2_Display/add92/c19 ),
    .fx({\u2_Display/n2945 [18],\u2_Display/n2945 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u19_al_u4938  (
    .a({\u2_Display/n2921 ,\u2_Display/n2923 }),
    .b({\u2_Display/n2920 ,\u2_Display/n2922 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add92/c19 ),
    .f({\u2_Display/n2945 [21],\u2_Display/n2945 [19]}),
    .fco(\u2_Display/add92/c23 ),
    .fx({\u2_Display/n2945 [22],\u2_Display/n2945 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u23_al_u4939  (
    .a({\u2_Display/n2917 ,\u2_Display/n2919 }),
    .b({\u2_Display/n2916 ,\u2_Display/n2918 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add92/c23 ),
    .f({\u2_Display/n2945 [25],\u2_Display/n2945 [23]}),
    .fco(\u2_Display/add92/c27 ),
    .fx({\u2_Display/n2945 [26],\u2_Display/n2945 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u27_al_u4940  (
    .a({\u2_Display/n2913 ,\u2_Display/n2915 }),
    .b({\u2_Display/n2912 ,\u2_Display/n2914 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add92/c27 ),
    .f({\u2_Display/n2945 [29],\u2_Display/n2945 [27]}),
    .fco(\u2_Display/add92/c31 ),
    .fx({\u2_Display/n2945 [30],\u2_Display/n2945 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u31_al_u4941  (
    .a({open_n67968,\u2_Display/n2911 }),
    .c(2'b00),
    .d({open_n67973,1'b1}),
    .fci(\u2_Display/add92/c31 ),
    .f({open_n67990,\u2_Display/n2945 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u3_al_u4934  (
    .a({\u2_Display/n2937 ,\u2_Display/n2939 }),
    .b({\u2_Display/n2936 ,\u2_Display/n2938 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add92/c3 ),
    .f({\u2_Display/n2945 [5],\u2_Display/n2945 [3]}),
    .fco(\u2_Display/add92/c7 ),
    .fx({\u2_Display/n2945 [6],\u2_Display/n2945 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u7_al_u4935  (
    .a({\u2_Display/n2933 ,\u2_Display/n2935 }),
    .b({\u2_Display/n2932 ,\u2_Display/n2934 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add92/c7 ),
    .f({\u2_Display/n2945 [9],\u2_Display/n2945 [7]}),
    .fco(\u2_Display/add92/c11 ),
    .fx({\u2_Display/n2945 [10],\u2_Display/n2945 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/ucin_al_u4933  (
    .a({\u2_Display/n2941 ,1'b1}),
    .b({\u2_Display/n2940 ,\u2_Display/n2942 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2945 [1],open_n68049}),
    .fco(\u2_Display/add92/c3 ),
    .fx({\u2_Display/n2945 [2],\u2_Display/n2945 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u11_al_u4945  (
    .a({\u2_Display/n2964 ,\u2_Display/n2966 }),
    .b({\u2_Display/n2963 ,\u2_Display/n2965 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add93/c11 ),
    .f({\u2_Display/n2980 [13],\u2_Display/n2980 [11]}),
    .fco(\u2_Display/add93/c15 ),
    .fx({\u2_Display/n2980 [14],\u2_Display/n2980 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u15_al_u4946  (
    .a({\u2_Display/n2960 ,\u2_Display/n2962 }),
    .b({\u2_Display/n2959 ,\u2_Display/n2961 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add93/c15 ),
    .f({\u2_Display/n2980 [17],\u2_Display/n2980 [15]}),
    .fco(\u2_Display/add93/c19 ),
    .fx({\u2_Display/n2980 [18],\u2_Display/n2980 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u19_al_u4947  (
    .a({\u2_Display/n2956 ,\u2_Display/n2958 }),
    .b({\u2_Display/n2955 ,\u2_Display/n2957 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add93/c19 ),
    .f({\u2_Display/n2980 [21],\u2_Display/n2980 [19]}),
    .fco(\u2_Display/add93/c23 ),
    .fx({\u2_Display/n2980 [22],\u2_Display/n2980 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u23_al_u4948  (
    .a({\u2_Display/n2952 ,\u2_Display/n2954 }),
    .b({\u2_Display/n2951 ,\u2_Display/n2953 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add93/c23 ),
    .f({\u2_Display/n2980 [25],\u2_Display/n2980 [23]}),
    .fco(\u2_Display/add93/c27 ),
    .fx({\u2_Display/n2980 [26],\u2_Display/n2980 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u27_al_u4949  (
    .a({\u2_Display/n2948 ,\u2_Display/n2950 }),
    .b({\u2_Display/n2947 ,\u2_Display/n2949 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add93/c27 ),
    .f({\u2_Display/n2980 [29],\u2_Display/n2980 [27]}),
    .fco(\u2_Display/add93/c31 ),
    .fx({\u2_Display/n2980 [30],\u2_Display/n2980 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u31_al_u4950  (
    .a({open_n68142,\u2_Display/n2946 }),
    .c(2'b00),
    .d({open_n68147,1'b1}),
    .fci(\u2_Display/add93/c31 ),
    .f({open_n68164,\u2_Display/n2980 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u3_al_u4943  (
    .a({\u2_Display/n2972 ,\u2_Display/n2974 }),
    .b({\u2_Display/n2971 ,\u2_Display/n2973 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add93/c3 ),
    .f({\u2_Display/n2980 [5],\u2_Display/n2980 [3]}),
    .fco(\u2_Display/add93/c7 ),
    .fx({\u2_Display/n2980 [6],\u2_Display/n2980 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u7_al_u4944  (
    .a({\u2_Display/n2968 ,\u2_Display/n2970 }),
    .b({\u2_Display/n2967 ,\u2_Display/n2969 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add93/c7 ),
    .f({\u2_Display/n2980 [9],\u2_Display/n2980 [7]}),
    .fco(\u2_Display/add93/c11 ),
    .fx({\u2_Display/n2980 [10],\u2_Display/n2980 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/ucin_al_u4942  (
    .a({\u2_Display/n2976 ,1'b1}),
    .b({\u2_Display/n2975 ,\u2_Display/n2977 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2980 [1],open_n68223}),
    .fco(\u2_Display/add93/c3 ),
    .fx({\u2_Display/n2980 [2],\u2_Display/n2980 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u11_al_u4954  (
    .a({\u2_Display/n2999 ,\u2_Display/n3001 }),
    .b({\u2_Display/n2998 ,\u2_Display/n3000 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add94/c11 ),
    .f({\u2_Display/n3015 [13],\u2_Display/n3015 [11]}),
    .fco(\u2_Display/add94/c15 ),
    .fx({\u2_Display/n3015 [14],\u2_Display/n3015 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u15_al_u4955  (
    .a({\u2_Display/n2995 ,\u2_Display/n2997 }),
    .b({\u2_Display/n2994 ,\u2_Display/n2996 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b00),
    .fci(\u2_Display/add94/c15 ),
    .f({\u2_Display/n3015 [17],\u2_Display/n3015 [15]}),
    .fco(\u2_Display/add94/c19 ),
    .fx({\u2_Display/n3015 [18],\u2_Display/n3015 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u19_al_u4956  (
    .a({\u2_Display/n2991 ,\u2_Display/n2993 }),
    .b({\u2_Display/n2990 ,\u2_Display/n2992 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add94/c19 ),
    .f({\u2_Display/n3015 [21],\u2_Display/n3015 [19]}),
    .fco(\u2_Display/add94/c23 ),
    .fx({\u2_Display/n3015 [22],\u2_Display/n3015 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u23_al_u4957  (
    .a({\u2_Display/n2987 ,\u2_Display/n2989 }),
    .b({\u2_Display/n2986 ,\u2_Display/n2988 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add94/c23 ),
    .f({\u2_Display/n3015 [25],\u2_Display/n3015 [23]}),
    .fco(\u2_Display/add94/c27 ),
    .fx({\u2_Display/n3015 [26],\u2_Display/n3015 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u27_al_u4958  (
    .a({\u2_Display/n2983 ,\u2_Display/n2985 }),
    .b({\u2_Display/n2982 ,\u2_Display/n2984 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add94/c27 ),
    .f({\u2_Display/n3015 [29],\u2_Display/n3015 [27]}),
    .fco(\u2_Display/add94/c31 ),
    .fx({\u2_Display/n3015 [30],\u2_Display/n3015 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u31_al_u4959  (
    .a({open_n68316,\u2_Display/n2981 }),
    .c(2'b00),
    .d({open_n68321,1'b1}),
    .fci(\u2_Display/add94/c31 ),
    .f({open_n68338,\u2_Display/n3015 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u3_al_u4952  (
    .a({\u2_Display/n3007 ,\u2_Display/n3009 }),
    .b({\u2_Display/n3006 ,\u2_Display/n3008 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add94/c3 ),
    .f({\u2_Display/n3015 [5],\u2_Display/n3015 [3]}),
    .fco(\u2_Display/add94/c7 ),
    .fx({\u2_Display/n3015 [6],\u2_Display/n3015 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u7_al_u4953  (
    .a({\u2_Display/n3003 ,\u2_Display/n3005 }),
    .b({\u2_Display/n3002 ,\u2_Display/n3004 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add94/c7 ),
    .f({\u2_Display/n3015 [9],\u2_Display/n3015 [7]}),
    .fco(\u2_Display/add94/c11 ),
    .fx({\u2_Display/n3015 [10],\u2_Display/n3015 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/ucin_al_u4951  (
    .a({\u2_Display/n3011 ,1'b1}),
    .b({\u2_Display/n3010 ,\u2_Display/n3012 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3015 [1],open_n68397}),
    .fco(\u2_Display/add94/c3 ),
    .fx({\u2_Display/n3015 [2],\u2_Display/n3015 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u11_al_u4963  (
    .a({\u2_Display/n3034 ,\u2_Display/n3036 }),
    .b({\u2_Display/n3033 ,\u2_Display/n3035 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add95/c11 ),
    .f({\u2_Display/n3050 [13],\u2_Display/n3050 [11]}),
    .fco(\u2_Display/add95/c15 ),
    .fx({\u2_Display/n3050 [14],\u2_Display/n3050 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u15_al_u4964  (
    .a({\u2_Display/n3030 ,\u2_Display/n3032 }),
    .b({\u2_Display/n3029 ,\u2_Display/n3031 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add95/c15 ),
    .f({\u2_Display/n3050 [17],\u2_Display/n3050 [15]}),
    .fco(\u2_Display/add95/c19 ),
    .fx({\u2_Display/n3050 [18],\u2_Display/n3050 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u19_al_u4965  (
    .a({\u2_Display/n3026 ,\u2_Display/n3028 }),
    .b({\u2_Display/n3025 ,\u2_Display/n3027 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add95/c19 ),
    .f({\u2_Display/n3050 [21],\u2_Display/n3050 [19]}),
    .fco(\u2_Display/add95/c23 ),
    .fx({\u2_Display/n3050 [22],\u2_Display/n3050 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u23_al_u4966  (
    .a({\u2_Display/n3022 ,\u2_Display/n3024 }),
    .b({\u2_Display/n3021 ,\u2_Display/n3023 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add95/c23 ),
    .f({\u2_Display/n3050 [25],\u2_Display/n3050 [23]}),
    .fco(\u2_Display/add95/c27 ),
    .fx({\u2_Display/n3050 [26],\u2_Display/n3050 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u27_al_u4967  (
    .a({\u2_Display/n3018 ,\u2_Display/n3020 }),
    .b({\u2_Display/n3017 ,\u2_Display/n3019 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add95/c27 ),
    .f({\u2_Display/n3050 [29],\u2_Display/n3050 [27]}),
    .fco(\u2_Display/add95/c31 ),
    .fx({\u2_Display/n3050 [30],\u2_Display/n3050 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u31_al_u4968  (
    .a({open_n68490,\u2_Display/n3016 }),
    .c(2'b00),
    .d({open_n68495,1'b1}),
    .fci(\u2_Display/add95/c31 ),
    .f({open_n68512,\u2_Display/n3050 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u3_al_u4961  (
    .a({\u2_Display/n3042 ,\u2_Display/n3044 }),
    .b({\u2_Display/n3041 ,\u2_Display/n3043 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add95/c3 ),
    .f({\u2_Display/n3050 [5],\u2_Display/n3050 [3]}),
    .fco(\u2_Display/add95/c7 ),
    .fx({\u2_Display/n3050 [6],\u2_Display/n3050 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u7_al_u4962  (
    .a({\u2_Display/n3038 ,\u2_Display/n3040 }),
    .b({\u2_Display/n3037 ,\u2_Display/n3039 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add95/c7 ),
    .f({\u2_Display/n3050 [9],\u2_Display/n3050 [7]}),
    .fco(\u2_Display/add95/c11 ),
    .fx({\u2_Display/n3050 [10],\u2_Display/n3050 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/ucin_al_u4960  (
    .a({\u2_Display/n3046 ,1'b1}),
    .b({\u2_Display/n3045 ,\u2_Display/n3047 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3050 [1],open_n68571}),
    .fco(\u2_Display/add95/c3 ),
    .fx({\u2_Display/n3050 [2],\u2_Display/n3050 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u11_al_u4972  (
    .a({\u2_Display/n3069 ,\u2_Display/n3071 }),
    .b({\u2_Display/n3068 ,\u2_Display/n3070 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add96/c11 ),
    .f({\u2_Display/n3085 [13],\u2_Display/n3085 [11]}),
    .fco(\u2_Display/add96/c15 ),
    .fx({\u2_Display/n3085 [14],\u2_Display/n3085 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u15_al_u4973  (
    .a({\u2_Display/n3065 ,\u2_Display/n3067 }),
    .b({\u2_Display/n3064 ,\u2_Display/n3066 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add96/c15 ),
    .f({\u2_Display/n3085 [17],\u2_Display/n3085 [15]}),
    .fco(\u2_Display/add96/c19 ),
    .fx({\u2_Display/n3085 [18],\u2_Display/n3085 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u19_al_u4974  (
    .a({\u2_Display/n3061 ,\u2_Display/n3063 }),
    .b({\u2_Display/n3060 ,\u2_Display/n3062 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add96/c19 ),
    .f({\u2_Display/n3085 [21],\u2_Display/n3085 [19]}),
    .fco(\u2_Display/add96/c23 ),
    .fx({\u2_Display/n3085 [22],\u2_Display/n3085 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u23_al_u4975  (
    .a({\u2_Display/n3057 ,\u2_Display/n3059 }),
    .b({\u2_Display/n3056 ,\u2_Display/n3058 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add96/c23 ),
    .f({\u2_Display/n3085 [25],\u2_Display/n3085 [23]}),
    .fco(\u2_Display/add96/c27 ),
    .fx({\u2_Display/n3085 [26],\u2_Display/n3085 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u27_al_u4976  (
    .a({\u2_Display/n3053 ,\u2_Display/n3055 }),
    .b({\u2_Display/n3052 ,\u2_Display/n3054 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add96/c27 ),
    .f({\u2_Display/n3085 [29],\u2_Display/n3085 [27]}),
    .fco(\u2_Display/add96/c31 ),
    .fx({\u2_Display/n3085 [30],\u2_Display/n3085 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u31_al_u4977  (
    .a({open_n68664,\u2_Display/n3051 }),
    .c(2'b00),
    .d({open_n68669,1'b1}),
    .fci(\u2_Display/add96/c31 ),
    .f({open_n68686,\u2_Display/n3085 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u3_al_u4970  (
    .a({\u2_Display/n3077 ,\u2_Display/n3079 }),
    .b({\u2_Display/n3076 ,\u2_Display/n3078 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add96/c3 ),
    .f({\u2_Display/n3085 [5],\u2_Display/n3085 [3]}),
    .fco(\u2_Display/add96/c7 ),
    .fx({\u2_Display/n3085 [6],\u2_Display/n3085 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u7_al_u4971  (
    .a({\u2_Display/n3073 ,\u2_Display/n3075 }),
    .b({\u2_Display/n3072 ,\u2_Display/n3074 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add96/c7 ),
    .f({\u2_Display/n3085 [9],\u2_Display/n3085 [7]}),
    .fco(\u2_Display/add96/c11 ),
    .fx({\u2_Display/n3085 [10],\u2_Display/n3085 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/ucin_al_u4969  (
    .a({\u2_Display/n3081 ,1'b1}),
    .b({\u2_Display/n3080 ,\u2_Display/n3082 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3085 [1],open_n68745}),
    .fco(\u2_Display/add96/c3 ),
    .fx({\u2_Display/n3085 [2],\u2_Display/n3085 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u11_al_u4981  (
    .a({\u2_Display/n3104 ,\u2_Display/n3106 }),
    .b({\u2_Display/n3103 ,\u2_Display/n3105 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add97/c11 ),
    .f({\u2_Display/n3120 [13],\u2_Display/n3120 [11]}),
    .fco(\u2_Display/add97/c15 ),
    .fx({\u2_Display/n3120 [14],\u2_Display/n3120 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u15_al_u4982  (
    .a({\u2_Display/n3100 ,\u2_Display/n3102 }),
    .b({\u2_Display/n3099 ,\u2_Display/n3101 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add97/c15 ),
    .f({\u2_Display/n3120 [17],\u2_Display/n3120 [15]}),
    .fco(\u2_Display/add97/c19 ),
    .fx({\u2_Display/n3120 [18],\u2_Display/n3120 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u19_al_u4983  (
    .a({\u2_Display/n3096 ,\u2_Display/n3098 }),
    .b({\u2_Display/n3095 ,\u2_Display/n3097 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add97/c19 ),
    .f({\u2_Display/n3120 [21],\u2_Display/n3120 [19]}),
    .fco(\u2_Display/add97/c23 ),
    .fx({\u2_Display/n3120 [22],\u2_Display/n3120 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u23_al_u4984  (
    .a({\u2_Display/n3092 ,\u2_Display/n3094 }),
    .b({\u2_Display/n3091 ,\u2_Display/n3093 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add97/c23 ),
    .f({\u2_Display/n3120 [25],\u2_Display/n3120 [23]}),
    .fco(\u2_Display/add97/c27 ),
    .fx({\u2_Display/n3120 [26],\u2_Display/n3120 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u27_al_u4985  (
    .a({\u2_Display/n3088 ,\u2_Display/n3090 }),
    .b({\u2_Display/n3087 ,\u2_Display/n3089 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add97/c27 ),
    .f({\u2_Display/n3120 [29],\u2_Display/n3120 [27]}),
    .fco(\u2_Display/add97/c31 ),
    .fx({\u2_Display/n3120 [30],\u2_Display/n3120 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u31_al_u4986  (
    .a({open_n68838,\u2_Display/n3086 }),
    .c(2'b00),
    .d({open_n68843,1'b1}),
    .fci(\u2_Display/add97/c31 ),
    .f({open_n68860,\u2_Display/n3120 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u3_al_u4979  (
    .a({\u2_Display/n3112 ,\u2_Display/n3114 }),
    .b({\u2_Display/n3111 ,\u2_Display/n3113 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add97/c3 ),
    .f({\u2_Display/n3120 [5],\u2_Display/n3120 [3]}),
    .fco(\u2_Display/add97/c7 ),
    .fx({\u2_Display/n3120 [6],\u2_Display/n3120 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u7_al_u4980  (
    .a({\u2_Display/n3108 ,\u2_Display/n3110 }),
    .b({\u2_Display/n3107 ,\u2_Display/n3109 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add97/c7 ),
    .f({\u2_Display/n3120 [9],\u2_Display/n3120 [7]}),
    .fco(\u2_Display/add97/c11 ),
    .fx({\u2_Display/n3120 [10],\u2_Display/n3120 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/ucin_al_u4978  (
    .a({\u2_Display/n3116 ,1'b1}),
    .b({\u2_Display/n3115 ,\u2_Display/n3117 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3120 [1],open_n68919}),
    .fco(\u2_Display/add97/c3 ),
    .fx({\u2_Display/n3120 [2],\u2_Display/n3120 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u11_al_u4990  (
    .a({\u2_Display/n3139 ,\u2_Display/n3141 }),
    .b({\u2_Display/n3138 ,\u2_Display/n3140 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b00),
    .fci(\u2_Display/add98/c11 ),
    .f({\u2_Display/n3155 [13],\u2_Display/n3155 [11]}),
    .fco(\u2_Display/add98/c15 ),
    .fx({\u2_Display/n3155 [14],\u2_Display/n3155 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u15_al_u4991  (
    .a({\u2_Display/n3135 ,\u2_Display/n3137 }),
    .b({\u2_Display/n3134 ,\u2_Display/n3136 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add98/c15 ),
    .f({\u2_Display/n3155 [17],\u2_Display/n3155 [15]}),
    .fco(\u2_Display/add98/c19 ),
    .fx({\u2_Display/n3155 [18],\u2_Display/n3155 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u19_al_u4992  (
    .a({\u2_Display/n3131 ,\u2_Display/n3133 }),
    .b({\u2_Display/n3130 ,\u2_Display/n3132 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add98/c19 ),
    .f({\u2_Display/n3155 [21],\u2_Display/n3155 [19]}),
    .fco(\u2_Display/add98/c23 ),
    .fx({\u2_Display/n3155 [22],\u2_Display/n3155 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u23_al_u4993  (
    .a({\u2_Display/n3127 ,\u2_Display/n3129 }),
    .b({\u2_Display/n3126 ,\u2_Display/n3128 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add98/c23 ),
    .f({\u2_Display/n3155 [25],\u2_Display/n3155 [23]}),
    .fco(\u2_Display/add98/c27 ),
    .fx({\u2_Display/n3155 [26],\u2_Display/n3155 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u27_al_u4994  (
    .a({\u2_Display/n3123 ,\u2_Display/n3125 }),
    .b({\u2_Display/n3122 ,\u2_Display/n3124 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add98/c27 ),
    .f({\u2_Display/n3155 [29],\u2_Display/n3155 [27]}),
    .fco(\u2_Display/add98/c31 ),
    .fx({\u2_Display/n3155 [30],\u2_Display/n3155 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u31_al_u4995  (
    .a({open_n69012,\u2_Display/n3121 }),
    .c(2'b00),
    .d({open_n69017,1'b1}),
    .fci(\u2_Display/add98/c31 ),
    .f({open_n69034,\u2_Display/n3155 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u3_al_u4988  (
    .a({\u2_Display/n3147 ,\u2_Display/n3149 }),
    .b({\u2_Display/n3146 ,\u2_Display/n3148 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add98/c3 ),
    .f({\u2_Display/n3155 [5],\u2_Display/n3155 [3]}),
    .fco(\u2_Display/add98/c7 ),
    .fx({\u2_Display/n3155 [6],\u2_Display/n3155 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u7_al_u4989  (
    .a({\u2_Display/n3143 ,\u2_Display/n3145 }),
    .b({\u2_Display/n3142 ,\u2_Display/n3144 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add98/c7 ),
    .f({\u2_Display/n3155 [9],\u2_Display/n3155 [7]}),
    .fco(\u2_Display/add98/c11 ),
    .fx({\u2_Display/n3155 [10],\u2_Display/n3155 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/ucin_al_u4987  (
    .a({\u2_Display/n3151 ,1'b1}),
    .b({\u2_Display/n3150 ,\u2_Display/n3152 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3155 [1],open_n69093}),
    .fco(\u2_Display/add98/c3 ),
    .fx({\u2_Display/n3155 [2],\u2_Display/n3155 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u11_al_u4999  (
    .a({\u2_Display/n3174 ,\u2_Display/n3176 }),
    .b({\u2_Display/n3173 ,\u2_Display/n3175 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add99/c11 ),
    .f({\u2_Display/n3190 [13],\u2_Display/n3190 [11]}),
    .fco(\u2_Display/add99/c15 ),
    .fx({\u2_Display/n3190 [14],\u2_Display/n3190 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u15_al_u5000  (
    .a({\u2_Display/n3170 ,\u2_Display/n3172 }),
    .b({\u2_Display/n3169 ,\u2_Display/n3171 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add99/c15 ),
    .f({\u2_Display/n3190 [17],\u2_Display/n3190 [15]}),
    .fco(\u2_Display/add99/c19 ),
    .fx({\u2_Display/n3190 [18],\u2_Display/n3190 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u19_al_u5001  (
    .a({\u2_Display/n3166 ,\u2_Display/n3168 }),
    .b({\u2_Display/n3165 ,\u2_Display/n3167 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add99/c19 ),
    .f({\u2_Display/n3190 [21],\u2_Display/n3190 [19]}),
    .fco(\u2_Display/add99/c23 ),
    .fx({\u2_Display/n3190 [22],\u2_Display/n3190 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u23_al_u5002  (
    .a({\u2_Display/n3162 ,\u2_Display/n3164 }),
    .b({\u2_Display/n3161 ,\u2_Display/n3163 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add99/c23 ),
    .f({\u2_Display/n3190 [25],\u2_Display/n3190 [23]}),
    .fco(\u2_Display/add99/c27 ),
    .fx({\u2_Display/n3190 [26],\u2_Display/n3190 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u27_al_u5003  (
    .a({\u2_Display/n3158 ,\u2_Display/n3160 }),
    .b({\u2_Display/n3157 ,\u2_Display/n3159 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add99/c27 ),
    .f({\u2_Display/n3190 [29],\u2_Display/n3190 [27]}),
    .fco(\u2_Display/add99/c31 ),
    .fx({\u2_Display/n3190 [30],\u2_Display/n3190 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u31_al_u5004  (
    .a({open_n69186,\u2_Display/n3156 }),
    .c(2'b00),
    .d({open_n69191,1'b1}),
    .fci(\u2_Display/add99/c31 ),
    .f({open_n69208,\u2_Display/n3190 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u3_al_u4997  (
    .a({\u2_Display/n3182 ,\u2_Display/n3184 }),
    .b({\u2_Display/n3181 ,\u2_Display/n3183 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add99/c3 ),
    .f({\u2_Display/n3190 [5],\u2_Display/n3190 [3]}),
    .fco(\u2_Display/add99/c7 ),
    .fx({\u2_Display/n3190 [6],\u2_Display/n3190 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u7_al_u4998  (
    .a({\u2_Display/n3178 ,\u2_Display/n3180 }),
    .b({\u2_Display/n3177 ,\u2_Display/n3179 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add99/c7 ),
    .f({\u2_Display/n3190 [9],\u2_Display/n3190 [7]}),
    .fco(\u2_Display/add99/c11 ),
    .fx({\u2_Display/n3190 [10],\u2_Display/n3190 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/ucin_al_u4996  (
    .a({\u2_Display/n3186 ,1'b1}),
    .b({\u2_Display/n3185 ,\u2_Display/n3187 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3190 [1],open_n69267}),
    .fco(\u2_Display/add99/c3 ),
    .fx({\u2_Display/n3190 [2],\u2_Display/n3190 [0]}));
  EG_PHY_GCLK \u2_Display/clk1s_gclk_inst  (
    .clki(\u2_Display/clk1s ),
    .clko(\u2_Display/clk1s_gclk_net ));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A)"),
    //.LUTG0("(~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010101010101),
    .INIT_LUTG0(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/clk1s_reg  (
    .a({open_n69270,\u2_Display/clk1s }),
    .ce(\u2_Display/n35 ),
    .clk(clk_vga),
    .q({open_n69299,\u2_Display/clk1s }));  // source/rtl/Display.v(61)
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_0|u2_Display/lt0_2_cin  (
    .a({lcd_xpos[0],1'b0}),
    .b({\u2_Display/i [0],open_n69300}),
    .fco(\u2_Display/lt0_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_10|u2_Display/lt0_2_9  (
    .a(lcd_xpos[10:9]),
    .b(\u2_Display/n43 [2:1]),
    .fci(\u2_Display/lt0_2_c9 ),
    .fco(\u2_Display/lt0_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_2|u2_Display/lt0_2_1  (
    .a(lcd_xpos[2:1]),
    .b(\u2_Display/i [2:1]),
    .fci(\u2_Display/lt0_2_c1 ),
    .fco(\u2_Display/lt0_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_4|u2_Display/lt0_2_3  (
    .a(lcd_xpos[4:3]),
    .b(\u2_Display/i [4:3]),
    .fci(\u2_Display/lt0_2_c3 ),
    .fco(\u2_Display/lt0_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_6|u2_Display/lt0_2_5  (
    .a(lcd_xpos[6:5]),
    .b(\u2_Display/i [6:5]),
    .fci(\u2_Display/lt0_2_c5 ),
    .fco(\u2_Display/lt0_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_8|u2_Display/lt0_2_7  (
    .a(lcd_xpos[8:7]),
    .b({\u2_Display/n43 [0],\u2_Display/i [7]}),
    .fci(\u2_Display/lt0_2_c7 ),
    .fco(\u2_Display/lt0_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_cout|u2_Display/lt0_2_11  (
    .a({1'b0,lcd_xpos[11]}),
    .b({1'b1,\u2_Display/add2_2_co }),
    .fci(\u2_Display/lt0_2_c11 ),
    .f({\u2_Display/n44 ,open_n69464}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_0|u2_Display/lt100_cin  (
    .a({\u2_Display/n3082 ,1'b0}),
    .b({1'b0,open_n69470}),
    .fco(\u2_Display/lt100_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_10|u2_Display/lt100_9  (
    .a({\u2_Display/n3072 ,\u2_Display/n3073 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c9 ),
    .fco(\u2_Display/lt100_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_12|u2_Display/lt100_11  (
    .a({\u2_Display/n3070 ,\u2_Display/n3071 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c11 ),
    .fco(\u2_Display/lt100_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_14|u2_Display/lt100_13  (
    .a({\u2_Display/n3068 ,\u2_Display/n3069 }),
    .b(2'b11),
    .fci(\u2_Display/lt100_c13 ),
    .fco(\u2_Display/lt100_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_16|u2_Display/lt100_15  (
    .a({\u2_Display/n3066 ,\u2_Display/n3067 }),
    .b(2'b10),
    .fci(\u2_Display/lt100_c15 ),
    .fco(\u2_Display/lt100_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_18|u2_Display/lt100_17  (
    .a({\u2_Display/n3064 ,\u2_Display/n3065 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c17 ),
    .fco(\u2_Display/lt100_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_20|u2_Display/lt100_19  (
    .a({\u2_Display/n3062 ,\u2_Display/n3063 }),
    .b(2'b01),
    .fci(\u2_Display/lt100_c19 ),
    .fco(\u2_Display/lt100_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_22|u2_Display/lt100_21  (
    .a({\u2_Display/n3060 ,\u2_Display/n3061 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c21 ),
    .fco(\u2_Display/lt100_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_24|u2_Display/lt100_23  (
    .a({\u2_Display/n3058 ,\u2_Display/n3059 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c23 ),
    .fco(\u2_Display/lt100_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_26|u2_Display/lt100_25  (
    .a({\u2_Display/n3056 ,\u2_Display/n3057 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c25 ),
    .fco(\u2_Display/lt100_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_28|u2_Display/lt100_27  (
    .a({\u2_Display/n3054 ,\u2_Display/n3055 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c27 ),
    .fco(\u2_Display/lt100_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_2|u2_Display/lt100_1  (
    .a({\u2_Display/n3080 ,\u2_Display/n3081 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c1 ),
    .fco(\u2_Display/lt100_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_30|u2_Display/lt100_29  (
    .a({\u2_Display/n3052 ,\u2_Display/n3053 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c29 ),
    .fco(\u2_Display/lt100_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_4|u2_Display/lt100_3  (
    .a({\u2_Display/n3078 ,\u2_Display/n3079 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c3 ),
    .fco(\u2_Display/lt100_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_6|u2_Display/lt100_5  (
    .a({\u2_Display/n3076 ,\u2_Display/n3077 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c5 ),
    .fco(\u2_Display/lt100_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_8|u2_Display/lt100_7  (
    .a({\u2_Display/n3074 ,\u2_Display/n3075 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c7 ),
    .fco(\u2_Display/lt100_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_cout|u2_Display/lt100_31  (
    .a({1'b0,\u2_Display/n3051 }),
    .b(2'b10),
    .fci(\u2_Display/lt100_c31 ),
    .f({\u2_Display/n3083 ,open_n69874}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_0|u2_Display/lt101_cin  (
    .a({\u2_Display/n3117 ,1'b0}),
    .b({1'b0,open_n69880}),
    .fco(\u2_Display/lt101_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_10|u2_Display/lt101_9  (
    .a({\u2_Display/n3107 ,\u2_Display/n3108 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c9 ),
    .fco(\u2_Display/lt101_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_12|u2_Display/lt101_11  (
    .a({\u2_Display/n3105 ,\u2_Display/n3106 }),
    .b(2'b10),
    .fci(\u2_Display/lt101_c11 ),
    .fco(\u2_Display/lt101_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_14|u2_Display/lt101_13  (
    .a({\u2_Display/n3103 ,\u2_Display/n3104 }),
    .b(2'b01),
    .fci(\u2_Display/lt101_c13 ),
    .fco(\u2_Display/lt101_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_16|u2_Display/lt101_15  (
    .a({\u2_Display/n3101 ,\u2_Display/n3102 }),
    .b(2'b01),
    .fci(\u2_Display/lt101_c15 ),
    .fco(\u2_Display/lt101_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_18|u2_Display/lt101_17  (
    .a({\u2_Display/n3099 ,\u2_Display/n3100 }),
    .b(2'b10),
    .fci(\u2_Display/lt101_c17 ),
    .fco(\u2_Display/lt101_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_20|u2_Display/lt101_19  (
    .a({\u2_Display/n3097 ,\u2_Display/n3098 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c19 ),
    .fco(\u2_Display/lt101_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_22|u2_Display/lt101_21  (
    .a({\u2_Display/n3095 ,\u2_Display/n3096 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c21 ),
    .fco(\u2_Display/lt101_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_24|u2_Display/lt101_23  (
    .a({\u2_Display/n3093 ,\u2_Display/n3094 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c23 ),
    .fco(\u2_Display/lt101_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_26|u2_Display/lt101_25  (
    .a({\u2_Display/n3091 ,\u2_Display/n3092 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c25 ),
    .fco(\u2_Display/lt101_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_28|u2_Display/lt101_27  (
    .a({\u2_Display/n3089 ,\u2_Display/n3090 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c27 ),
    .fco(\u2_Display/lt101_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_2|u2_Display/lt101_1  (
    .a({\u2_Display/n3115 ,\u2_Display/n3116 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c1 ),
    .fco(\u2_Display/lt101_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_30|u2_Display/lt101_29  (
    .a({\u2_Display/n3087 ,\u2_Display/n3088 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c29 ),
    .fco(\u2_Display/lt101_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_4|u2_Display/lt101_3  (
    .a({\u2_Display/n3113 ,\u2_Display/n3114 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c3 ),
    .fco(\u2_Display/lt101_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_6|u2_Display/lt101_5  (
    .a({\u2_Display/n3111 ,\u2_Display/n3112 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c5 ),
    .fco(\u2_Display/lt101_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_8|u2_Display/lt101_7  (
    .a({\u2_Display/n3109 ,\u2_Display/n3110 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c7 ),
    .fco(\u2_Display/lt101_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_cout|u2_Display/lt101_31  (
    .a({1'b0,\u2_Display/n3086 }),
    .b(2'b10),
    .fci(\u2_Display/lt101_c31 ),
    .f({\u2_Display/n3118 ,open_n70284}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_0|u2_Display/lt102_cin  (
    .a({\u2_Display/n3152 ,1'b0}),
    .b({1'b0,open_n70290}),
    .fco(\u2_Display/lt102_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_10|u2_Display/lt102_9  (
    .a({\u2_Display/n3142 ,\u2_Display/n3143 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c9 ),
    .fco(\u2_Display/lt102_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_12|u2_Display/lt102_11  (
    .a({\u2_Display/n3140 ,\u2_Display/n3141 }),
    .b(2'b11),
    .fci(\u2_Display/lt102_c11 ),
    .fco(\u2_Display/lt102_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_14|u2_Display/lt102_13  (
    .a({\u2_Display/n3138 ,\u2_Display/n3139 }),
    .b(2'b10),
    .fci(\u2_Display/lt102_c13 ),
    .fco(\u2_Display/lt102_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_16|u2_Display/lt102_15  (
    .a({\u2_Display/n3136 ,\u2_Display/n3137 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c15 ),
    .fco(\u2_Display/lt102_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_18|u2_Display/lt102_17  (
    .a({\u2_Display/n3134 ,\u2_Display/n3135 }),
    .b(2'b01),
    .fci(\u2_Display/lt102_c17 ),
    .fco(\u2_Display/lt102_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_20|u2_Display/lt102_19  (
    .a({\u2_Display/n3132 ,\u2_Display/n3133 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c19 ),
    .fco(\u2_Display/lt102_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_22|u2_Display/lt102_21  (
    .a({\u2_Display/n3130 ,\u2_Display/n3131 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c21 ),
    .fco(\u2_Display/lt102_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_24|u2_Display/lt102_23  (
    .a({\u2_Display/n3128 ,\u2_Display/n3129 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c23 ),
    .fco(\u2_Display/lt102_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_26|u2_Display/lt102_25  (
    .a({\u2_Display/n3126 ,\u2_Display/n3127 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c25 ),
    .fco(\u2_Display/lt102_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_28|u2_Display/lt102_27  (
    .a({\u2_Display/n3124 ,\u2_Display/n3125 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c27 ),
    .fco(\u2_Display/lt102_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_2|u2_Display/lt102_1  (
    .a({\u2_Display/n3150 ,\u2_Display/n3151 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c1 ),
    .fco(\u2_Display/lt102_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_30|u2_Display/lt102_29  (
    .a({\u2_Display/n3122 ,\u2_Display/n3123 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c29 ),
    .fco(\u2_Display/lt102_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_4|u2_Display/lt102_3  (
    .a({\u2_Display/n3148 ,\u2_Display/n3149 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c3 ),
    .fco(\u2_Display/lt102_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_6|u2_Display/lt102_5  (
    .a({\u2_Display/n3146 ,\u2_Display/n3147 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c5 ),
    .fco(\u2_Display/lt102_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_8|u2_Display/lt102_7  (
    .a({\u2_Display/n3144 ,\u2_Display/n3145 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c7 ),
    .fco(\u2_Display/lt102_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_cout|u2_Display/lt102_31  (
    .a({1'b0,\u2_Display/n3121 }),
    .b(2'b10),
    .fci(\u2_Display/lt102_c31 ),
    .f({\u2_Display/n3153 ,open_n70694}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_0|u2_Display/lt103_cin  (
    .a({\u2_Display/n3187 ,1'b0}),
    .b({1'b0,open_n70700}),
    .fco(\u2_Display/lt103_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_10|u2_Display/lt103_9  (
    .a({\u2_Display/n3177 ,\u2_Display/n3178 }),
    .b(2'b10),
    .fci(\u2_Display/lt103_c9 ),
    .fco(\u2_Display/lt103_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_12|u2_Display/lt103_11  (
    .a({\u2_Display/n3175 ,\u2_Display/n3176 }),
    .b(2'b01),
    .fci(\u2_Display/lt103_c11 ),
    .fco(\u2_Display/lt103_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_14|u2_Display/lt103_13  (
    .a({\u2_Display/n3173 ,\u2_Display/n3174 }),
    .b(2'b01),
    .fci(\u2_Display/lt103_c13 ),
    .fco(\u2_Display/lt103_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_16|u2_Display/lt103_15  (
    .a({\u2_Display/n3171 ,\u2_Display/n3172 }),
    .b(2'b10),
    .fci(\u2_Display/lt103_c15 ),
    .fco(\u2_Display/lt103_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_18|u2_Display/lt103_17  (
    .a({\u2_Display/n3169 ,\u2_Display/n3170 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c17 ),
    .fco(\u2_Display/lt103_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_20|u2_Display/lt103_19  (
    .a({\u2_Display/n3167 ,\u2_Display/n3168 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c19 ),
    .fco(\u2_Display/lt103_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_22|u2_Display/lt103_21  (
    .a({\u2_Display/n3165 ,\u2_Display/n3166 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c21 ),
    .fco(\u2_Display/lt103_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_24|u2_Display/lt103_23  (
    .a({\u2_Display/n3163 ,\u2_Display/n3164 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c23 ),
    .fco(\u2_Display/lt103_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_26|u2_Display/lt103_25  (
    .a({\u2_Display/n3161 ,\u2_Display/n3162 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c25 ),
    .fco(\u2_Display/lt103_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_28|u2_Display/lt103_27  (
    .a({\u2_Display/n3159 ,\u2_Display/n3160 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c27 ),
    .fco(\u2_Display/lt103_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_2|u2_Display/lt103_1  (
    .a({\u2_Display/n3185 ,\u2_Display/n3186 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c1 ),
    .fco(\u2_Display/lt103_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_30|u2_Display/lt103_29  (
    .a({\u2_Display/n3157 ,\u2_Display/n3158 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c29 ),
    .fco(\u2_Display/lt103_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_4|u2_Display/lt103_3  (
    .a({\u2_Display/n3183 ,\u2_Display/n3184 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c3 ),
    .fco(\u2_Display/lt103_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_6|u2_Display/lt103_5  (
    .a({\u2_Display/n3181 ,\u2_Display/n3182 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c5 ),
    .fco(\u2_Display/lt103_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_8|u2_Display/lt103_7  (
    .a({\u2_Display/n3179 ,\u2_Display/n3180 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c7 ),
    .fco(\u2_Display/lt103_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_cout|u2_Display/lt103_31  (
    .a({1'b0,\u2_Display/n3156 }),
    .b(2'b10),
    .fci(\u2_Display/lt103_c31 ),
    .f({\u2_Display/n3188 ,open_n71104}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_0|u2_Display/lt104_cin  (
    .a({\u2_Display/n3222 ,1'b0}),
    .b({1'b0,open_n71110}),
    .fco(\u2_Display/lt104_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_10|u2_Display/lt104_9  (
    .a({\u2_Display/n3212 ,\u2_Display/n3213 }),
    .b(2'b11),
    .fci(\u2_Display/lt104_c9 ),
    .fco(\u2_Display/lt104_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_12|u2_Display/lt104_11  (
    .a({\u2_Display/n3210 ,\u2_Display/n3211 }),
    .b(2'b10),
    .fci(\u2_Display/lt104_c11 ),
    .fco(\u2_Display/lt104_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_14|u2_Display/lt104_13  (
    .a({\u2_Display/n3208 ,\u2_Display/n3209 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c13 ),
    .fco(\u2_Display/lt104_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_16|u2_Display/lt104_15  (
    .a({\u2_Display/n3206 ,\u2_Display/n3207 }),
    .b(2'b01),
    .fci(\u2_Display/lt104_c15 ),
    .fco(\u2_Display/lt104_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_18|u2_Display/lt104_17  (
    .a({\u2_Display/n3204 ,\u2_Display/n3205 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c17 ),
    .fco(\u2_Display/lt104_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_20|u2_Display/lt104_19  (
    .a({\u2_Display/n3202 ,\u2_Display/n3203 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c19 ),
    .fco(\u2_Display/lt104_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_22|u2_Display/lt104_21  (
    .a({\u2_Display/n3200 ,\u2_Display/n3201 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c21 ),
    .fco(\u2_Display/lt104_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_24|u2_Display/lt104_23  (
    .a({\u2_Display/n3198 ,\u2_Display/n3199 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c23 ),
    .fco(\u2_Display/lt104_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_26|u2_Display/lt104_25  (
    .a({\u2_Display/n3196 ,\u2_Display/n3197 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c25 ),
    .fco(\u2_Display/lt104_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_28|u2_Display/lt104_27  (
    .a({\u2_Display/n3194 ,\u2_Display/n3195 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c27 ),
    .fco(\u2_Display/lt104_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_2|u2_Display/lt104_1  (
    .a({\u2_Display/n3220 ,\u2_Display/n3221 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c1 ),
    .fco(\u2_Display/lt104_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_30|u2_Display/lt104_29  (
    .a({\u2_Display/n3192 ,\u2_Display/n3193 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c29 ),
    .fco(\u2_Display/lt104_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_4|u2_Display/lt104_3  (
    .a({\u2_Display/n3218 ,\u2_Display/n3219 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c3 ),
    .fco(\u2_Display/lt104_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_6|u2_Display/lt104_5  (
    .a({\u2_Display/n3216 ,\u2_Display/n3217 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c5 ),
    .fco(\u2_Display/lt104_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_8|u2_Display/lt104_7  (
    .a({\u2_Display/n3214 ,\u2_Display/n3215 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c7 ),
    .fco(\u2_Display/lt104_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_cout|u2_Display/lt104_31  (
    .a({1'b0,\u2_Display/n3191 }),
    .b(2'b10),
    .fci(\u2_Display/lt104_c31 ),
    .f({\u2_Display/n3223 ,open_n71514}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_0|u2_Display/lt105_cin  (
    .a({\u2_Display/n3257 ,1'b0}),
    .b({1'b0,open_n71520}),
    .fco(\u2_Display/lt105_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_10|u2_Display/lt105_9  (
    .a({\u2_Display/n3247 ,\u2_Display/n3248 }),
    .b(2'b01),
    .fci(\u2_Display/lt105_c9 ),
    .fco(\u2_Display/lt105_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_12|u2_Display/lt105_11  (
    .a({\u2_Display/n3245 ,\u2_Display/n3246 }),
    .b(2'b01),
    .fci(\u2_Display/lt105_c11 ),
    .fco(\u2_Display/lt105_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_14|u2_Display/lt105_13  (
    .a({\u2_Display/n3243 ,\u2_Display/n3244 }),
    .b(2'b10),
    .fci(\u2_Display/lt105_c13 ),
    .fco(\u2_Display/lt105_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_16|u2_Display/lt105_15  (
    .a({\u2_Display/n3241 ,\u2_Display/n3242 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c15 ),
    .fco(\u2_Display/lt105_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_18|u2_Display/lt105_17  (
    .a({\u2_Display/n3239 ,\u2_Display/n3240 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c17 ),
    .fco(\u2_Display/lt105_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_20|u2_Display/lt105_19  (
    .a({\u2_Display/n3237 ,\u2_Display/n3238 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c19 ),
    .fco(\u2_Display/lt105_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_22|u2_Display/lt105_21  (
    .a({\u2_Display/n3235 ,\u2_Display/n3236 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c21 ),
    .fco(\u2_Display/lt105_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_24|u2_Display/lt105_23  (
    .a({\u2_Display/n3233 ,\u2_Display/n3234 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c23 ),
    .fco(\u2_Display/lt105_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_26|u2_Display/lt105_25  (
    .a({\u2_Display/n3231 ,\u2_Display/n3232 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c25 ),
    .fco(\u2_Display/lt105_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_28|u2_Display/lt105_27  (
    .a({\u2_Display/n3229 ,\u2_Display/n3230 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c27 ),
    .fco(\u2_Display/lt105_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_2|u2_Display/lt105_1  (
    .a({\u2_Display/n3255 ,\u2_Display/n3256 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c1 ),
    .fco(\u2_Display/lt105_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_30|u2_Display/lt105_29  (
    .a({\u2_Display/n3227 ,\u2_Display/n3228 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c29 ),
    .fco(\u2_Display/lt105_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_4|u2_Display/lt105_3  (
    .a({\u2_Display/n3253 ,\u2_Display/n3254 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c3 ),
    .fco(\u2_Display/lt105_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_6|u2_Display/lt105_5  (
    .a({\u2_Display/n3251 ,\u2_Display/n3252 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c5 ),
    .fco(\u2_Display/lt105_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_8|u2_Display/lt105_7  (
    .a({\u2_Display/n3249 ,\u2_Display/n3250 }),
    .b(2'b10),
    .fci(\u2_Display/lt105_c7 ),
    .fco(\u2_Display/lt105_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_cout|u2_Display/lt105_31  (
    .a({1'b0,\u2_Display/n3226 }),
    .b(2'b10),
    .fci(\u2_Display/lt105_c31 ),
    .f({\u2_Display/n3258 ,open_n71924}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_0|u2_Display/lt106_cin  (
    .a({\u2_Display/n3292 ,1'b0}),
    .b({1'b0,open_n71930}),
    .fco(\u2_Display/lt106_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_10|u2_Display/lt106_9  (
    .a({\u2_Display/n3282 ,\u2_Display/n3283 }),
    .b(2'b10),
    .fci(\u2_Display/lt106_c9 ),
    .fco(\u2_Display/lt106_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_12|u2_Display/lt106_11  (
    .a({\u2_Display/n3280 ,\u2_Display/n3281 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c11 ),
    .fco(\u2_Display/lt106_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_14|u2_Display/lt106_13  (
    .a({\u2_Display/n3278 ,\u2_Display/n3279 }),
    .b(2'b01),
    .fci(\u2_Display/lt106_c13 ),
    .fco(\u2_Display/lt106_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_16|u2_Display/lt106_15  (
    .a({\u2_Display/n3276 ,\u2_Display/n3277 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c15 ),
    .fco(\u2_Display/lt106_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_18|u2_Display/lt106_17  (
    .a({\u2_Display/n3274 ,\u2_Display/n3275 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c17 ),
    .fco(\u2_Display/lt106_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_20|u2_Display/lt106_19  (
    .a({\u2_Display/n3272 ,\u2_Display/n3273 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c19 ),
    .fco(\u2_Display/lt106_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_22|u2_Display/lt106_21  (
    .a({\u2_Display/n3270 ,\u2_Display/n3271 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c21 ),
    .fco(\u2_Display/lt106_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_24|u2_Display/lt106_23  (
    .a({\u2_Display/n3268 ,\u2_Display/n3269 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c23 ),
    .fco(\u2_Display/lt106_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_26|u2_Display/lt106_25  (
    .a({\u2_Display/n3266 ,\u2_Display/n3267 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c25 ),
    .fco(\u2_Display/lt106_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_28|u2_Display/lt106_27  (
    .a({\u2_Display/n3264 ,\u2_Display/n3265 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c27 ),
    .fco(\u2_Display/lt106_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_2|u2_Display/lt106_1  (
    .a({\u2_Display/n3290 ,\u2_Display/n3291 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c1 ),
    .fco(\u2_Display/lt106_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_30|u2_Display/lt106_29  (
    .a({\u2_Display/n3262 ,\u2_Display/n3263 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c29 ),
    .fco(\u2_Display/lt106_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_4|u2_Display/lt106_3  (
    .a({\u2_Display/n3288 ,\u2_Display/n3289 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c3 ),
    .fco(\u2_Display/lt106_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_6|u2_Display/lt106_5  (
    .a({\u2_Display/n3286 ,\u2_Display/n3287 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c5 ),
    .fco(\u2_Display/lt106_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_8|u2_Display/lt106_7  (
    .a({\u2_Display/n3284 ,\u2_Display/n3285 }),
    .b(2'b11),
    .fci(\u2_Display/lt106_c7 ),
    .fco(\u2_Display/lt106_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_cout|u2_Display/lt106_31  (
    .a({1'b0,\u2_Display/n3261 }),
    .b(2'b10),
    .fci(\u2_Display/lt106_c31 ),
    .f({\u2_Display/n3293 ,open_n72334}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_0|u2_Display/lt107_cin  (
    .a({\u2_Display/n3327 ,1'b0}),
    .b({1'b0,open_n72340}),
    .fco(\u2_Display/lt107_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_10|u2_Display/lt107_9  (
    .a({\u2_Display/n3317 ,\u2_Display/n3318 }),
    .b(2'b01),
    .fci(\u2_Display/lt107_c9 ),
    .fco(\u2_Display/lt107_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_12|u2_Display/lt107_11  (
    .a({\u2_Display/n3315 ,\u2_Display/n3316 }),
    .b(2'b10),
    .fci(\u2_Display/lt107_c11 ),
    .fco(\u2_Display/lt107_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_14|u2_Display/lt107_13  (
    .a({\u2_Display/n3313 ,\u2_Display/n3314 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c13 ),
    .fco(\u2_Display/lt107_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_16|u2_Display/lt107_15  (
    .a({\u2_Display/n3311 ,\u2_Display/n3312 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c15 ),
    .fco(\u2_Display/lt107_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_18|u2_Display/lt107_17  (
    .a({\u2_Display/n3309 ,\u2_Display/n3310 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c17 ),
    .fco(\u2_Display/lt107_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_20|u2_Display/lt107_19  (
    .a({\u2_Display/n3307 ,\u2_Display/n3308 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c19 ),
    .fco(\u2_Display/lt107_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_22|u2_Display/lt107_21  (
    .a({\u2_Display/n3305 ,\u2_Display/n3306 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c21 ),
    .fco(\u2_Display/lt107_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_24|u2_Display/lt107_23  (
    .a({\u2_Display/n3303 ,\u2_Display/n3304 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c23 ),
    .fco(\u2_Display/lt107_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_26|u2_Display/lt107_25  (
    .a({\u2_Display/n3301 ,\u2_Display/n3302 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c25 ),
    .fco(\u2_Display/lt107_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_28|u2_Display/lt107_27  (
    .a({\u2_Display/n3299 ,\u2_Display/n3300 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c27 ),
    .fco(\u2_Display/lt107_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_2|u2_Display/lt107_1  (
    .a({\u2_Display/n3325 ,\u2_Display/n3326 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c1 ),
    .fco(\u2_Display/lt107_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_30|u2_Display/lt107_29  (
    .a({\u2_Display/n3297 ,\u2_Display/n3298 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c29 ),
    .fco(\u2_Display/lt107_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_4|u2_Display/lt107_3  (
    .a({\u2_Display/n3323 ,\u2_Display/n3324 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c3 ),
    .fco(\u2_Display/lt107_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_6|u2_Display/lt107_5  (
    .a({\u2_Display/n3321 ,\u2_Display/n3322 }),
    .b(2'b10),
    .fci(\u2_Display/lt107_c5 ),
    .fco(\u2_Display/lt107_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_8|u2_Display/lt107_7  (
    .a({\u2_Display/n3319 ,\u2_Display/n3320 }),
    .b(2'b01),
    .fci(\u2_Display/lt107_c7 ),
    .fco(\u2_Display/lt107_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_cout|u2_Display/lt107_31  (
    .a({1'b0,\u2_Display/n3296 }),
    .b(2'b10),
    .fci(\u2_Display/lt107_c31 ),
    .f({\u2_Display/n3328 ,open_n72744}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_0|u2_Display/lt108_cin  (
    .a({\u2_Display/n3362 ,1'b0}),
    .b({1'b0,open_n72750}),
    .fco(\u2_Display/lt108_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_10|u2_Display/lt108_9  (
    .a({\u2_Display/n3352 ,\u2_Display/n3353 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c9 ),
    .fco(\u2_Display/lt108_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_12|u2_Display/lt108_11  (
    .a({\u2_Display/n3350 ,\u2_Display/n3351 }),
    .b(2'b01),
    .fci(\u2_Display/lt108_c11 ),
    .fco(\u2_Display/lt108_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_14|u2_Display/lt108_13  (
    .a({\u2_Display/n3348 ,\u2_Display/n3349 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c13 ),
    .fco(\u2_Display/lt108_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_16|u2_Display/lt108_15  (
    .a({\u2_Display/n3346 ,\u2_Display/n3347 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c15 ),
    .fco(\u2_Display/lt108_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_18|u2_Display/lt108_17  (
    .a({\u2_Display/n3344 ,\u2_Display/n3345 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c17 ),
    .fco(\u2_Display/lt108_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_20|u2_Display/lt108_19  (
    .a({\u2_Display/n3342 ,\u2_Display/n3343 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c19 ),
    .fco(\u2_Display/lt108_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_22|u2_Display/lt108_21  (
    .a({\u2_Display/n3340 ,\u2_Display/n3341 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c21 ),
    .fco(\u2_Display/lt108_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_24|u2_Display/lt108_23  (
    .a({\u2_Display/n3338 ,\u2_Display/n3339 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c23 ),
    .fco(\u2_Display/lt108_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_26|u2_Display/lt108_25  (
    .a({\u2_Display/n3336 ,\u2_Display/n3337 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c25 ),
    .fco(\u2_Display/lt108_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_28|u2_Display/lt108_27  (
    .a({\u2_Display/n3334 ,\u2_Display/n3335 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c27 ),
    .fco(\u2_Display/lt108_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_2|u2_Display/lt108_1  (
    .a({\u2_Display/n3360 ,\u2_Display/n3361 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c1 ),
    .fco(\u2_Display/lt108_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_30|u2_Display/lt108_29  (
    .a({\u2_Display/n3332 ,\u2_Display/n3333 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c29 ),
    .fco(\u2_Display/lt108_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_4|u2_Display/lt108_3  (
    .a({\u2_Display/n3358 ,\u2_Display/n3359 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c3 ),
    .fco(\u2_Display/lt108_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_6|u2_Display/lt108_5  (
    .a({\u2_Display/n3356 ,\u2_Display/n3357 }),
    .b(2'b11),
    .fci(\u2_Display/lt108_c5 ),
    .fco(\u2_Display/lt108_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_8|u2_Display/lt108_7  (
    .a({\u2_Display/n3354 ,\u2_Display/n3355 }),
    .b(2'b10),
    .fci(\u2_Display/lt108_c7 ),
    .fco(\u2_Display/lt108_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_cout|u2_Display/lt108_31  (
    .a({1'b0,\u2_Display/n3331 }),
    .b(2'b10),
    .fci(\u2_Display/lt108_c31 ),
    .f({\u2_Display/n3363 ,open_n73154}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_0|u2_Display/lt109_cin  (
    .a({\u2_Display/n3397 ,1'b0}),
    .b({1'b0,open_n73160}),
    .fco(\u2_Display/lt109_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_10|u2_Display/lt109_9  (
    .a({\u2_Display/n3387 ,\u2_Display/n3388 }),
    .b(2'b10),
    .fci(\u2_Display/lt109_c9 ),
    .fco(\u2_Display/lt109_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_12|u2_Display/lt109_11  (
    .a({\u2_Display/n3385 ,\u2_Display/n3386 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c11 ),
    .fco(\u2_Display/lt109_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_14|u2_Display/lt109_13  (
    .a({\u2_Display/n3383 ,\u2_Display/n3384 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c13 ),
    .fco(\u2_Display/lt109_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_16|u2_Display/lt109_15  (
    .a({\u2_Display/n3381 ,\u2_Display/n3382 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c15 ),
    .fco(\u2_Display/lt109_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_18|u2_Display/lt109_17  (
    .a({\u2_Display/n3379 ,\u2_Display/n3380 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c17 ),
    .fco(\u2_Display/lt109_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_20|u2_Display/lt109_19  (
    .a({\u2_Display/n3377 ,\u2_Display/n3378 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c19 ),
    .fco(\u2_Display/lt109_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_22|u2_Display/lt109_21  (
    .a({\u2_Display/n3375 ,\u2_Display/n3376 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c21 ),
    .fco(\u2_Display/lt109_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_24|u2_Display/lt109_23  (
    .a({\u2_Display/n3373 ,\u2_Display/n3374 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c23 ),
    .fco(\u2_Display/lt109_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_26|u2_Display/lt109_25  (
    .a({\u2_Display/n3371 ,\u2_Display/n3372 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c25 ),
    .fco(\u2_Display/lt109_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_28|u2_Display/lt109_27  (
    .a({\u2_Display/n3369 ,\u2_Display/n3370 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c27 ),
    .fco(\u2_Display/lt109_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_2|u2_Display/lt109_1  (
    .a({\u2_Display/n3395 ,\u2_Display/n3396 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c1 ),
    .fco(\u2_Display/lt109_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_30|u2_Display/lt109_29  (
    .a({\u2_Display/n3367 ,\u2_Display/n3368 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c29 ),
    .fco(\u2_Display/lt109_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_4|u2_Display/lt109_3  (
    .a({\u2_Display/n3393 ,\u2_Display/n3394 }),
    .b(2'b10),
    .fci(\u2_Display/lt109_c3 ),
    .fco(\u2_Display/lt109_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_6|u2_Display/lt109_5  (
    .a({\u2_Display/n3391 ,\u2_Display/n3392 }),
    .b(2'b01),
    .fci(\u2_Display/lt109_c5 ),
    .fco(\u2_Display/lt109_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_8|u2_Display/lt109_7  (
    .a({\u2_Display/n3389 ,\u2_Display/n3390 }),
    .b(2'b01),
    .fci(\u2_Display/lt109_c7 ),
    .fco(\u2_Display/lt109_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_cout|u2_Display/lt109_31  (
    .a({1'b0,\u2_Display/n3366 }),
    .b(2'b10),
    .fci(\u2_Display/lt109_c31 ),
    .f({\u2_Display/n3398 ,open_n73564}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_0|u2_Display/lt10_2_cin  (
    .a({lcd_ypos[0],1'b0}),
    .b({\u2_Display/i [0],open_n73570}),
    .fco(\u2_Display/lt10_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_10|u2_Display/lt10_2_9  (
    .a(lcd_ypos[10:9]),
    .b(\u2_Display/n140 [1:0]),
    .fci(\u2_Display/lt10_2_c9 ),
    .fco(\u2_Display/lt10_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_2|u2_Display/lt10_2_1  (
    .a(lcd_ypos[2:1]),
    .b(\u2_Display/i [2:1]),
    .fci(\u2_Display/lt10_2_c1 ),
    .fco(\u2_Display/lt10_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_4|u2_Display/lt10_2_3  (
    .a(lcd_ypos[4:3]),
    .b(\u2_Display/i [4:3]),
    .fci(\u2_Display/lt10_2_c3 ),
    .fco(\u2_Display/lt10_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_6|u2_Display/lt10_2_5  (
    .a(lcd_ypos[6:5]),
    .b(\u2_Display/i [6:5]),
    .fci(\u2_Display/lt10_2_c5 ),
    .fco(\u2_Display/lt10_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_8|u2_Display/lt10_2_7  (
    .a(lcd_ypos[8:7]),
    .b(\u2_Display/i [8:7]),
    .fci(\u2_Display/lt10_2_c7 ),
    .fco(\u2_Display/lt10_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_cout|u2_Display/lt10_2_11  (
    .a({1'b0,lcd_ypos[11]}),
    .b({1'b1,\u2_Display/add7_2_co }),
    .fci(\u2_Display/lt10_2_c11 ),
    .f({\u2_Display/n141 ,open_n73734}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_0|u2_Display/lt110_cin  (
    .a({\u2_Display/n3432 ,1'b0}),
    .b({1'b0,open_n73740}),
    .fco(\u2_Display/lt110_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_10|u2_Display/lt110_9  (
    .a({\u2_Display/n3422 ,\u2_Display/n3423 }),
    .b(2'b01),
    .fci(\u2_Display/lt110_c9 ),
    .fco(\u2_Display/lt110_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_12|u2_Display/lt110_11  (
    .a({\u2_Display/n3420 ,\u2_Display/n3421 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c11 ),
    .fco(\u2_Display/lt110_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_14|u2_Display/lt110_13  (
    .a({\u2_Display/n3418 ,\u2_Display/n3419 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c13 ),
    .fco(\u2_Display/lt110_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_16|u2_Display/lt110_15  (
    .a({\u2_Display/n3416 ,\u2_Display/n3417 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c15 ),
    .fco(\u2_Display/lt110_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_18|u2_Display/lt110_17  (
    .a({\u2_Display/n3414 ,\u2_Display/n3415 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c17 ),
    .fco(\u2_Display/lt110_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_20|u2_Display/lt110_19  (
    .a({\u2_Display/n3412 ,\u2_Display/n3413 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c19 ),
    .fco(\u2_Display/lt110_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_22|u2_Display/lt110_21  (
    .a({\u2_Display/n3410 ,\u2_Display/n3411 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c21 ),
    .fco(\u2_Display/lt110_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_24|u2_Display/lt110_23  (
    .a({\u2_Display/n3408 ,\u2_Display/n3409 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c23 ),
    .fco(\u2_Display/lt110_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_26|u2_Display/lt110_25  (
    .a({\u2_Display/n3406 ,\u2_Display/n3407 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c25 ),
    .fco(\u2_Display/lt110_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_28|u2_Display/lt110_27  (
    .a({\u2_Display/n3404 ,\u2_Display/n3405 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c27 ),
    .fco(\u2_Display/lt110_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_2|u2_Display/lt110_1  (
    .a({\u2_Display/n3430 ,\u2_Display/n3431 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c1 ),
    .fco(\u2_Display/lt110_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_30|u2_Display/lt110_29  (
    .a({\u2_Display/n3402 ,\u2_Display/n3403 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c29 ),
    .fco(\u2_Display/lt110_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_4|u2_Display/lt110_3  (
    .a({\u2_Display/n3428 ,\u2_Display/n3429 }),
    .b(2'b11),
    .fci(\u2_Display/lt110_c3 ),
    .fco(\u2_Display/lt110_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_6|u2_Display/lt110_5  (
    .a({\u2_Display/n3426 ,\u2_Display/n3427 }),
    .b(2'b10),
    .fci(\u2_Display/lt110_c5 ),
    .fco(\u2_Display/lt110_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_8|u2_Display/lt110_7  (
    .a({\u2_Display/n3424 ,\u2_Display/n3425 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c7 ),
    .fco(\u2_Display/lt110_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_cout|u2_Display/lt110_31  (
    .a({1'b0,\u2_Display/n3401 }),
    .b(2'b10),
    .fci(\u2_Display/lt110_c31 ),
    .f({\u2_Display/n3433 ,open_n74144}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_0|u2_Display/lt11_2_cin  (
    .a({\u2_Display/n143 [0],1'b0}),
    .b({lcd_ypos[0],open_n74150}),
    .fco(\u2_Display/lt11_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_10|u2_Display/lt11_2_9  (
    .a(\u2_Display/n143 [10:9]),
    .b(lcd_ypos[10:9]),
    .fci(\u2_Display/lt11_2_c9 ),
    .fco(\u2_Display/lt11_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_12|u2_Display/lt11_2_11  (
    .a({\u2_Display/n143 [31],\u2_Display/n143 [31]}),
    .b({1'b0,lcd_ypos[11]}),
    .fci(\u2_Display/lt11_2_c11 ),
    .fco(\u2_Display/lt11_2_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_2|u2_Display/lt11_2_1  (
    .a(\u2_Display/n143 [2:1]),
    .b(lcd_ypos[2:1]),
    .fci(\u2_Display/lt11_2_c1 ),
    .fco(\u2_Display/lt11_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_4|u2_Display/lt11_2_3  (
    .a(\u2_Display/n143 [4:3]),
    .b(lcd_ypos[4:3]),
    .fci(\u2_Display/lt11_2_c3 ),
    .fco(\u2_Display/lt11_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_6|u2_Display/lt11_2_5  (
    .a(\u2_Display/n143 [6:5]),
    .b(lcd_ypos[6:5]),
    .fci(\u2_Display/lt11_2_c5 ),
    .fco(\u2_Display/lt11_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_8|u2_Display/lt11_2_7  (
    .a(\u2_Display/n143 [8:7]),
    .b(lcd_ypos[8:7]),
    .fci(\u2_Display/lt11_2_c7 ),
    .fco(\u2_Display/lt11_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_cout_al_u5060  (
    .a({open_n74320,1'b0}),
    .b({open_n74321,1'b1}),
    .fci(\u2_Display/lt11_2_c13 ),
    .f({open_n74340,\u2_Display/n144 }));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_0|u2_Display/lt121_cin  (
    .a({\u2_Display/counta [0],1'b0}),
    .b({1'b0,open_n74346}),
    .fco(\u2_Display/lt121_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_10|u2_Display/lt121_9  (
    .a(\u2_Display/counta [10:9]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c9 ),
    .fco(\u2_Display/lt121_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_12|u2_Display/lt121_11  (
    .a(\u2_Display/counta [12:11]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c11 ),
    .fco(\u2_Display/lt121_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_14|u2_Display/lt121_13  (
    .a(\u2_Display/counta [14:13]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c13 ),
    .fco(\u2_Display/lt121_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_16|u2_Display/lt121_15  (
    .a(\u2_Display/counta [16:15]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c15 ),
    .fco(\u2_Display/lt121_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_18|u2_Display/lt121_17  (
    .a(\u2_Display/counta [18:17]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c17 ),
    .fco(\u2_Display/lt121_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_20|u2_Display/lt121_19  (
    .a(\u2_Display/counta [20:19]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c19 ),
    .fco(\u2_Display/lt121_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_22|u2_Display/lt121_21  (
    .a(\u2_Display/counta [22:21]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c21 ),
    .fco(\u2_Display/lt121_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_24|u2_Display/lt121_23  (
    .a(\u2_Display/counta [24:23]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c23 ),
    .fco(\u2_Display/lt121_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_26|u2_Display/lt121_25  (
    .a(\u2_Display/counta [26:25]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c25 ),
    .fco(\u2_Display/lt121_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_28|u2_Display/lt121_27  (
    .a(\u2_Display/counta [28:27]),
    .b(2'b01),
    .fci(\u2_Display/lt121_c27 ),
    .fco(\u2_Display/lt121_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_2|u2_Display/lt121_1  (
    .a(\u2_Display/counta [2:1]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c1 ),
    .fco(\u2_Display/lt121_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_30|u2_Display/lt121_29  (
    .a(\u2_Display/counta [30:29]),
    .b(2'b10),
    .fci(\u2_Display/lt121_c29 ),
    .fco(\u2_Display/lt121_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_4|u2_Display/lt121_3  (
    .a(\u2_Display/counta [4:3]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c3 ),
    .fco(\u2_Display/lt121_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_6|u2_Display/lt121_5  (
    .a(\u2_Display/counta [6:5]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c5 ),
    .fco(\u2_Display/lt121_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_8|u2_Display/lt121_7  (
    .a(\u2_Display/counta [8:7]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c7 ),
    .fco(\u2_Display/lt121_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_cout|u2_Display/lt121_31  (
    .a({1'b0,\u2_Display/counta [31]}),
    .b(2'b11),
    .fci(\u2_Display/lt121_c31 ),
    .f({\u2_Display/n3786 ,open_n74750}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_0|u2_Display/lt122_cin  (
    .a({\u2_Display/n3820 ,1'b0}),
    .b({1'b0,open_n74756}),
    .fco(\u2_Display/lt122_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_10|u2_Display/lt122_9  (
    .a({\u2_Display/n3810 ,\u2_Display/n3811 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c9 ),
    .fco(\u2_Display/lt122_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_12|u2_Display/lt122_11  (
    .a({\u2_Display/n3808 ,\u2_Display/n3809 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c11 ),
    .fco(\u2_Display/lt122_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_14|u2_Display/lt122_13  (
    .a({\u2_Display/n3806 ,\u2_Display/n3807 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c13 ),
    .fco(\u2_Display/lt122_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_16|u2_Display/lt122_15  (
    .a({\u2_Display/n3804 ,\u2_Display/n3805 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c15 ),
    .fco(\u2_Display/lt122_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_18|u2_Display/lt122_17  (
    .a({\u2_Display/n3802 ,\u2_Display/n3803 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c17 ),
    .fco(\u2_Display/lt122_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_20|u2_Display/lt122_19  (
    .a({\u2_Display/n3800 ,\u2_Display/n3801 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c19 ),
    .fco(\u2_Display/lt122_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_22|u2_Display/lt122_21  (
    .a({\u2_Display/n3798 ,\u2_Display/n3799 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c21 ),
    .fco(\u2_Display/lt122_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_24|u2_Display/lt122_23  (
    .a({\u2_Display/n3796 ,\u2_Display/n3797 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c23 ),
    .fco(\u2_Display/lt122_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_26|u2_Display/lt122_25  (
    .a({\u2_Display/n3794 ,\u2_Display/n3795 }),
    .b(2'b10),
    .fci(\u2_Display/lt122_c25 ),
    .fco(\u2_Display/lt122_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_28|u2_Display/lt122_27  (
    .a({\u2_Display/n3792 ,\u2_Display/n3793 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c27 ),
    .fco(\u2_Display/lt122_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_2|u2_Display/lt122_1  (
    .a({\u2_Display/n3818 ,\u2_Display/n3819 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c1 ),
    .fco(\u2_Display/lt122_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_30|u2_Display/lt122_29  (
    .a({\u2_Display/n3790 ,\u2_Display/n3791 }),
    .b(2'b11),
    .fci(\u2_Display/lt122_c29 ),
    .fco(\u2_Display/lt122_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_4|u2_Display/lt122_3  (
    .a({\u2_Display/n3816 ,\u2_Display/n3817 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c3 ),
    .fco(\u2_Display/lt122_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_6|u2_Display/lt122_5  (
    .a({\u2_Display/n3814 ,\u2_Display/n3815 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c5 ),
    .fco(\u2_Display/lt122_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_8|u2_Display/lt122_7  (
    .a({\u2_Display/n3812 ,\u2_Display/n3813 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c7 ),
    .fco(\u2_Display/lt122_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_cout|u2_Display/lt122_31  (
    .a({1'b0,\u2_Display/n3789 }),
    .b(2'b10),
    .fci(\u2_Display/lt122_c31 ),
    .f({\u2_Display/n3821 ,open_n75160}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_0|u2_Display/lt123_cin  (
    .a({\u2_Display/n3855 ,1'b0}),
    .b({1'b0,open_n75166}),
    .fco(\u2_Display/lt123_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_10|u2_Display/lt123_9  (
    .a({\u2_Display/n3845 ,\u2_Display/n3846 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c9 ),
    .fco(\u2_Display/lt123_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_12|u2_Display/lt123_11  (
    .a({\u2_Display/n3843 ,\u2_Display/n3844 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c11 ),
    .fco(\u2_Display/lt123_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_14|u2_Display/lt123_13  (
    .a({\u2_Display/n3841 ,\u2_Display/n3842 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c13 ),
    .fco(\u2_Display/lt123_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_16|u2_Display/lt123_15  (
    .a({\u2_Display/n3839 ,\u2_Display/n3840 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c15 ),
    .fco(\u2_Display/lt123_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_18|u2_Display/lt123_17  (
    .a({\u2_Display/n3837 ,\u2_Display/n3838 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c17 ),
    .fco(\u2_Display/lt123_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_20|u2_Display/lt123_19  (
    .a({\u2_Display/n3835 ,\u2_Display/n3836 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c19 ),
    .fco(\u2_Display/lt123_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_22|u2_Display/lt123_21  (
    .a({\u2_Display/n3833 ,\u2_Display/n3834 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c21 ),
    .fco(\u2_Display/lt123_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_24|u2_Display/lt123_23  (
    .a({\u2_Display/n3831 ,\u2_Display/n3832 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c23 ),
    .fco(\u2_Display/lt123_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_26|u2_Display/lt123_25  (
    .a({\u2_Display/n3829 ,\u2_Display/n3830 }),
    .b(2'b01),
    .fci(\u2_Display/lt123_c25 ),
    .fco(\u2_Display/lt123_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_28|u2_Display/lt123_27  (
    .a({\u2_Display/n3827 ,\u2_Display/n3828 }),
    .b(2'b10),
    .fci(\u2_Display/lt123_c27 ),
    .fco(\u2_Display/lt123_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_2|u2_Display/lt123_1  (
    .a({\u2_Display/n3853 ,\u2_Display/n3854 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c1 ),
    .fco(\u2_Display/lt123_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_30|u2_Display/lt123_29  (
    .a({\u2_Display/n3825 ,\u2_Display/n3826 }),
    .b(2'b01),
    .fci(\u2_Display/lt123_c29 ),
    .fco(\u2_Display/lt123_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_4|u2_Display/lt123_3  (
    .a({\u2_Display/n3851 ,\u2_Display/n3852 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c3 ),
    .fco(\u2_Display/lt123_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_6|u2_Display/lt123_5  (
    .a({\u2_Display/n3849 ,\u2_Display/n3850 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c5 ),
    .fco(\u2_Display/lt123_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_8|u2_Display/lt123_7  (
    .a({\u2_Display/n3847 ,\u2_Display/n3848 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c7 ),
    .fco(\u2_Display/lt123_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_cout|u2_Display/lt123_31  (
    .a({1'b0,\u2_Display/n3824 }),
    .b(2'b10),
    .fci(\u2_Display/lt123_c31 ),
    .f({\u2_Display/n3856 ,open_n75570}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_0|u2_Display/lt124_cin  (
    .a({\u2_Display/n3890 ,1'b0}),
    .b({1'b0,open_n75576}),
    .fco(\u2_Display/lt124_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_10|u2_Display/lt124_9  (
    .a({\u2_Display/n3880 ,\u2_Display/n3881 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c9 ),
    .fco(\u2_Display/lt124_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_12|u2_Display/lt124_11  (
    .a({\u2_Display/n3878 ,\u2_Display/n3879 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c11 ),
    .fco(\u2_Display/lt124_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_14|u2_Display/lt124_13  (
    .a({\u2_Display/n3876 ,\u2_Display/n3877 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c13 ),
    .fco(\u2_Display/lt124_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_16|u2_Display/lt124_15  (
    .a({\u2_Display/n3874 ,\u2_Display/n3875 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c15 ),
    .fco(\u2_Display/lt124_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_18|u2_Display/lt124_17  (
    .a({\u2_Display/n3872 ,\u2_Display/n3873 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c17 ),
    .fco(\u2_Display/lt124_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_20|u2_Display/lt124_19  (
    .a({\u2_Display/n3870 ,\u2_Display/n3871 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c19 ),
    .fco(\u2_Display/lt124_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_22|u2_Display/lt124_21  (
    .a({\u2_Display/n3868 ,\u2_Display/n3869 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c21 ),
    .fco(\u2_Display/lt124_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_24|u2_Display/lt124_23  (
    .a({\u2_Display/n3866 ,\u2_Display/n3867 }),
    .b(2'b10),
    .fci(\u2_Display/lt124_c23 ),
    .fco(\u2_Display/lt124_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_26|u2_Display/lt124_25  (
    .a({\u2_Display/n3864 ,\u2_Display/n3865 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c25 ),
    .fco(\u2_Display/lt124_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_28|u2_Display/lt124_27  (
    .a({\u2_Display/n3862 ,\u2_Display/n3863 }),
    .b(2'b11),
    .fci(\u2_Display/lt124_c27 ),
    .fco(\u2_Display/lt124_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_2|u2_Display/lt124_1  (
    .a({\u2_Display/n3888 ,\u2_Display/n3889 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c1 ),
    .fco(\u2_Display/lt124_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_30|u2_Display/lt124_29  (
    .a({\u2_Display/n3860 ,\u2_Display/n3861 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c29 ),
    .fco(\u2_Display/lt124_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_4|u2_Display/lt124_3  (
    .a({\u2_Display/n3886 ,\u2_Display/n3887 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c3 ),
    .fco(\u2_Display/lt124_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_6|u2_Display/lt124_5  (
    .a({\u2_Display/n3884 ,\u2_Display/n3885 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c5 ),
    .fco(\u2_Display/lt124_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_8|u2_Display/lt124_7  (
    .a({\u2_Display/n3882 ,\u2_Display/n3883 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c7 ),
    .fco(\u2_Display/lt124_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_cout|u2_Display/lt124_31  (
    .a({1'b0,\u2_Display/n3859 }),
    .b(2'b10),
    .fci(\u2_Display/lt124_c31 ),
    .f({\u2_Display/n3891 ,open_n75980}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_0|u2_Display/lt125_cin  (
    .a({\u2_Display/n3925 ,1'b0}),
    .b({1'b0,open_n75986}),
    .fco(\u2_Display/lt125_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_10|u2_Display/lt125_9  (
    .a({\u2_Display/n3915 ,\u2_Display/n3916 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c9 ),
    .fco(\u2_Display/lt125_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_12|u2_Display/lt125_11  (
    .a({\u2_Display/n3913 ,\u2_Display/n3914 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c11 ),
    .fco(\u2_Display/lt125_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_14|u2_Display/lt125_13  (
    .a({\u2_Display/n3911 ,\u2_Display/n3912 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c13 ),
    .fco(\u2_Display/lt125_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_16|u2_Display/lt125_15  (
    .a({\u2_Display/n3909 ,\u2_Display/n3910 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c15 ),
    .fco(\u2_Display/lt125_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_18|u2_Display/lt125_17  (
    .a({\u2_Display/n3907 ,\u2_Display/n3908 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c17 ),
    .fco(\u2_Display/lt125_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_20|u2_Display/lt125_19  (
    .a({\u2_Display/n3905 ,\u2_Display/n3906 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c19 ),
    .fco(\u2_Display/lt125_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_22|u2_Display/lt125_21  (
    .a({\u2_Display/n3903 ,\u2_Display/n3904 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c21 ),
    .fco(\u2_Display/lt125_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_24|u2_Display/lt125_23  (
    .a({\u2_Display/n3901 ,\u2_Display/n3902 }),
    .b(2'b01),
    .fci(\u2_Display/lt125_c23 ),
    .fco(\u2_Display/lt125_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_26|u2_Display/lt125_25  (
    .a({\u2_Display/n3899 ,\u2_Display/n3900 }),
    .b(2'b10),
    .fci(\u2_Display/lt125_c25 ),
    .fco(\u2_Display/lt125_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_28|u2_Display/lt125_27  (
    .a({\u2_Display/n3897 ,\u2_Display/n3898 }),
    .b(2'b01),
    .fci(\u2_Display/lt125_c27 ),
    .fco(\u2_Display/lt125_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_2|u2_Display/lt125_1  (
    .a({\u2_Display/n3923 ,\u2_Display/n3924 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c1 ),
    .fco(\u2_Display/lt125_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_30|u2_Display/lt125_29  (
    .a({\u2_Display/n3895 ,\u2_Display/n3896 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c29 ),
    .fco(\u2_Display/lt125_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_4|u2_Display/lt125_3  (
    .a({\u2_Display/n3921 ,\u2_Display/n3922 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c3 ),
    .fco(\u2_Display/lt125_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_6|u2_Display/lt125_5  (
    .a({\u2_Display/n3919 ,\u2_Display/n3920 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c5 ),
    .fco(\u2_Display/lt125_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_8|u2_Display/lt125_7  (
    .a({\u2_Display/n3917 ,\u2_Display/n3918 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c7 ),
    .fco(\u2_Display/lt125_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_cout|u2_Display/lt125_31  (
    .a({1'b0,\u2_Display/n3894 }),
    .b(2'b10),
    .fci(\u2_Display/lt125_c31 ),
    .f({\u2_Display/n3926 ,open_n76390}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_0|u2_Display/lt126_cin  (
    .a({\u2_Display/n3960 ,1'b0}),
    .b({1'b0,open_n76396}),
    .fco(\u2_Display/lt126_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_10|u2_Display/lt126_9  (
    .a({\u2_Display/n3950 ,\u2_Display/n3951 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c9 ),
    .fco(\u2_Display/lt126_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_12|u2_Display/lt126_11  (
    .a({\u2_Display/n3948 ,\u2_Display/n3949 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c11 ),
    .fco(\u2_Display/lt126_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_14|u2_Display/lt126_13  (
    .a({\u2_Display/n3946 ,\u2_Display/n3947 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c13 ),
    .fco(\u2_Display/lt126_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_16|u2_Display/lt126_15  (
    .a({\u2_Display/n3944 ,\u2_Display/n3945 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c15 ),
    .fco(\u2_Display/lt126_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_18|u2_Display/lt126_17  (
    .a({\u2_Display/n3942 ,\u2_Display/n3943 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c17 ),
    .fco(\u2_Display/lt126_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_20|u2_Display/lt126_19  (
    .a({\u2_Display/n3940 ,\u2_Display/n3941 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c19 ),
    .fco(\u2_Display/lt126_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_22|u2_Display/lt126_21  (
    .a({\u2_Display/n3938 ,\u2_Display/n3939 }),
    .b(2'b10),
    .fci(\u2_Display/lt126_c21 ),
    .fco(\u2_Display/lt126_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_24|u2_Display/lt126_23  (
    .a({\u2_Display/n3936 ,\u2_Display/n3937 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c23 ),
    .fco(\u2_Display/lt126_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_26|u2_Display/lt126_25  (
    .a({\u2_Display/n3934 ,\u2_Display/n3935 }),
    .b(2'b11),
    .fci(\u2_Display/lt126_c25 ),
    .fco(\u2_Display/lt126_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_28|u2_Display/lt126_27  (
    .a({\u2_Display/n3932 ,\u2_Display/n3933 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c27 ),
    .fco(\u2_Display/lt126_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_2|u2_Display/lt126_1  (
    .a({\u2_Display/n3958 ,\u2_Display/n3959 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c1 ),
    .fco(\u2_Display/lt126_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_30|u2_Display/lt126_29  (
    .a({\u2_Display/n3930 ,\u2_Display/n3931 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c29 ),
    .fco(\u2_Display/lt126_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_4|u2_Display/lt126_3  (
    .a({\u2_Display/n3956 ,\u2_Display/n3957 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c3 ),
    .fco(\u2_Display/lt126_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_6|u2_Display/lt126_5  (
    .a({\u2_Display/n3954 ,\u2_Display/n3955 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c5 ),
    .fco(\u2_Display/lt126_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_8|u2_Display/lt126_7  (
    .a({\u2_Display/n3952 ,\u2_Display/n3953 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c7 ),
    .fco(\u2_Display/lt126_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_cout|u2_Display/lt126_31  (
    .a({1'b0,\u2_Display/n3929 }),
    .b(2'b10),
    .fci(\u2_Display/lt126_c31 ),
    .f({\u2_Display/n3961 ,open_n76800}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_0|u2_Display/lt127_cin  (
    .a({\u2_Display/n3995 ,1'b0}),
    .b({1'b0,open_n76806}),
    .fco(\u2_Display/lt127_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_10|u2_Display/lt127_9  (
    .a({\u2_Display/n3985 ,\u2_Display/n3986 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c9 ),
    .fco(\u2_Display/lt127_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_12|u2_Display/lt127_11  (
    .a({\u2_Display/n3983 ,\u2_Display/n3984 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c11 ),
    .fco(\u2_Display/lt127_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_14|u2_Display/lt127_13  (
    .a({\u2_Display/n3981 ,\u2_Display/n3982 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c13 ),
    .fco(\u2_Display/lt127_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_16|u2_Display/lt127_15  (
    .a({\u2_Display/n3979 ,\u2_Display/n3980 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c15 ),
    .fco(\u2_Display/lt127_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_18|u2_Display/lt127_17  (
    .a({\u2_Display/n3977 ,\u2_Display/n3978 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c17 ),
    .fco(\u2_Display/lt127_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_20|u2_Display/lt127_19  (
    .a({\u2_Display/n3975 ,\u2_Display/n3976 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c19 ),
    .fco(\u2_Display/lt127_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_22|u2_Display/lt127_21  (
    .a({\u2_Display/n3973 ,\u2_Display/n3974 }),
    .b(2'b01),
    .fci(\u2_Display/lt127_c21 ),
    .fco(\u2_Display/lt127_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_24|u2_Display/lt127_23  (
    .a({\u2_Display/n3971 ,\u2_Display/n3972 }),
    .b(2'b10),
    .fci(\u2_Display/lt127_c23 ),
    .fco(\u2_Display/lt127_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_26|u2_Display/lt127_25  (
    .a({\u2_Display/n3969 ,\u2_Display/n3970 }),
    .b(2'b01),
    .fci(\u2_Display/lt127_c25 ),
    .fco(\u2_Display/lt127_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_28|u2_Display/lt127_27  (
    .a({\u2_Display/n3967 ,\u2_Display/n3968 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c27 ),
    .fco(\u2_Display/lt127_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_2|u2_Display/lt127_1  (
    .a({\u2_Display/n3993 ,\u2_Display/n3994 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c1 ),
    .fco(\u2_Display/lt127_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_30|u2_Display/lt127_29  (
    .a({\u2_Display/n3965 ,\u2_Display/n3966 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c29 ),
    .fco(\u2_Display/lt127_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_4|u2_Display/lt127_3  (
    .a({\u2_Display/n3991 ,\u2_Display/n3992 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c3 ),
    .fco(\u2_Display/lt127_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_6|u2_Display/lt127_5  (
    .a({\u2_Display/n3989 ,\u2_Display/n3990 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c5 ),
    .fco(\u2_Display/lt127_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_8|u2_Display/lt127_7  (
    .a({\u2_Display/n3987 ,\u2_Display/n3988 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c7 ),
    .fco(\u2_Display/lt127_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_cout|u2_Display/lt127_31  (
    .a({1'b0,\u2_Display/n3964 }),
    .b(2'b10),
    .fci(\u2_Display/lt127_c31 ),
    .f({\u2_Display/n3996 ,open_n77210}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_0|u2_Display/lt128_cin  (
    .a({\u2_Display/n4030 ,1'b0}),
    .b({1'b0,open_n77216}),
    .fco(\u2_Display/lt128_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_10|u2_Display/lt128_9  (
    .a({\u2_Display/n4020 ,\u2_Display/n4021 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c9 ),
    .fco(\u2_Display/lt128_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_12|u2_Display/lt128_11  (
    .a({\u2_Display/n4018 ,\u2_Display/n4019 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c11 ),
    .fco(\u2_Display/lt128_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_14|u2_Display/lt128_13  (
    .a({\u2_Display/n4016 ,\u2_Display/n4017 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c13 ),
    .fco(\u2_Display/lt128_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_16|u2_Display/lt128_15  (
    .a({\u2_Display/n4014 ,\u2_Display/n4015 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c15 ),
    .fco(\u2_Display/lt128_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_18|u2_Display/lt128_17  (
    .a({\u2_Display/n4012 ,\u2_Display/n4013 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c17 ),
    .fco(\u2_Display/lt128_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_20|u2_Display/lt128_19  (
    .a({\u2_Display/n4010 ,\u2_Display/n4011 }),
    .b(2'b10),
    .fci(\u2_Display/lt128_c19 ),
    .fco(\u2_Display/lt128_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_22|u2_Display/lt128_21  (
    .a({\u2_Display/n4008 ,\u2_Display/n4009 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c21 ),
    .fco(\u2_Display/lt128_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_24|u2_Display/lt128_23  (
    .a({\u2_Display/n4006 ,\u2_Display/n4007 }),
    .b(2'b11),
    .fci(\u2_Display/lt128_c23 ),
    .fco(\u2_Display/lt128_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_26|u2_Display/lt128_25  (
    .a({\u2_Display/n4004 ,\u2_Display/n4005 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c25 ),
    .fco(\u2_Display/lt128_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_28|u2_Display/lt128_27  (
    .a({\u2_Display/n4002 ,\u2_Display/n4003 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c27 ),
    .fco(\u2_Display/lt128_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_2|u2_Display/lt128_1  (
    .a({\u2_Display/n4028 ,\u2_Display/n4029 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c1 ),
    .fco(\u2_Display/lt128_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_30|u2_Display/lt128_29  (
    .a({\u2_Display/n4000 ,\u2_Display/n4001 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c29 ),
    .fco(\u2_Display/lt128_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_4|u2_Display/lt128_3  (
    .a({\u2_Display/n4026 ,\u2_Display/n4027 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c3 ),
    .fco(\u2_Display/lt128_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_6|u2_Display/lt128_5  (
    .a({\u2_Display/n4024 ,\u2_Display/n4025 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c5 ),
    .fco(\u2_Display/lt128_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_8|u2_Display/lt128_7  (
    .a({\u2_Display/n4022 ,\u2_Display/n4023 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c7 ),
    .fco(\u2_Display/lt128_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_cout|u2_Display/lt128_31  (
    .a({1'b0,\u2_Display/n3999 }),
    .b(2'b10),
    .fci(\u2_Display/lt128_c31 ),
    .f({\u2_Display/n4031 ,open_n77620}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_0|u2_Display/lt129_cin  (
    .a({\u2_Display/n4065 ,1'b0}),
    .b({1'b0,open_n77626}),
    .fco(\u2_Display/lt129_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_10|u2_Display/lt129_9  (
    .a({\u2_Display/n4055 ,\u2_Display/n4056 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c9 ),
    .fco(\u2_Display/lt129_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_12|u2_Display/lt129_11  (
    .a({\u2_Display/n4053 ,\u2_Display/n4054 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c11 ),
    .fco(\u2_Display/lt129_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_14|u2_Display/lt129_13  (
    .a({\u2_Display/n4051 ,\u2_Display/n4052 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c13 ),
    .fco(\u2_Display/lt129_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_16|u2_Display/lt129_15  (
    .a({\u2_Display/n4049 ,\u2_Display/n4050 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c15 ),
    .fco(\u2_Display/lt129_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_18|u2_Display/lt129_17  (
    .a({\u2_Display/n4047 ,\u2_Display/n4048 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c17 ),
    .fco(\u2_Display/lt129_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_20|u2_Display/lt129_19  (
    .a({\u2_Display/n4045 ,\u2_Display/n4046 }),
    .b(2'b01),
    .fci(\u2_Display/lt129_c19 ),
    .fco(\u2_Display/lt129_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_22|u2_Display/lt129_21  (
    .a({\u2_Display/n4043 ,\u2_Display/n4044 }),
    .b(2'b10),
    .fci(\u2_Display/lt129_c21 ),
    .fco(\u2_Display/lt129_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_24|u2_Display/lt129_23  (
    .a({\u2_Display/n4041 ,\u2_Display/n4042 }),
    .b(2'b01),
    .fci(\u2_Display/lt129_c23 ),
    .fco(\u2_Display/lt129_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_26|u2_Display/lt129_25  (
    .a({\u2_Display/n4039 ,\u2_Display/n4040 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c25 ),
    .fco(\u2_Display/lt129_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_28|u2_Display/lt129_27  (
    .a({\u2_Display/n4037 ,\u2_Display/n4038 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c27 ),
    .fco(\u2_Display/lt129_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_2|u2_Display/lt129_1  (
    .a({\u2_Display/n4063 ,\u2_Display/n4064 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c1 ),
    .fco(\u2_Display/lt129_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_30|u2_Display/lt129_29  (
    .a({\u2_Display/n4035 ,\u2_Display/n4036 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c29 ),
    .fco(\u2_Display/lt129_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_4|u2_Display/lt129_3  (
    .a({\u2_Display/n4061 ,\u2_Display/n4062 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c3 ),
    .fco(\u2_Display/lt129_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_6|u2_Display/lt129_5  (
    .a({\u2_Display/n4059 ,\u2_Display/n4060 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c5 ),
    .fco(\u2_Display/lt129_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_8|u2_Display/lt129_7  (
    .a({\u2_Display/n4057 ,\u2_Display/n4058 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c7 ),
    .fco(\u2_Display/lt129_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_cout|u2_Display/lt129_31  (
    .a({1'b0,\u2_Display/n4034 }),
    .b(2'b10),
    .fci(\u2_Display/lt129_c31 ),
    .f({\u2_Display/n4066 ,open_n78030}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_0|u2_Display/lt130_cin  (
    .a({\u2_Display/n4100 ,1'b0}),
    .b({1'b0,open_n78036}),
    .fco(\u2_Display/lt130_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_10|u2_Display/lt130_9  (
    .a({\u2_Display/n4090 ,\u2_Display/n4091 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c9 ),
    .fco(\u2_Display/lt130_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_12|u2_Display/lt130_11  (
    .a({\u2_Display/n4088 ,\u2_Display/n4089 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c11 ),
    .fco(\u2_Display/lt130_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_14|u2_Display/lt130_13  (
    .a({\u2_Display/n4086 ,\u2_Display/n4087 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c13 ),
    .fco(\u2_Display/lt130_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_16|u2_Display/lt130_15  (
    .a({\u2_Display/n4084 ,\u2_Display/n4085 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c15 ),
    .fco(\u2_Display/lt130_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_18|u2_Display/lt130_17  (
    .a({\u2_Display/n4082 ,\u2_Display/n4083 }),
    .b(2'b10),
    .fci(\u2_Display/lt130_c17 ),
    .fco(\u2_Display/lt130_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_20|u2_Display/lt130_19  (
    .a({\u2_Display/n4080 ,\u2_Display/n4081 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c19 ),
    .fco(\u2_Display/lt130_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_22|u2_Display/lt130_21  (
    .a({\u2_Display/n4078 ,\u2_Display/n4079 }),
    .b(2'b11),
    .fci(\u2_Display/lt130_c21 ),
    .fco(\u2_Display/lt130_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_24|u2_Display/lt130_23  (
    .a({\u2_Display/n4076 ,\u2_Display/n4077 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c23 ),
    .fco(\u2_Display/lt130_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_26|u2_Display/lt130_25  (
    .a({\u2_Display/n4074 ,\u2_Display/n4075 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c25 ),
    .fco(\u2_Display/lt130_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_28|u2_Display/lt130_27  (
    .a({\u2_Display/n4072 ,\u2_Display/n4073 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c27 ),
    .fco(\u2_Display/lt130_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_2|u2_Display/lt130_1  (
    .a({\u2_Display/n4098 ,\u2_Display/n4099 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c1 ),
    .fco(\u2_Display/lt130_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_30|u2_Display/lt130_29  (
    .a({\u2_Display/n4070 ,\u2_Display/n4071 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c29 ),
    .fco(\u2_Display/lt130_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_4|u2_Display/lt130_3  (
    .a({\u2_Display/n4096 ,\u2_Display/n4097 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c3 ),
    .fco(\u2_Display/lt130_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_6|u2_Display/lt130_5  (
    .a({\u2_Display/n4094 ,\u2_Display/n4095 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c5 ),
    .fco(\u2_Display/lt130_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_8|u2_Display/lt130_7  (
    .a({\u2_Display/n4092 ,\u2_Display/n4093 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c7 ),
    .fco(\u2_Display/lt130_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_cout|u2_Display/lt130_31  (
    .a({1'b0,\u2_Display/n4069 }),
    .b(2'b10),
    .fci(\u2_Display/lt130_c31 ),
    .f({\u2_Display/n4101 ,open_n78440}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_0|u2_Display/lt131_cin  (
    .a({\u2_Display/n4135 ,1'b0}),
    .b({1'b0,open_n78446}),
    .fco(\u2_Display/lt131_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_10|u2_Display/lt131_9  (
    .a({\u2_Display/n4125 ,\u2_Display/n4126 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c9 ),
    .fco(\u2_Display/lt131_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_12|u2_Display/lt131_11  (
    .a({\u2_Display/n4123 ,\u2_Display/n4124 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c11 ),
    .fco(\u2_Display/lt131_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_14|u2_Display/lt131_13  (
    .a({\u2_Display/n4121 ,\u2_Display/n4122 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c13 ),
    .fco(\u2_Display/lt131_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_16|u2_Display/lt131_15  (
    .a({\u2_Display/n4119 ,\u2_Display/n4120 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c15 ),
    .fco(\u2_Display/lt131_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_18|u2_Display/lt131_17  (
    .a({\u2_Display/n4117 ,\u2_Display/n4118 }),
    .b(2'b01),
    .fci(\u2_Display/lt131_c17 ),
    .fco(\u2_Display/lt131_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_20|u2_Display/lt131_19  (
    .a({\u2_Display/n4115 ,\u2_Display/n4116 }),
    .b(2'b10),
    .fci(\u2_Display/lt131_c19 ),
    .fco(\u2_Display/lt131_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_22|u2_Display/lt131_21  (
    .a({\u2_Display/n4113 ,\u2_Display/n4114 }),
    .b(2'b01),
    .fci(\u2_Display/lt131_c21 ),
    .fco(\u2_Display/lt131_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_24|u2_Display/lt131_23  (
    .a({\u2_Display/n4111 ,\u2_Display/n4112 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c23 ),
    .fco(\u2_Display/lt131_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_26|u2_Display/lt131_25  (
    .a({\u2_Display/n4109 ,\u2_Display/n4110 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c25 ),
    .fco(\u2_Display/lt131_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_28|u2_Display/lt131_27  (
    .a({\u2_Display/n4107 ,\u2_Display/n4108 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c27 ),
    .fco(\u2_Display/lt131_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_2|u2_Display/lt131_1  (
    .a({\u2_Display/n4133 ,\u2_Display/n4134 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c1 ),
    .fco(\u2_Display/lt131_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_30|u2_Display/lt131_29  (
    .a({\u2_Display/n4105 ,\u2_Display/n4106 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c29 ),
    .fco(\u2_Display/lt131_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_4|u2_Display/lt131_3  (
    .a({\u2_Display/n4131 ,\u2_Display/n4132 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c3 ),
    .fco(\u2_Display/lt131_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_6|u2_Display/lt131_5  (
    .a({\u2_Display/n4129 ,\u2_Display/n4130 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c5 ),
    .fco(\u2_Display/lt131_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_8|u2_Display/lt131_7  (
    .a({\u2_Display/n4127 ,\u2_Display/n4128 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c7 ),
    .fco(\u2_Display/lt131_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_cout|u2_Display/lt131_31  (
    .a({1'b0,\u2_Display/n4104 }),
    .b(2'b10),
    .fci(\u2_Display/lt131_c31 ),
    .f({\u2_Display/n4136 ,open_n78850}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_0|u2_Display/lt132_cin  (
    .a({\u2_Display/n4170 ,1'b0}),
    .b({1'b0,open_n78856}),
    .fco(\u2_Display/lt132_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_10|u2_Display/lt132_9  (
    .a({\u2_Display/n4160 ,\u2_Display/n4161 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c9 ),
    .fco(\u2_Display/lt132_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_12|u2_Display/lt132_11  (
    .a({\u2_Display/n4158 ,\u2_Display/n4159 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c11 ),
    .fco(\u2_Display/lt132_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_14|u2_Display/lt132_13  (
    .a({\u2_Display/n4156 ,\u2_Display/n4157 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c13 ),
    .fco(\u2_Display/lt132_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_16|u2_Display/lt132_15  (
    .a({\u2_Display/n4154 ,\u2_Display/n4155 }),
    .b(2'b10),
    .fci(\u2_Display/lt132_c15 ),
    .fco(\u2_Display/lt132_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_18|u2_Display/lt132_17  (
    .a({\u2_Display/n4152 ,\u2_Display/n4153 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c17 ),
    .fco(\u2_Display/lt132_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_20|u2_Display/lt132_19  (
    .a({\u2_Display/n4150 ,\u2_Display/n4151 }),
    .b(2'b11),
    .fci(\u2_Display/lt132_c19 ),
    .fco(\u2_Display/lt132_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_22|u2_Display/lt132_21  (
    .a({\u2_Display/n4148 ,\u2_Display/n4149 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c21 ),
    .fco(\u2_Display/lt132_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_24|u2_Display/lt132_23  (
    .a({\u2_Display/n4146 ,\u2_Display/n4147 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c23 ),
    .fco(\u2_Display/lt132_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_26|u2_Display/lt132_25  (
    .a({\u2_Display/n4144 ,\u2_Display/n4145 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c25 ),
    .fco(\u2_Display/lt132_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_28|u2_Display/lt132_27  (
    .a({\u2_Display/n4142 ,\u2_Display/n4143 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c27 ),
    .fco(\u2_Display/lt132_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_2|u2_Display/lt132_1  (
    .a({\u2_Display/n4168 ,\u2_Display/n4169 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c1 ),
    .fco(\u2_Display/lt132_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_30|u2_Display/lt132_29  (
    .a({\u2_Display/n4140 ,\u2_Display/n4141 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c29 ),
    .fco(\u2_Display/lt132_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_4|u2_Display/lt132_3  (
    .a({\u2_Display/n4166 ,\u2_Display/n4167 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c3 ),
    .fco(\u2_Display/lt132_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_6|u2_Display/lt132_5  (
    .a({\u2_Display/n4164 ,\u2_Display/n4165 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c5 ),
    .fco(\u2_Display/lt132_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_8|u2_Display/lt132_7  (
    .a({\u2_Display/n4162 ,\u2_Display/n4163 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c7 ),
    .fco(\u2_Display/lt132_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_cout|u2_Display/lt132_31  (
    .a({1'b0,\u2_Display/n4139 }),
    .b(2'b10),
    .fci(\u2_Display/lt132_c31 ),
    .f({\u2_Display/n4171 ,open_n79260}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_0|u2_Display/lt133_cin  (
    .a({\u2_Display/n4205 ,1'b0}),
    .b({1'b0,open_n79266}),
    .fco(\u2_Display/lt133_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_10|u2_Display/lt133_9  (
    .a({\u2_Display/n4195 ,\u2_Display/n4196 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c9 ),
    .fco(\u2_Display/lt133_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_12|u2_Display/lt133_11  (
    .a({\u2_Display/n4193 ,\u2_Display/n4194 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c11 ),
    .fco(\u2_Display/lt133_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_14|u2_Display/lt133_13  (
    .a({\u2_Display/n4191 ,\u2_Display/n4192 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c13 ),
    .fco(\u2_Display/lt133_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_16|u2_Display/lt133_15  (
    .a({\u2_Display/n4189 ,\u2_Display/n4190 }),
    .b(2'b01),
    .fci(\u2_Display/lt133_c15 ),
    .fco(\u2_Display/lt133_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_18|u2_Display/lt133_17  (
    .a({\u2_Display/n4187 ,\u2_Display/n4188 }),
    .b(2'b10),
    .fci(\u2_Display/lt133_c17 ),
    .fco(\u2_Display/lt133_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_20|u2_Display/lt133_19  (
    .a({\u2_Display/n4185 ,\u2_Display/n4186 }),
    .b(2'b01),
    .fci(\u2_Display/lt133_c19 ),
    .fco(\u2_Display/lt133_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_22|u2_Display/lt133_21  (
    .a({\u2_Display/n4183 ,\u2_Display/n4184 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c21 ),
    .fco(\u2_Display/lt133_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_24|u2_Display/lt133_23  (
    .a({\u2_Display/n4181 ,\u2_Display/n4182 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c23 ),
    .fco(\u2_Display/lt133_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_26|u2_Display/lt133_25  (
    .a({\u2_Display/n4179 ,\u2_Display/n4180 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c25 ),
    .fco(\u2_Display/lt133_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_28|u2_Display/lt133_27  (
    .a({\u2_Display/n4177 ,\u2_Display/n4178 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c27 ),
    .fco(\u2_Display/lt133_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_2|u2_Display/lt133_1  (
    .a({\u2_Display/n4203 ,\u2_Display/n4204 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c1 ),
    .fco(\u2_Display/lt133_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_30|u2_Display/lt133_29  (
    .a({\u2_Display/n4175 ,\u2_Display/n4176 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c29 ),
    .fco(\u2_Display/lt133_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_4|u2_Display/lt133_3  (
    .a({\u2_Display/n4201 ,\u2_Display/n4202 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c3 ),
    .fco(\u2_Display/lt133_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_6|u2_Display/lt133_5  (
    .a({\u2_Display/n4199 ,\u2_Display/n4200 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c5 ),
    .fco(\u2_Display/lt133_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_8|u2_Display/lt133_7  (
    .a({\u2_Display/n4197 ,\u2_Display/n4198 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c7 ),
    .fco(\u2_Display/lt133_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_cout|u2_Display/lt133_31  (
    .a({1'b0,\u2_Display/n4174 }),
    .b(2'b10),
    .fci(\u2_Display/lt133_c31 ),
    .f({\u2_Display/n4206 ,open_n79670}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_0|u2_Display/lt134_cin  (
    .a({\u2_Display/n4240 ,1'b0}),
    .b({1'b0,open_n79676}),
    .fco(\u2_Display/lt134_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_10|u2_Display/lt134_9  (
    .a({\u2_Display/n4230 ,\u2_Display/n4231 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c9 ),
    .fco(\u2_Display/lt134_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_12|u2_Display/lt134_11  (
    .a({\u2_Display/n4228 ,\u2_Display/n4229 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c11 ),
    .fco(\u2_Display/lt134_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_14|u2_Display/lt134_13  (
    .a({\u2_Display/n4226 ,\u2_Display/n4227 }),
    .b(2'b10),
    .fci(\u2_Display/lt134_c13 ),
    .fco(\u2_Display/lt134_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_16|u2_Display/lt134_15  (
    .a({\u2_Display/n4224 ,\u2_Display/n4225 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c15 ),
    .fco(\u2_Display/lt134_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_18|u2_Display/lt134_17  (
    .a({\u2_Display/n4222 ,\u2_Display/n4223 }),
    .b(2'b11),
    .fci(\u2_Display/lt134_c17 ),
    .fco(\u2_Display/lt134_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_20|u2_Display/lt134_19  (
    .a({\u2_Display/n4220 ,\u2_Display/n4221 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c19 ),
    .fco(\u2_Display/lt134_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_22|u2_Display/lt134_21  (
    .a({\u2_Display/n4218 ,\u2_Display/n4219 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c21 ),
    .fco(\u2_Display/lt134_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_24|u2_Display/lt134_23  (
    .a({\u2_Display/n4216 ,\u2_Display/n4217 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c23 ),
    .fco(\u2_Display/lt134_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_26|u2_Display/lt134_25  (
    .a({\u2_Display/n4214 ,\u2_Display/n4215 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c25 ),
    .fco(\u2_Display/lt134_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_28|u2_Display/lt134_27  (
    .a({\u2_Display/n4212 ,\u2_Display/n4213 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c27 ),
    .fco(\u2_Display/lt134_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_2|u2_Display/lt134_1  (
    .a({\u2_Display/n4238 ,\u2_Display/n4239 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c1 ),
    .fco(\u2_Display/lt134_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_30|u2_Display/lt134_29  (
    .a({\u2_Display/n4210 ,\u2_Display/n4211 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c29 ),
    .fco(\u2_Display/lt134_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_4|u2_Display/lt134_3  (
    .a({\u2_Display/n4236 ,\u2_Display/n4237 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c3 ),
    .fco(\u2_Display/lt134_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_6|u2_Display/lt134_5  (
    .a({\u2_Display/n4234 ,\u2_Display/n4235 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c5 ),
    .fco(\u2_Display/lt134_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_8|u2_Display/lt134_7  (
    .a({\u2_Display/n4232 ,\u2_Display/n4233 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c7 ),
    .fco(\u2_Display/lt134_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_cout|u2_Display/lt134_31  (
    .a({1'b0,\u2_Display/n4209 }),
    .b(2'b10),
    .fci(\u2_Display/lt134_c31 ),
    .f({\u2_Display/n4241 ,open_n80080}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_0|u2_Display/lt135_cin  (
    .a({\u2_Display/n4275 ,1'b0}),
    .b({1'b0,open_n80086}),
    .fco(\u2_Display/lt135_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_10|u2_Display/lt135_9  (
    .a({\u2_Display/n4265 ,\u2_Display/n4266 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c9 ),
    .fco(\u2_Display/lt135_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_12|u2_Display/lt135_11  (
    .a({\u2_Display/n4263 ,\u2_Display/n4264 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c11 ),
    .fco(\u2_Display/lt135_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_14|u2_Display/lt135_13  (
    .a({\u2_Display/n4261 ,\u2_Display/n4262 }),
    .b(2'b01),
    .fci(\u2_Display/lt135_c13 ),
    .fco(\u2_Display/lt135_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_16|u2_Display/lt135_15  (
    .a({\u2_Display/n4259 ,\u2_Display/n4260 }),
    .b(2'b10),
    .fci(\u2_Display/lt135_c15 ),
    .fco(\u2_Display/lt135_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_18|u2_Display/lt135_17  (
    .a({\u2_Display/n4257 ,\u2_Display/n4258 }),
    .b(2'b01),
    .fci(\u2_Display/lt135_c17 ),
    .fco(\u2_Display/lt135_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_20|u2_Display/lt135_19  (
    .a({\u2_Display/n4255 ,\u2_Display/n4256 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c19 ),
    .fco(\u2_Display/lt135_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_22|u2_Display/lt135_21  (
    .a({\u2_Display/n4253 ,\u2_Display/n4254 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c21 ),
    .fco(\u2_Display/lt135_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_24|u2_Display/lt135_23  (
    .a({\u2_Display/n4251 ,\u2_Display/n4252 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c23 ),
    .fco(\u2_Display/lt135_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_26|u2_Display/lt135_25  (
    .a({\u2_Display/n4249 ,\u2_Display/n4250 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c25 ),
    .fco(\u2_Display/lt135_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_28|u2_Display/lt135_27  (
    .a({\u2_Display/n4247 ,\u2_Display/n4248 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c27 ),
    .fco(\u2_Display/lt135_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_2|u2_Display/lt135_1  (
    .a({\u2_Display/n4273 ,\u2_Display/n4274 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c1 ),
    .fco(\u2_Display/lt135_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_30|u2_Display/lt135_29  (
    .a({\u2_Display/n4245 ,\u2_Display/n4246 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c29 ),
    .fco(\u2_Display/lt135_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_4|u2_Display/lt135_3  (
    .a({\u2_Display/n4271 ,\u2_Display/n4272 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c3 ),
    .fco(\u2_Display/lt135_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_6|u2_Display/lt135_5  (
    .a({\u2_Display/n4269 ,\u2_Display/n4270 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c5 ),
    .fco(\u2_Display/lt135_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_8|u2_Display/lt135_7  (
    .a({\u2_Display/n4267 ,\u2_Display/n4268 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c7 ),
    .fco(\u2_Display/lt135_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_cout|u2_Display/lt135_31  (
    .a({1'b0,\u2_Display/n4244 }),
    .b(2'b10),
    .fci(\u2_Display/lt135_c31 ),
    .f({\u2_Display/n4276 ,open_n80490}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_0|u2_Display/lt136_cin  (
    .a({\u2_Display/n4310 ,1'b0}),
    .b({1'b0,open_n80496}),
    .fco(\u2_Display/lt136_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_10|u2_Display/lt136_9  (
    .a({\u2_Display/n4300 ,\u2_Display/n4301 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c9 ),
    .fco(\u2_Display/lt136_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_12|u2_Display/lt136_11  (
    .a({\u2_Display/n4298 ,\u2_Display/n4299 }),
    .b(2'b10),
    .fci(\u2_Display/lt136_c11 ),
    .fco(\u2_Display/lt136_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_14|u2_Display/lt136_13  (
    .a({\u2_Display/n4296 ,\u2_Display/n4297 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c13 ),
    .fco(\u2_Display/lt136_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_16|u2_Display/lt136_15  (
    .a({\u2_Display/n4294 ,\u2_Display/n4295 }),
    .b(2'b11),
    .fci(\u2_Display/lt136_c15 ),
    .fco(\u2_Display/lt136_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_18|u2_Display/lt136_17  (
    .a({\u2_Display/n4292 ,\u2_Display/n4293 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c17 ),
    .fco(\u2_Display/lt136_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_20|u2_Display/lt136_19  (
    .a({\u2_Display/n4290 ,\u2_Display/n4291 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c19 ),
    .fco(\u2_Display/lt136_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_22|u2_Display/lt136_21  (
    .a({\u2_Display/n4288 ,\u2_Display/n4289 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c21 ),
    .fco(\u2_Display/lt136_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_24|u2_Display/lt136_23  (
    .a({\u2_Display/n4286 ,\u2_Display/n4287 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c23 ),
    .fco(\u2_Display/lt136_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_26|u2_Display/lt136_25  (
    .a({\u2_Display/n4284 ,\u2_Display/n4285 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c25 ),
    .fco(\u2_Display/lt136_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_28|u2_Display/lt136_27  (
    .a({\u2_Display/n4282 ,\u2_Display/n4283 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c27 ),
    .fco(\u2_Display/lt136_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_2|u2_Display/lt136_1  (
    .a({\u2_Display/n4308 ,\u2_Display/n4309 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c1 ),
    .fco(\u2_Display/lt136_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_30|u2_Display/lt136_29  (
    .a({\u2_Display/n4280 ,\u2_Display/n4281 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c29 ),
    .fco(\u2_Display/lt136_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_4|u2_Display/lt136_3  (
    .a({\u2_Display/n4306 ,\u2_Display/n4307 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c3 ),
    .fco(\u2_Display/lt136_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_6|u2_Display/lt136_5  (
    .a({\u2_Display/n4304 ,\u2_Display/n4305 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c5 ),
    .fco(\u2_Display/lt136_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_8|u2_Display/lt136_7  (
    .a({\u2_Display/n4302 ,\u2_Display/n4303 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c7 ),
    .fco(\u2_Display/lt136_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_cout|u2_Display/lt136_31  (
    .a({1'b0,\u2_Display/n4279 }),
    .b(2'b10),
    .fci(\u2_Display/lt136_c31 ),
    .f({\u2_Display/n4311 ,open_n80900}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/lt137_0|u2_Display/lt137_cin  (
    .a({\u2_Display/n4345 ,1'b0}),
    .b({1'b0,open_n80906}),
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .mi(\u2_Display/n41 [31:30]),
    .fco(\u2_Display/lt137_c1 ),
    .q(\u2_Display/counta [31:30]));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_10|u2_Display/lt137_9  (
    .a({\u2_Display/n4335 ,\u2_Display/n4336 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c9 ),
    .fco(\u2_Display/lt137_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_12|u2_Display/lt137_11  (
    .a({\u2_Display/n4333 ,\u2_Display/n4334 }),
    .b(2'b01),
    .fci(\u2_Display/lt137_c11 ),
    .fco(\u2_Display/lt137_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_14|u2_Display/lt137_13  (
    .a({\u2_Display/n4331 ,\u2_Display/n4332 }),
    .b(2'b10),
    .fci(\u2_Display/lt137_c13 ),
    .fco(\u2_Display/lt137_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_16|u2_Display/lt137_15  (
    .a({\u2_Display/n4329 ,\u2_Display/n4330 }),
    .b(2'b01),
    .fci(\u2_Display/lt137_c15 ),
    .fco(\u2_Display/lt137_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_18|u2_Display/lt137_17  (
    .a({\u2_Display/n4327 ,\u2_Display/n4328 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c17 ),
    .fco(\u2_Display/lt137_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_20|u2_Display/lt137_19  (
    .a({\u2_Display/n4325 ,\u2_Display/n4326 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c19 ),
    .fco(\u2_Display/lt137_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_22|u2_Display/lt137_21  (
    .a({\u2_Display/n4323 ,\u2_Display/n4324 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c21 ),
    .fco(\u2_Display/lt137_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_24|u2_Display/lt137_23  (
    .a({\u2_Display/n4321 ,\u2_Display/n4322 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c23 ),
    .fco(\u2_Display/lt137_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_26|u2_Display/lt137_25  (
    .a({\u2_Display/n4319 ,\u2_Display/n4320 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c25 ),
    .fco(\u2_Display/lt137_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_28|u2_Display/lt137_27  (
    .a({\u2_Display/n4317 ,\u2_Display/n4318 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c27 ),
    .fco(\u2_Display/lt137_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_2|u2_Display/lt137_1  (
    .a({\u2_Display/n4343 ,\u2_Display/n4344 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c1 ),
    .fco(\u2_Display/lt137_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_30|u2_Display/lt137_29  (
    .a({\u2_Display/n4315 ,\u2_Display/n4316 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c29 ),
    .fco(\u2_Display/lt137_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_4|u2_Display/lt137_3  (
    .a({\u2_Display/n4341 ,\u2_Display/n4342 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c3 ),
    .fco(\u2_Display/lt137_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_6|u2_Display/lt137_5  (
    .a({\u2_Display/n4339 ,\u2_Display/n4340 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c5 ),
    .fco(\u2_Display/lt137_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_8|u2_Display/lt137_7  (
    .a({\u2_Display/n4337 ,\u2_Display/n4338 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c7 ),
    .fco(\u2_Display/lt137_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_cout|u2_Display/lt137_31  (
    .a({1'b0,\u2_Display/n4314 }),
    .b(2'b10),
    .fci(\u2_Display/lt137_c31 ),
    .f({\u2_Display/n4346 ,open_n81304}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_0|u2_Display/lt138_cin  (
    .a({\u2_Display/n4380 ,1'b0}),
    .b({1'b0,open_n81310}),
    .fco(\u2_Display/lt138_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_10|u2_Display/lt138_9  (
    .a({\u2_Display/n4370 ,\u2_Display/n4371 }),
    .b(2'b10),
    .fci(\u2_Display/lt138_c9 ),
    .fco(\u2_Display/lt138_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_12|u2_Display/lt138_11  (
    .a({\u2_Display/n4368 ,\u2_Display/n4369 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c11 ),
    .fco(\u2_Display/lt138_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_14|u2_Display/lt138_13  (
    .a({\u2_Display/n4366 ,\u2_Display/n4367 }),
    .b(2'b11),
    .fci(\u2_Display/lt138_c13 ),
    .fco(\u2_Display/lt138_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_16|u2_Display/lt138_15  (
    .a({\u2_Display/n4364 ,\u2_Display/n4365 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c15 ),
    .fco(\u2_Display/lt138_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_18|u2_Display/lt138_17  (
    .a({\u2_Display/n4362 ,\u2_Display/n4363 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c17 ),
    .fco(\u2_Display/lt138_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_20|u2_Display/lt138_19  (
    .a({\u2_Display/n4360 ,\u2_Display/n4361 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c19 ),
    .fco(\u2_Display/lt138_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_22|u2_Display/lt138_21  (
    .a({\u2_Display/n4358 ,\u2_Display/n4359 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c21 ),
    .fco(\u2_Display/lt138_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_24|u2_Display/lt138_23  (
    .a({\u2_Display/n4356 ,\u2_Display/n4357 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c23 ),
    .fco(\u2_Display/lt138_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_26|u2_Display/lt138_25  (
    .a({\u2_Display/n4354 ,\u2_Display/n4355 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c25 ),
    .fco(\u2_Display/lt138_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_28|u2_Display/lt138_27  (
    .a({\u2_Display/n4352 ,\u2_Display/n4353 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c27 ),
    .fco(\u2_Display/lt138_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_2|u2_Display/lt138_1  (
    .a({\u2_Display/n4378 ,\u2_Display/n4379 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c1 ),
    .fco(\u2_Display/lt138_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_30|u2_Display/lt138_29  (
    .a({\u2_Display/n4350 ,\u2_Display/n4351 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c29 ),
    .fco(\u2_Display/lt138_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_4|u2_Display/lt138_3  (
    .a({\u2_Display/n4376 ,\u2_Display/n4377 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c3 ),
    .fco(\u2_Display/lt138_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_6|u2_Display/lt138_5  (
    .a({\u2_Display/n4374 ,\u2_Display/n4375 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c5 ),
    .fco(\u2_Display/lt138_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_8|u2_Display/lt138_7  (
    .a({\u2_Display/n4372 ,\u2_Display/n4373 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c7 ),
    .fco(\u2_Display/lt138_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_cout|u2_Display/lt138_31  (
    .a({1'b0,\u2_Display/n4349 }),
    .b(2'b10),
    .fci(\u2_Display/lt138_c31 ),
    .f({\u2_Display/n4381 ,open_n81714}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_0|u2_Display/lt139_cin  (
    .a({\u2_Display/n4415 ,1'b0}),
    .b({1'b0,open_n81720}),
    .fco(\u2_Display/lt139_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_10|u2_Display/lt139_9  (
    .a({\u2_Display/n4405 ,\u2_Display/n4406 }),
    .b(2'b01),
    .fci(\u2_Display/lt139_c9 ),
    .fco(\u2_Display/lt139_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_12|u2_Display/lt139_11  (
    .a({\u2_Display/n4403 ,\u2_Display/n4404 }),
    .b(2'b10),
    .fci(\u2_Display/lt139_c11 ),
    .fco(\u2_Display/lt139_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_14|u2_Display/lt139_13  (
    .a({\u2_Display/n4401 ,\u2_Display/n4402 }),
    .b(2'b01),
    .fci(\u2_Display/lt139_c13 ),
    .fco(\u2_Display/lt139_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_16|u2_Display/lt139_15  (
    .a({\u2_Display/n4399 ,\u2_Display/n4400 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c15 ),
    .fco(\u2_Display/lt139_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_18|u2_Display/lt139_17  (
    .a({\u2_Display/n4397 ,\u2_Display/n4398 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c17 ),
    .fco(\u2_Display/lt139_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_20|u2_Display/lt139_19  (
    .a({\u2_Display/n4395 ,\u2_Display/n4396 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c19 ),
    .fco(\u2_Display/lt139_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_22|u2_Display/lt139_21  (
    .a({\u2_Display/n4393 ,\u2_Display/n4394 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c21 ),
    .fco(\u2_Display/lt139_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_24|u2_Display/lt139_23  (
    .a({\u2_Display/n4391 ,\u2_Display/n4392 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c23 ),
    .fco(\u2_Display/lt139_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_26|u2_Display/lt139_25  (
    .a({\u2_Display/n4389 ,\u2_Display/n4390 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c25 ),
    .fco(\u2_Display/lt139_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_28|u2_Display/lt139_27  (
    .a({\u2_Display/n4387 ,\u2_Display/n4388 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c27 ),
    .fco(\u2_Display/lt139_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_2|u2_Display/lt139_1  (
    .a({\u2_Display/n4413 ,\u2_Display/n4414 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c1 ),
    .fco(\u2_Display/lt139_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_30|u2_Display/lt139_29  (
    .a({\u2_Display/n4385 ,\u2_Display/n4386 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c29 ),
    .fco(\u2_Display/lt139_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_4|u2_Display/lt139_3  (
    .a({\u2_Display/n4411 ,\u2_Display/n4412 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c3 ),
    .fco(\u2_Display/lt139_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_6|u2_Display/lt139_5  (
    .a({\u2_Display/n4409 ,\u2_Display/n4410 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c5 ),
    .fco(\u2_Display/lt139_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_8|u2_Display/lt139_7  (
    .a({\u2_Display/n4407 ,\u2_Display/n4408 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c7 ),
    .fco(\u2_Display/lt139_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_cout|u2_Display/lt139_31  (
    .a({1'b0,\u2_Display/n4384 }),
    .b(2'b10),
    .fci(\u2_Display/lt139_c31 ),
    .f({\u2_Display/n4416 ,open_n82124}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_0|u2_Display/lt140_cin  (
    .a({\u2_Display/n4450 ,1'b0}),
    .b({1'b0,open_n82130}),
    .fco(\u2_Display/lt140_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_10|u2_Display/lt140_9  (
    .a({\u2_Display/n4440 ,\u2_Display/n4441 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c9 ),
    .fco(\u2_Display/lt140_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_12|u2_Display/lt140_11  (
    .a({\u2_Display/n4438 ,\u2_Display/n4439 }),
    .b(2'b11),
    .fci(\u2_Display/lt140_c11 ),
    .fco(\u2_Display/lt140_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_14|u2_Display/lt140_13  (
    .a({\u2_Display/n4436 ,\u2_Display/n4437 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c13 ),
    .fco(\u2_Display/lt140_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_16|u2_Display/lt140_15  (
    .a({\u2_Display/n4434 ,\u2_Display/n4435 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c15 ),
    .fco(\u2_Display/lt140_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_18|u2_Display/lt140_17  (
    .a({\u2_Display/n4432 ,\u2_Display/n4433 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c17 ),
    .fco(\u2_Display/lt140_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_20|u2_Display/lt140_19  (
    .a({\u2_Display/n4430 ,\u2_Display/n4431 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c19 ),
    .fco(\u2_Display/lt140_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_22|u2_Display/lt140_21  (
    .a({\u2_Display/n4428 ,\u2_Display/n4429 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c21 ),
    .fco(\u2_Display/lt140_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_24|u2_Display/lt140_23  (
    .a({\u2_Display/n4426 ,\u2_Display/n4427 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c23 ),
    .fco(\u2_Display/lt140_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_26|u2_Display/lt140_25  (
    .a({\u2_Display/n4424 ,\u2_Display/n4425 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c25 ),
    .fco(\u2_Display/lt140_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_28|u2_Display/lt140_27  (
    .a({\u2_Display/n4422 ,\u2_Display/n4423 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c27 ),
    .fco(\u2_Display/lt140_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_2|u2_Display/lt140_1  (
    .a({\u2_Display/n4448 ,\u2_Display/n4449 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c1 ),
    .fco(\u2_Display/lt140_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_30|u2_Display/lt140_29  (
    .a({\u2_Display/n4420 ,\u2_Display/n4421 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c29 ),
    .fco(\u2_Display/lt140_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_4|u2_Display/lt140_3  (
    .a({\u2_Display/n4446 ,\u2_Display/n4447 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c3 ),
    .fco(\u2_Display/lt140_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_6|u2_Display/lt140_5  (
    .a({\u2_Display/n4444 ,\u2_Display/n4445 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c5 ),
    .fco(\u2_Display/lt140_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_8|u2_Display/lt140_7  (
    .a({\u2_Display/n4442 ,\u2_Display/n4443 }),
    .b(2'b10),
    .fci(\u2_Display/lt140_c7 ),
    .fco(\u2_Display/lt140_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_cout|u2_Display/lt140_31  (
    .a({1'b0,\u2_Display/n4419 }),
    .b(2'b10),
    .fci(\u2_Display/lt140_c31 ),
    .f({\u2_Display/n4451 ,open_n82534}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_0|u2_Display/lt141_cin  (
    .a({\u2_Display/n4485 ,1'b0}),
    .b({1'b0,open_n82540}),
    .fco(\u2_Display/lt141_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_10|u2_Display/lt141_9  (
    .a({\u2_Display/n4475 ,\u2_Display/n4476 }),
    .b(2'b10),
    .fci(\u2_Display/lt141_c9 ),
    .fco(\u2_Display/lt141_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_12|u2_Display/lt141_11  (
    .a({\u2_Display/n4473 ,\u2_Display/n4474 }),
    .b(2'b01),
    .fci(\u2_Display/lt141_c11 ),
    .fco(\u2_Display/lt141_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_14|u2_Display/lt141_13  (
    .a({\u2_Display/n4471 ,\u2_Display/n4472 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c13 ),
    .fco(\u2_Display/lt141_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_16|u2_Display/lt141_15  (
    .a({\u2_Display/n4469 ,\u2_Display/n4470 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c15 ),
    .fco(\u2_Display/lt141_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_18|u2_Display/lt141_17  (
    .a({\u2_Display/n4467 ,\u2_Display/n4468 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c17 ),
    .fco(\u2_Display/lt141_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_20|u2_Display/lt141_19  (
    .a({\u2_Display/n4465 ,\u2_Display/n4466 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c19 ),
    .fco(\u2_Display/lt141_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_22|u2_Display/lt141_21  (
    .a({\u2_Display/n4463 ,\u2_Display/n4464 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c21 ),
    .fco(\u2_Display/lt141_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_24|u2_Display/lt141_23  (
    .a({\u2_Display/n4461 ,\u2_Display/n4462 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c23 ),
    .fco(\u2_Display/lt141_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_26|u2_Display/lt141_25  (
    .a({\u2_Display/n4459 ,\u2_Display/n4460 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c25 ),
    .fco(\u2_Display/lt141_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_28|u2_Display/lt141_27  (
    .a({\u2_Display/n4457 ,\u2_Display/n4458 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c27 ),
    .fco(\u2_Display/lt141_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_2|u2_Display/lt141_1  (
    .a({\u2_Display/n4483 ,\u2_Display/n4484 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c1 ),
    .fco(\u2_Display/lt141_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_30|u2_Display/lt141_29  (
    .a({\u2_Display/n4455 ,\u2_Display/n4456 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c29 ),
    .fco(\u2_Display/lt141_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_4|u2_Display/lt141_3  (
    .a({\u2_Display/n4481 ,\u2_Display/n4482 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c3 ),
    .fco(\u2_Display/lt141_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_6|u2_Display/lt141_5  (
    .a({\u2_Display/n4479 ,\u2_Display/n4480 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c5 ),
    .fco(\u2_Display/lt141_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_8|u2_Display/lt141_7  (
    .a({\u2_Display/n4477 ,\u2_Display/n4478 }),
    .b(2'b01),
    .fci(\u2_Display/lt141_c7 ),
    .fco(\u2_Display/lt141_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_cout|u2_Display/lt141_31  (
    .a({1'b0,\u2_Display/n4454 }),
    .b(2'b10),
    .fci(\u2_Display/lt141_c31 ),
    .f({\u2_Display/n4486 ,open_n82944}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_0|u2_Display/lt142_cin  (
    .a({\u2_Display/n4520 ,1'b0}),
    .b({1'b0,open_n82950}),
    .fco(\u2_Display/lt142_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_10|u2_Display/lt142_9  (
    .a({\u2_Display/n4510 ,\u2_Display/n4511 }),
    .b(2'b11),
    .fci(\u2_Display/lt142_c9 ),
    .fco(\u2_Display/lt142_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_12|u2_Display/lt142_11  (
    .a({\u2_Display/n4508 ,\u2_Display/n4509 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c11 ),
    .fco(\u2_Display/lt142_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_14|u2_Display/lt142_13  (
    .a({\u2_Display/n4506 ,\u2_Display/n4507 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c13 ),
    .fco(\u2_Display/lt142_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_16|u2_Display/lt142_15  (
    .a({\u2_Display/n4504 ,\u2_Display/n4505 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c15 ),
    .fco(\u2_Display/lt142_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_18|u2_Display/lt142_17  (
    .a({\u2_Display/n4502 ,\u2_Display/n4503 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c17 ),
    .fco(\u2_Display/lt142_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_20|u2_Display/lt142_19  (
    .a({\u2_Display/n4500 ,\u2_Display/n4501 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c19 ),
    .fco(\u2_Display/lt142_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_22|u2_Display/lt142_21  (
    .a({\u2_Display/n4498 ,\u2_Display/n4499 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c21 ),
    .fco(\u2_Display/lt142_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_24|u2_Display/lt142_23  (
    .a({\u2_Display/n4496 ,\u2_Display/n4497 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c23 ),
    .fco(\u2_Display/lt142_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_26|u2_Display/lt142_25  (
    .a({\u2_Display/n4494 ,\u2_Display/n4495 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c25 ),
    .fco(\u2_Display/lt142_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_28|u2_Display/lt142_27  (
    .a({\u2_Display/n4492 ,\u2_Display/n4493 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c27 ),
    .fco(\u2_Display/lt142_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_2|u2_Display/lt142_1  (
    .a({\u2_Display/n4518 ,\u2_Display/n4519 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c1 ),
    .fco(\u2_Display/lt142_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_30|u2_Display/lt142_29  (
    .a({\u2_Display/n4490 ,\u2_Display/n4491 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c29 ),
    .fco(\u2_Display/lt142_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_4|u2_Display/lt142_3  (
    .a({\u2_Display/n4516 ,\u2_Display/n4517 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c3 ),
    .fco(\u2_Display/lt142_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_6|u2_Display/lt142_5  (
    .a({\u2_Display/n4514 ,\u2_Display/n4515 }),
    .b(2'b10),
    .fci(\u2_Display/lt142_c5 ),
    .fco(\u2_Display/lt142_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_8|u2_Display/lt142_7  (
    .a({\u2_Display/n4512 ,\u2_Display/n4513 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c7 ),
    .fco(\u2_Display/lt142_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_cout|u2_Display/lt142_31  (
    .a({1'b0,\u2_Display/n4489 }),
    .b(2'b10),
    .fci(\u2_Display/lt142_c31 ),
    .f({\u2_Display/n4521 ,open_n83354}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_0|u2_Display/lt143_cin  (
    .a({\u2_Display/n4555 ,1'b0}),
    .b({1'b0,open_n83360}),
    .fco(\u2_Display/lt143_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_10|u2_Display/lt143_9  (
    .a({\u2_Display/n4545 ,\u2_Display/n4546 }),
    .b(2'b01),
    .fci(\u2_Display/lt143_c9 ),
    .fco(\u2_Display/lt143_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_12|u2_Display/lt143_11  (
    .a({\u2_Display/n4543 ,\u2_Display/n4544 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c11 ),
    .fco(\u2_Display/lt143_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_14|u2_Display/lt143_13  (
    .a({\u2_Display/n4541 ,\u2_Display/n4542 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c13 ),
    .fco(\u2_Display/lt143_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_16|u2_Display/lt143_15  (
    .a({\u2_Display/n4539 ,\u2_Display/n4540 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c15 ),
    .fco(\u2_Display/lt143_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_18|u2_Display/lt143_17  (
    .a({\u2_Display/n4537 ,\u2_Display/n4538 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c17 ),
    .fco(\u2_Display/lt143_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_20|u2_Display/lt143_19  (
    .a({\u2_Display/n4535 ,\u2_Display/n4536 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c19 ),
    .fco(\u2_Display/lt143_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_22|u2_Display/lt143_21  (
    .a({\u2_Display/n4533 ,\u2_Display/n4534 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c21 ),
    .fco(\u2_Display/lt143_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_24|u2_Display/lt143_23  (
    .a({\u2_Display/n4531 ,\u2_Display/n4532 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c23 ),
    .fco(\u2_Display/lt143_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_26|u2_Display/lt143_25  (
    .a({\u2_Display/n4529 ,\u2_Display/n4530 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c25 ),
    .fco(\u2_Display/lt143_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_28|u2_Display/lt143_27  (
    .a({\u2_Display/n4527 ,\u2_Display/n4528 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c27 ),
    .fco(\u2_Display/lt143_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_2|u2_Display/lt143_1  (
    .a({\u2_Display/n4553 ,\u2_Display/n4554 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c1 ),
    .fco(\u2_Display/lt143_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_30|u2_Display/lt143_29  (
    .a({\u2_Display/n4525 ,\u2_Display/n4526 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c29 ),
    .fco(\u2_Display/lt143_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_4|u2_Display/lt143_3  (
    .a({\u2_Display/n4551 ,\u2_Display/n4552 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c3 ),
    .fco(\u2_Display/lt143_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_6|u2_Display/lt143_5  (
    .a({\u2_Display/n4549 ,\u2_Display/n4550 }),
    .b(2'b01),
    .fci(\u2_Display/lt143_c5 ),
    .fco(\u2_Display/lt143_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_8|u2_Display/lt143_7  (
    .a({\u2_Display/n4547 ,\u2_Display/n4548 }),
    .b(2'b10),
    .fci(\u2_Display/lt143_c7 ),
    .fco(\u2_Display/lt143_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_cout|u2_Display/lt143_31  (
    .a({1'b0,\u2_Display/n4524 }),
    .b(2'b10),
    .fci(\u2_Display/lt143_c31 ),
    .f({\u2_Display/n4556 ,open_n83764}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_0|u2_Display/lt154_cin  (
    .a({\u2_Display/counta [0],1'b0}),
    .b({1'b0,open_n83770}),
    .fco(\u2_Display/lt154_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_10|u2_Display/lt154_9  (
    .a(\u2_Display/counta [10:9]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c9 ),
    .fco(\u2_Display/lt154_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_12|u2_Display/lt154_11  (
    .a(\u2_Display/counta [12:11]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c11 ),
    .fco(\u2_Display/lt154_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_14|u2_Display/lt154_13  (
    .a(\u2_Display/counta [14:13]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c13 ),
    .fco(\u2_Display/lt154_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_16|u2_Display/lt154_15  (
    .a(\u2_Display/counta [16:15]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c15 ),
    .fco(\u2_Display/lt154_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_18|u2_Display/lt154_17  (
    .a(\u2_Display/counta [18:17]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c17 ),
    .fco(\u2_Display/lt154_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_20|u2_Display/lt154_19  (
    .a(\u2_Display/counta [20:19]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c19 ),
    .fco(\u2_Display/lt154_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_22|u2_Display/lt154_21  (
    .a(\u2_Display/counta [22:21]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c21 ),
    .fco(\u2_Display/lt154_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_24|u2_Display/lt154_23  (
    .a(\u2_Display/counta [24:23]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c23 ),
    .fco(\u2_Display/lt154_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_26|u2_Display/lt154_25  (
    .a(\u2_Display/counta [26:25]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c25 ),
    .fco(\u2_Display/lt154_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_28|u2_Display/lt154_27  (
    .a(\u2_Display/counta [28:27]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c27 ),
    .fco(\u2_Display/lt154_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_2|u2_Display/lt154_1  (
    .a(\u2_Display/counta [2:1]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c1 ),
    .fco(\u2_Display/lt154_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_30|u2_Display/lt154_29  (
    .a(\u2_Display/counta [30:29]),
    .b(2'b01),
    .fci(\u2_Display/lt154_c29 ),
    .fco(\u2_Display/lt154_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_4|u2_Display/lt154_3  (
    .a(\u2_Display/counta [4:3]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c3 ),
    .fco(\u2_Display/lt154_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_6|u2_Display/lt154_5  (
    .a(\u2_Display/counta [6:5]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c5 ),
    .fco(\u2_Display/lt154_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_8|u2_Display/lt154_7  (
    .a(\u2_Display/counta [8:7]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c7 ),
    .fco(\u2_Display/lt154_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_cout|u2_Display/lt154_31  (
    .a({1'b0,\u2_Display/counta [31]}),
    .b(2'b11),
    .fci(\u2_Display/lt154_c31 ),
    .f({\u2_Display/n4909 ,open_n84174}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_0|u2_Display/lt155_cin  (
    .a({\u2_Display/n6101 ,1'b0}),
    .b({1'b0,open_n84180}),
    .fco(\u2_Display/lt155_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_10|u2_Display/lt155_9  (
    .a({\u2_Display/n6091 ,\u2_Display/n6092 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c9 ),
    .fco(\u2_Display/lt155_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_12|u2_Display/lt155_11  (
    .a({\u2_Display/n6089 ,\u2_Display/n6090 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c11 ),
    .fco(\u2_Display/lt155_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_14|u2_Display/lt155_13  (
    .a({\u2_Display/n6087 ,\u2_Display/n6088 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c13 ),
    .fco(\u2_Display/lt155_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_16|u2_Display/lt155_15  (
    .a({\u2_Display/n6085 ,\u2_Display/n6086 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c15 ),
    .fco(\u2_Display/lt155_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_18|u2_Display/lt155_17  (
    .a({\u2_Display/n6083 ,\u2_Display/n6084 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c17 ),
    .fco(\u2_Display/lt155_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_20|u2_Display/lt155_19  (
    .a({\u2_Display/n6081 ,\u2_Display/n6082 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c19 ),
    .fco(\u2_Display/lt155_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_22|u2_Display/lt155_21  (
    .a({\u2_Display/n6079 ,\u2_Display/n6080 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c21 ),
    .fco(\u2_Display/lt155_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_24|u2_Display/lt155_23  (
    .a({\u2_Display/n6077 ,\u2_Display/n6078 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c23 ),
    .fco(\u2_Display/lt155_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_26|u2_Display/lt155_25  (
    .a({\u2_Display/n6075 ,\u2_Display/n6076 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c25 ),
    .fco(\u2_Display/lt155_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_28|u2_Display/lt155_27  (
    .a({\u2_Display/n6073 ,\u2_Display/n6074 }),
    .b(2'b10),
    .fci(\u2_Display/lt155_c27 ),
    .fco(\u2_Display/lt155_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_2|u2_Display/lt155_1  (
    .a({\u2_Display/n6099 ,\u2_Display/n6100 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c1 ),
    .fco(\u2_Display/lt155_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_30|u2_Display/lt155_29  (
    .a({\u2_Display/n6071 ,\u2_Display/n6072 }),
    .b(2'b10),
    .fci(\u2_Display/lt155_c29 ),
    .fco(\u2_Display/lt155_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_4|u2_Display/lt155_3  (
    .a({\u2_Display/n6097 ,\u2_Display/n6098 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c3 ),
    .fco(\u2_Display/lt155_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_6|u2_Display/lt155_5  (
    .a({\u2_Display/n6095 ,\u2_Display/n6096 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c5 ),
    .fco(\u2_Display/lt155_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_8|u2_Display/lt155_7  (
    .a({\u2_Display/n6093 ,\u2_Display/n6094 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c7 ),
    .fco(\u2_Display/lt155_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_cout|u2_Display/lt155_31  (
    .a({1'b0,\u2_Display/n6070 }),
    .b(2'b10),
    .fci(\u2_Display/lt155_c31 ),
    .f({\u2_Display/n4944 ,open_n84584}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_0|u2_Display/lt156_cin  (
    .a({\u2_Display/n6136 ,1'b0}),
    .b({1'b0,open_n84590}),
    .fco(\u2_Display/lt156_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_10|u2_Display/lt156_9  (
    .a({\u2_Display/n6126 ,\u2_Display/n6127 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c9 ),
    .fco(\u2_Display/lt156_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_12|u2_Display/lt156_11  (
    .a({\u2_Display/n6124 ,\u2_Display/n6125 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c11 ),
    .fco(\u2_Display/lt156_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_14|u2_Display/lt156_13  (
    .a({\u2_Display/n6122 ,\u2_Display/n6123 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c13 ),
    .fco(\u2_Display/lt156_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_16|u2_Display/lt156_15  (
    .a({\u2_Display/n6120 ,\u2_Display/n6121 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c15 ),
    .fco(\u2_Display/lt156_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_18|u2_Display/lt156_17  (
    .a({\u2_Display/n6118 ,\u2_Display/n6119 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c17 ),
    .fco(\u2_Display/lt156_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_20|u2_Display/lt156_19  (
    .a({\u2_Display/n6116 ,\u2_Display/n6117 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c19 ),
    .fco(\u2_Display/lt156_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_22|u2_Display/lt156_21  (
    .a({\u2_Display/n6114 ,\u2_Display/n6115 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c21 ),
    .fco(\u2_Display/lt156_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_24|u2_Display/lt156_23  (
    .a({\u2_Display/n6112 ,\u2_Display/n6113 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c23 ),
    .fco(\u2_Display/lt156_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_26|u2_Display/lt156_25  (
    .a({\u2_Display/n6110 ,\u2_Display/n6111 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c25 ),
    .fco(\u2_Display/lt156_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_28|u2_Display/lt156_27  (
    .a({\u2_Display/n6108 ,\u2_Display/n6109 }),
    .b(2'b01),
    .fci(\u2_Display/lt156_c27 ),
    .fco(\u2_Display/lt156_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_2|u2_Display/lt156_1  (
    .a({\u2_Display/n6134 ,\u2_Display/n6135 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c1 ),
    .fco(\u2_Display/lt156_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_30|u2_Display/lt156_29  (
    .a({\u2_Display/n6106 ,\u2_Display/n6107 }),
    .b(2'b01),
    .fci(\u2_Display/lt156_c29 ),
    .fco(\u2_Display/lt156_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_4|u2_Display/lt156_3  (
    .a({\u2_Display/n6132 ,\u2_Display/n6133 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c3 ),
    .fco(\u2_Display/lt156_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_6|u2_Display/lt156_5  (
    .a({\u2_Display/n6130 ,\u2_Display/n6131 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c5 ),
    .fco(\u2_Display/lt156_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_8|u2_Display/lt156_7  (
    .a({\u2_Display/n6128 ,\u2_Display/n6129 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c7 ),
    .fco(\u2_Display/lt156_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_cout|u2_Display/lt156_31  (
    .a({1'b0,\u2_Display/n6105 }),
    .b(2'b10),
    .fci(\u2_Display/lt156_c31 ),
    .f({\u2_Display/n4979 ,open_n84994}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_0|u2_Display/lt157_cin  (
    .a({\u2_Display/n6171 ,1'b0}),
    .b({1'b0,open_n85000}),
    .fco(\u2_Display/lt157_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_10|u2_Display/lt157_9  (
    .a({\u2_Display/n6161 ,\u2_Display/n6162 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c9 ),
    .fco(\u2_Display/lt157_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_12|u2_Display/lt157_11  (
    .a({\u2_Display/n6159 ,\u2_Display/n6160 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c11 ),
    .fco(\u2_Display/lt157_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_14|u2_Display/lt157_13  (
    .a({\u2_Display/n6157 ,\u2_Display/n6158 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c13 ),
    .fco(\u2_Display/lt157_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_16|u2_Display/lt157_15  (
    .a({\u2_Display/n6155 ,\u2_Display/n6156 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c15 ),
    .fco(\u2_Display/lt157_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_18|u2_Display/lt157_17  (
    .a({\u2_Display/n6153 ,\u2_Display/n6154 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c17 ),
    .fco(\u2_Display/lt157_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_20|u2_Display/lt157_19  (
    .a({\u2_Display/n6151 ,\u2_Display/n6152 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c19 ),
    .fco(\u2_Display/lt157_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_22|u2_Display/lt157_21  (
    .a({\u2_Display/n6149 ,\u2_Display/n6150 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c21 ),
    .fco(\u2_Display/lt157_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_24|u2_Display/lt157_23  (
    .a({\u2_Display/n6147 ,\u2_Display/n6148 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c23 ),
    .fco(\u2_Display/lt157_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_26|u2_Display/lt157_25  (
    .a({\u2_Display/n6145 ,\u2_Display/n6146 }),
    .b(2'b10),
    .fci(\u2_Display/lt157_c25 ),
    .fco(\u2_Display/lt157_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_28|u2_Display/lt157_27  (
    .a({\u2_Display/n6143 ,\u2_Display/n6144 }),
    .b(2'b10),
    .fci(\u2_Display/lt157_c27 ),
    .fco(\u2_Display/lt157_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_2|u2_Display/lt157_1  (
    .a({\u2_Display/n6169 ,\u2_Display/n6170 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c1 ),
    .fco(\u2_Display/lt157_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_30|u2_Display/lt157_29  (
    .a({\u2_Display/n6141 ,\u2_Display/n6142 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c29 ),
    .fco(\u2_Display/lt157_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_4|u2_Display/lt157_3  (
    .a({\u2_Display/n6167 ,\u2_Display/n6168 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c3 ),
    .fco(\u2_Display/lt157_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_6|u2_Display/lt157_5  (
    .a({\u2_Display/n6165 ,\u2_Display/n6166 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c5 ),
    .fco(\u2_Display/lt157_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_8|u2_Display/lt157_7  (
    .a({\u2_Display/n6163 ,\u2_Display/n6164 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c7 ),
    .fco(\u2_Display/lt157_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_cout|u2_Display/lt157_31  (
    .a({1'b0,\u2_Display/n6140 }),
    .b(2'b10),
    .fci(\u2_Display/lt157_c31 ),
    .f({\u2_Display/n5014 ,open_n85404}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_0|u2_Display/lt158_cin  (
    .a({\u2_Display/n6206 ,1'b0}),
    .b({1'b0,open_n85410}),
    .fco(\u2_Display/lt158_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_10|u2_Display/lt158_9  (
    .a({\u2_Display/n6196 ,\u2_Display/n6197 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c9 ),
    .fco(\u2_Display/lt158_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_12|u2_Display/lt158_11  (
    .a({\u2_Display/n6194 ,\u2_Display/n6195 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c11 ),
    .fco(\u2_Display/lt158_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_14|u2_Display/lt158_13  (
    .a({\u2_Display/n6192 ,\u2_Display/n6193 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c13 ),
    .fco(\u2_Display/lt158_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_16|u2_Display/lt158_15  (
    .a({\u2_Display/n6190 ,\u2_Display/n6191 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c15 ),
    .fco(\u2_Display/lt158_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_18|u2_Display/lt158_17  (
    .a({\u2_Display/n6188 ,\u2_Display/n6189 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c17 ),
    .fco(\u2_Display/lt158_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_20|u2_Display/lt158_19  (
    .a({\u2_Display/n6186 ,\u2_Display/n6187 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c19 ),
    .fco(\u2_Display/lt158_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_22|u2_Display/lt158_21  (
    .a({\u2_Display/n6184 ,\u2_Display/n6185 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c21 ),
    .fco(\u2_Display/lt158_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_24|u2_Display/lt158_23  (
    .a({\u2_Display/n6182 ,\u2_Display/n6183 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c23 ),
    .fco(\u2_Display/lt158_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_26|u2_Display/lt158_25  (
    .a({\u2_Display/n6180 ,\u2_Display/n6181 }),
    .b(2'b01),
    .fci(\u2_Display/lt158_c25 ),
    .fco(\u2_Display/lt158_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_28|u2_Display/lt158_27  (
    .a({\u2_Display/n6178 ,\u2_Display/n6179 }),
    .b(2'b01),
    .fci(\u2_Display/lt158_c27 ),
    .fco(\u2_Display/lt158_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_2|u2_Display/lt158_1  (
    .a({\u2_Display/n6204 ,\u2_Display/n6205 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c1 ),
    .fco(\u2_Display/lt158_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_30|u2_Display/lt158_29  (
    .a({\u2_Display/n6176 ,\u2_Display/n6177 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c29 ),
    .fco(\u2_Display/lt158_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_4|u2_Display/lt158_3  (
    .a({\u2_Display/n6202 ,\u2_Display/n6203 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c3 ),
    .fco(\u2_Display/lt158_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_6|u2_Display/lt158_5  (
    .a({\u2_Display/n6200 ,\u2_Display/n6201 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c5 ),
    .fco(\u2_Display/lt158_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_8|u2_Display/lt158_7  (
    .a({\u2_Display/n6198 ,\u2_Display/n6199 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c7 ),
    .fco(\u2_Display/lt158_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_cout|u2_Display/lt158_31  (
    .a({1'b0,\u2_Display/n6175 }),
    .b(2'b10),
    .fci(\u2_Display/lt158_c31 ),
    .f({\u2_Display/n5049 ,open_n85814}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_0|u2_Display/lt159_cin  (
    .a({\u2_Display/n6241 ,1'b0}),
    .b({1'b0,open_n85820}),
    .fco(\u2_Display/lt159_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_10|u2_Display/lt159_9  (
    .a({\u2_Display/n6231 ,\u2_Display/n6232 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c9 ),
    .fco(\u2_Display/lt159_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_12|u2_Display/lt159_11  (
    .a({\u2_Display/n6229 ,\u2_Display/n6230 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c11 ),
    .fco(\u2_Display/lt159_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_14|u2_Display/lt159_13  (
    .a({\u2_Display/n6227 ,\u2_Display/n6228 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c13 ),
    .fco(\u2_Display/lt159_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_16|u2_Display/lt159_15  (
    .a({\u2_Display/n6225 ,\u2_Display/n6226 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c15 ),
    .fco(\u2_Display/lt159_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_18|u2_Display/lt159_17  (
    .a({\u2_Display/n6223 ,\u2_Display/n6224 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c17 ),
    .fco(\u2_Display/lt159_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_20|u2_Display/lt159_19  (
    .a({\u2_Display/n6221 ,\u2_Display/n6222 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c19 ),
    .fco(\u2_Display/lt159_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_22|u2_Display/lt159_21  (
    .a({\u2_Display/n6219 ,\u2_Display/n6220 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c21 ),
    .fco(\u2_Display/lt159_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_24|u2_Display/lt159_23  (
    .a({\u2_Display/n6217 ,\u2_Display/n6218 }),
    .b(2'b10),
    .fci(\u2_Display/lt159_c23 ),
    .fco(\u2_Display/lt159_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_26|u2_Display/lt159_25  (
    .a({\u2_Display/n6215 ,\u2_Display/n6216 }),
    .b(2'b10),
    .fci(\u2_Display/lt159_c25 ),
    .fco(\u2_Display/lt159_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_28|u2_Display/lt159_27  (
    .a({\u2_Display/n6213 ,\u2_Display/n6214 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c27 ),
    .fco(\u2_Display/lt159_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_2|u2_Display/lt159_1  (
    .a({\u2_Display/n6239 ,\u2_Display/n6240 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c1 ),
    .fco(\u2_Display/lt159_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_30|u2_Display/lt159_29  (
    .a({\u2_Display/n6211 ,\u2_Display/n6212 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c29 ),
    .fco(\u2_Display/lt159_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_4|u2_Display/lt159_3  (
    .a({\u2_Display/n6237 ,\u2_Display/n6238 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c3 ),
    .fco(\u2_Display/lt159_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_6|u2_Display/lt159_5  (
    .a({\u2_Display/n6235 ,\u2_Display/n6236 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c5 ),
    .fco(\u2_Display/lt159_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_8|u2_Display/lt159_7  (
    .a({\u2_Display/n6233 ,\u2_Display/n6234 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c7 ),
    .fco(\u2_Display/lt159_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_cout|u2_Display/lt159_31  (
    .a({1'b0,\u2_Display/n6210 }),
    .b(2'b10),
    .fci(\u2_Display/lt159_c31 ),
    .f({\u2_Display/n5084 ,open_n86224}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_0|u2_Display/lt160_cin  (
    .a({\u2_Display/n6276 ,1'b0}),
    .b({1'b0,open_n86230}),
    .fco(\u2_Display/lt160_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_10|u2_Display/lt160_9  (
    .a({\u2_Display/n6266 ,\u2_Display/n6267 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c9 ),
    .fco(\u2_Display/lt160_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_12|u2_Display/lt160_11  (
    .a({\u2_Display/n6264 ,\u2_Display/n6265 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c11 ),
    .fco(\u2_Display/lt160_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_14|u2_Display/lt160_13  (
    .a({\u2_Display/n6262 ,\u2_Display/n6263 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c13 ),
    .fco(\u2_Display/lt160_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_16|u2_Display/lt160_15  (
    .a({\u2_Display/n6260 ,\u2_Display/n6261 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c15 ),
    .fco(\u2_Display/lt160_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_18|u2_Display/lt160_17  (
    .a({\u2_Display/n6258 ,\u2_Display/n6259 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c17 ),
    .fco(\u2_Display/lt160_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_20|u2_Display/lt160_19  (
    .a({\u2_Display/n6256 ,\u2_Display/n6257 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c19 ),
    .fco(\u2_Display/lt160_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_22|u2_Display/lt160_21  (
    .a({\u2_Display/n6254 ,\u2_Display/n6255 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c21 ),
    .fco(\u2_Display/lt160_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_24|u2_Display/lt160_23  (
    .a({\u2_Display/n6252 ,\u2_Display/n6253 }),
    .b(2'b01),
    .fci(\u2_Display/lt160_c23 ),
    .fco(\u2_Display/lt160_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_26|u2_Display/lt160_25  (
    .a({\u2_Display/n6250 ,\u2_Display/n6251 }),
    .b(2'b01),
    .fci(\u2_Display/lt160_c25 ),
    .fco(\u2_Display/lt160_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_28|u2_Display/lt160_27  (
    .a({\u2_Display/n6248 ,\u2_Display/n6249 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c27 ),
    .fco(\u2_Display/lt160_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_2|u2_Display/lt160_1  (
    .a({\u2_Display/n6274 ,\u2_Display/n6275 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c1 ),
    .fco(\u2_Display/lt160_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_30|u2_Display/lt160_29  (
    .a({\u2_Display/n6246 ,\u2_Display/n6247 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c29 ),
    .fco(\u2_Display/lt160_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_4|u2_Display/lt160_3  (
    .a({\u2_Display/n6272 ,\u2_Display/n6273 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c3 ),
    .fco(\u2_Display/lt160_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_6|u2_Display/lt160_5  (
    .a({\u2_Display/n6270 ,\u2_Display/n6271 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c5 ),
    .fco(\u2_Display/lt160_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_8|u2_Display/lt160_7  (
    .a({\u2_Display/n6268 ,\u2_Display/n6269 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c7 ),
    .fco(\u2_Display/lt160_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_cout|u2_Display/lt160_31  (
    .a({1'b0,\u2_Display/n6245 }),
    .b(2'b10),
    .fci(\u2_Display/lt160_c31 ),
    .f({\u2_Display/n5119 ,open_n86634}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_0|u2_Display/lt161_cin  (
    .a({\u2_Display/n6311 ,1'b0}),
    .b({1'b0,open_n86640}),
    .fco(\u2_Display/lt161_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_10|u2_Display/lt161_9  (
    .a({\u2_Display/n6301 ,\u2_Display/n6302 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c9 ),
    .fco(\u2_Display/lt161_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_12|u2_Display/lt161_11  (
    .a({\u2_Display/n6299 ,\u2_Display/n6300 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c11 ),
    .fco(\u2_Display/lt161_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_14|u2_Display/lt161_13  (
    .a({\u2_Display/n6297 ,\u2_Display/n6298 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c13 ),
    .fco(\u2_Display/lt161_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_16|u2_Display/lt161_15  (
    .a({\u2_Display/n6295 ,\u2_Display/n6296 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c15 ),
    .fco(\u2_Display/lt161_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_18|u2_Display/lt161_17  (
    .a({\u2_Display/n6293 ,\u2_Display/n6294 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c17 ),
    .fco(\u2_Display/lt161_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_20|u2_Display/lt161_19  (
    .a({\u2_Display/n6291 ,\u2_Display/n6292 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c19 ),
    .fco(\u2_Display/lt161_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_22|u2_Display/lt161_21  (
    .a({\u2_Display/n6289 ,\u2_Display/n6290 }),
    .b(2'b10),
    .fci(\u2_Display/lt161_c21 ),
    .fco(\u2_Display/lt161_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_24|u2_Display/lt161_23  (
    .a({\u2_Display/n6287 ,\u2_Display/n6288 }),
    .b(2'b10),
    .fci(\u2_Display/lt161_c23 ),
    .fco(\u2_Display/lt161_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_26|u2_Display/lt161_25  (
    .a({\u2_Display/n6285 ,\u2_Display/n6286 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c25 ),
    .fco(\u2_Display/lt161_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_28|u2_Display/lt161_27  (
    .a({\u2_Display/n6283 ,\u2_Display/n6284 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c27 ),
    .fco(\u2_Display/lt161_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_2|u2_Display/lt161_1  (
    .a({\u2_Display/n6309 ,\u2_Display/n6310 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c1 ),
    .fco(\u2_Display/lt161_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_30|u2_Display/lt161_29  (
    .a({\u2_Display/n6281 ,\u2_Display/n6282 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c29 ),
    .fco(\u2_Display/lt161_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_4|u2_Display/lt161_3  (
    .a({\u2_Display/n6307 ,\u2_Display/n6308 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c3 ),
    .fco(\u2_Display/lt161_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_6|u2_Display/lt161_5  (
    .a({\u2_Display/n6305 ,\u2_Display/n6306 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c5 ),
    .fco(\u2_Display/lt161_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_8|u2_Display/lt161_7  (
    .a({\u2_Display/n6303 ,\u2_Display/n6304 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c7 ),
    .fco(\u2_Display/lt161_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_cout|u2_Display/lt161_31  (
    .a({1'b0,\u2_Display/n6280 }),
    .b(2'b10),
    .fci(\u2_Display/lt161_c31 ),
    .f({\u2_Display/n5154 ,open_n87044}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_0|u2_Display/lt162_cin  (
    .a({\u2_Display/n6346 ,1'b0}),
    .b({1'b0,open_n87050}),
    .fco(\u2_Display/lt162_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_10|u2_Display/lt162_9  (
    .a({\u2_Display/n6336 ,\u2_Display/n6337 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c9 ),
    .fco(\u2_Display/lt162_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_12|u2_Display/lt162_11  (
    .a({\u2_Display/n6334 ,\u2_Display/n6335 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c11 ),
    .fco(\u2_Display/lt162_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_14|u2_Display/lt162_13  (
    .a({\u2_Display/n6332 ,\u2_Display/n6333 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c13 ),
    .fco(\u2_Display/lt162_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_16|u2_Display/lt162_15  (
    .a({\u2_Display/n6330 ,\u2_Display/n6331 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c15 ),
    .fco(\u2_Display/lt162_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_18|u2_Display/lt162_17  (
    .a({\u2_Display/n6328 ,\u2_Display/n6329 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c17 ),
    .fco(\u2_Display/lt162_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_20|u2_Display/lt162_19  (
    .a({\u2_Display/n6326 ,\u2_Display/n6327 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c19 ),
    .fco(\u2_Display/lt162_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_22|u2_Display/lt162_21  (
    .a({\u2_Display/n6324 ,\u2_Display/n6325 }),
    .b(2'b01),
    .fci(\u2_Display/lt162_c21 ),
    .fco(\u2_Display/lt162_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_24|u2_Display/lt162_23  (
    .a({\u2_Display/n6322 ,\u2_Display/n6323 }),
    .b(2'b01),
    .fci(\u2_Display/lt162_c23 ),
    .fco(\u2_Display/lt162_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_26|u2_Display/lt162_25  (
    .a({\u2_Display/n6320 ,\u2_Display/n6321 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c25 ),
    .fco(\u2_Display/lt162_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_28|u2_Display/lt162_27  (
    .a({\u2_Display/n6318 ,\u2_Display/n6319 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c27 ),
    .fco(\u2_Display/lt162_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_2|u2_Display/lt162_1  (
    .a({\u2_Display/n6344 ,\u2_Display/n6345 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c1 ),
    .fco(\u2_Display/lt162_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_30|u2_Display/lt162_29  (
    .a({\u2_Display/n6316 ,\u2_Display/n6317 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c29 ),
    .fco(\u2_Display/lt162_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_4|u2_Display/lt162_3  (
    .a({\u2_Display/n6342 ,\u2_Display/n6343 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c3 ),
    .fco(\u2_Display/lt162_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_6|u2_Display/lt162_5  (
    .a({\u2_Display/n6340 ,\u2_Display/n6341 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c5 ),
    .fco(\u2_Display/lt162_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_8|u2_Display/lt162_7  (
    .a({\u2_Display/n6338 ,\u2_Display/n6339 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c7 ),
    .fco(\u2_Display/lt162_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_cout|u2_Display/lt162_31  (
    .a({1'b0,\u2_Display/n6315 }),
    .b(2'b10),
    .fci(\u2_Display/lt162_c31 ),
    .f({\u2_Display/n5189 ,open_n87454}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_0|u2_Display/lt163_cin  (
    .a({\u2_Display/n5223 ,1'b0}),
    .b({1'b0,open_n87460}),
    .fco(\u2_Display/lt163_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_10|u2_Display/lt163_9  (
    .a({\u2_Display/n5213 ,\u2_Display/n5214 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c9 ),
    .fco(\u2_Display/lt163_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_12|u2_Display/lt163_11  (
    .a({\u2_Display/n5211 ,\u2_Display/n5212 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c11 ),
    .fco(\u2_Display/lt163_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_14|u2_Display/lt163_13  (
    .a({\u2_Display/n5209 ,\u2_Display/n5210 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c13 ),
    .fco(\u2_Display/lt163_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_16|u2_Display/lt163_15  (
    .a({\u2_Display/n5207 ,\u2_Display/n5208 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c15 ),
    .fco(\u2_Display/lt163_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_18|u2_Display/lt163_17  (
    .a({\u2_Display/n5205 ,\u2_Display/n5206 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c17 ),
    .fco(\u2_Display/lt163_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_20|u2_Display/lt163_19  (
    .a({\u2_Display/n5203 ,\u2_Display/n5204 }),
    .b(2'b10),
    .fci(\u2_Display/lt163_c19 ),
    .fco(\u2_Display/lt163_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_22|u2_Display/lt163_21  (
    .a({\u2_Display/n5201 ,\u2_Display/n5202 }),
    .b(2'b10),
    .fci(\u2_Display/lt163_c21 ),
    .fco(\u2_Display/lt163_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_24|u2_Display/lt163_23  (
    .a({\u2_Display/n5199 ,\u2_Display/n5200 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c23 ),
    .fco(\u2_Display/lt163_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_26|u2_Display/lt163_25  (
    .a({\u2_Display/n5197 ,\u2_Display/n5198 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c25 ),
    .fco(\u2_Display/lt163_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_28|u2_Display/lt163_27  (
    .a({\u2_Display/n6353 ,\u2_Display/n5196 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c27 ),
    .fco(\u2_Display/lt163_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_2|u2_Display/lt163_1  (
    .a({\u2_Display/n5221 ,\u2_Display/n5222 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c1 ),
    .fco(\u2_Display/lt163_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_30|u2_Display/lt163_29  (
    .a({\u2_Display/n6351 ,\u2_Display/n6352 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c29 ),
    .fco(\u2_Display/lt163_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_4|u2_Display/lt163_3  (
    .a({\u2_Display/n5219 ,\u2_Display/n5220 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c3 ),
    .fco(\u2_Display/lt163_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_6|u2_Display/lt163_5  (
    .a({\u2_Display/n5217 ,\u2_Display/n5218 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c5 ),
    .fco(\u2_Display/lt163_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_8|u2_Display/lt163_7  (
    .a({\u2_Display/n5215 ,\u2_Display/n5216 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c7 ),
    .fco(\u2_Display/lt163_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_cout|u2_Display/lt163_31  (
    .a({1'b0,\u2_Display/n6350 }),
    .b(2'b10),
    .fci(\u2_Display/lt163_c31 ),
    .f({\u2_Display/n5224 ,open_n87864}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_0|u2_Display/lt164_cin  (
    .a({\u2_Display/n5258 ,1'b0}),
    .b({1'b0,open_n87870}),
    .fco(\u2_Display/lt164_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_10|u2_Display/lt164_9  (
    .a({\u2_Display/n5248 ,\u2_Display/n5249 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c9 ),
    .fco(\u2_Display/lt164_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_12|u2_Display/lt164_11  (
    .a({\u2_Display/n5246 ,\u2_Display/n5247 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c11 ),
    .fco(\u2_Display/lt164_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_14|u2_Display/lt164_13  (
    .a({\u2_Display/n5244 ,\u2_Display/n5245 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c13 ),
    .fco(\u2_Display/lt164_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_16|u2_Display/lt164_15  (
    .a({\u2_Display/n5242 ,\u2_Display/n5243 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c15 ),
    .fco(\u2_Display/lt164_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_18|u2_Display/lt164_17  (
    .a({\u2_Display/n5240 ,\u2_Display/n5241 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c17 ),
    .fco(\u2_Display/lt164_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_20|u2_Display/lt164_19  (
    .a({\u2_Display/n5238 ,\u2_Display/n5239 }),
    .b(2'b01),
    .fci(\u2_Display/lt164_c19 ),
    .fco(\u2_Display/lt164_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_22|u2_Display/lt164_21  (
    .a({\u2_Display/n5236 ,\u2_Display/n5237 }),
    .b(2'b01),
    .fci(\u2_Display/lt164_c21 ),
    .fco(\u2_Display/lt164_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_24|u2_Display/lt164_23  (
    .a({\u2_Display/n5234 ,\u2_Display/n5235 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c23 ),
    .fco(\u2_Display/lt164_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_26|u2_Display/lt164_25  (
    .a({\u2_Display/n5232 ,\u2_Display/n5233 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c25 ),
    .fco(\u2_Display/lt164_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_28|u2_Display/lt164_27  (
    .a({\u2_Display/n5230 ,\u2_Display/n5231 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c27 ),
    .fco(\u2_Display/lt164_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_2|u2_Display/lt164_1  (
    .a({\u2_Display/n5256 ,\u2_Display/n5257 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c1 ),
    .fco(\u2_Display/lt164_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_30|u2_Display/lt164_29  (
    .a({\u2_Display/n5228 ,\u2_Display/n5229 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c29 ),
    .fco(\u2_Display/lt164_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_4|u2_Display/lt164_3  (
    .a({\u2_Display/n5254 ,\u2_Display/n5255 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c3 ),
    .fco(\u2_Display/lt164_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_6|u2_Display/lt164_5  (
    .a({\u2_Display/n5252 ,\u2_Display/n5253 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c5 ),
    .fco(\u2_Display/lt164_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_8|u2_Display/lt164_7  (
    .a({\u2_Display/n5250 ,\u2_Display/n5251 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c7 ),
    .fco(\u2_Display/lt164_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_cout|u2_Display/lt164_31  (
    .a({1'b0,\u2_Display/n5227 }),
    .b(2'b10),
    .fci(\u2_Display/lt164_c31 ),
    .f({\u2_Display/n5259 ,open_n88274}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_0|u2_Display/lt165_cin  (
    .a({\u2_Display/n5293 ,1'b0}),
    .b({1'b0,open_n88280}),
    .fco(\u2_Display/lt165_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_10|u2_Display/lt165_9  (
    .a({\u2_Display/n5283 ,\u2_Display/n5284 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c9 ),
    .fco(\u2_Display/lt165_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_12|u2_Display/lt165_11  (
    .a({\u2_Display/n5281 ,\u2_Display/n5282 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c11 ),
    .fco(\u2_Display/lt165_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_14|u2_Display/lt165_13  (
    .a({\u2_Display/n5279 ,\u2_Display/n5280 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c13 ),
    .fco(\u2_Display/lt165_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_16|u2_Display/lt165_15  (
    .a({\u2_Display/n5277 ,\u2_Display/n5278 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c15 ),
    .fco(\u2_Display/lt165_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_18|u2_Display/lt165_17  (
    .a({\u2_Display/n5275 ,\u2_Display/n5276 }),
    .b(2'b10),
    .fci(\u2_Display/lt165_c17 ),
    .fco(\u2_Display/lt165_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_20|u2_Display/lt165_19  (
    .a({\u2_Display/n5273 ,\u2_Display/n5274 }),
    .b(2'b10),
    .fci(\u2_Display/lt165_c19 ),
    .fco(\u2_Display/lt165_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_22|u2_Display/lt165_21  (
    .a({\u2_Display/n5271 ,\u2_Display/n5272 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c21 ),
    .fco(\u2_Display/lt165_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_24|u2_Display/lt165_23  (
    .a({\u2_Display/n5269 ,\u2_Display/n5270 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c23 ),
    .fco(\u2_Display/lt165_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_26|u2_Display/lt165_25  (
    .a({\u2_Display/n5267 ,\u2_Display/n5268 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c25 ),
    .fco(\u2_Display/lt165_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_28|u2_Display/lt165_27  (
    .a({\u2_Display/n5265 ,\u2_Display/n5266 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c27 ),
    .fco(\u2_Display/lt165_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_2|u2_Display/lt165_1  (
    .a({\u2_Display/n5291 ,\u2_Display/n5292 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c1 ),
    .fco(\u2_Display/lt165_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_30|u2_Display/lt165_29  (
    .a({\u2_Display/n5263 ,\u2_Display/n5264 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c29 ),
    .fco(\u2_Display/lt165_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_4|u2_Display/lt165_3  (
    .a({\u2_Display/n5289 ,\u2_Display/n5290 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c3 ),
    .fco(\u2_Display/lt165_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_6|u2_Display/lt165_5  (
    .a({\u2_Display/n5287 ,\u2_Display/n5288 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c5 ),
    .fco(\u2_Display/lt165_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_8|u2_Display/lt165_7  (
    .a({\u2_Display/n5285 ,\u2_Display/n5286 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c7 ),
    .fco(\u2_Display/lt165_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_cout|u2_Display/lt165_31  (
    .a({1'b0,\u2_Display/n5262 }),
    .b(2'b10),
    .fci(\u2_Display/lt165_c31 ),
    .f({\u2_Display/n5294 ,open_n88684}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_0|u2_Display/lt166_cin  (
    .a({\u2_Display/n5328 ,1'b0}),
    .b({1'b0,open_n88690}),
    .fco(\u2_Display/lt166_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_10|u2_Display/lt166_9  (
    .a({\u2_Display/n5318 ,\u2_Display/n5319 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c9 ),
    .fco(\u2_Display/lt166_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_12|u2_Display/lt166_11  (
    .a({\u2_Display/n5316 ,\u2_Display/n5317 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c11 ),
    .fco(\u2_Display/lt166_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_14|u2_Display/lt166_13  (
    .a({\u2_Display/n5314 ,\u2_Display/n5315 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c13 ),
    .fco(\u2_Display/lt166_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_16|u2_Display/lt166_15  (
    .a({\u2_Display/n5312 ,\u2_Display/n5313 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c15 ),
    .fco(\u2_Display/lt166_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_18|u2_Display/lt166_17  (
    .a({\u2_Display/n5310 ,\u2_Display/n5311 }),
    .b(2'b01),
    .fci(\u2_Display/lt166_c17 ),
    .fco(\u2_Display/lt166_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_20|u2_Display/lt166_19  (
    .a({\u2_Display/n5308 ,\u2_Display/n5309 }),
    .b(2'b01),
    .fci(\u2_Display/lt166_c19 ),
    .fco(\u2_Display/lt166_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_22|u2_Display/lt166_21  (
    .a({\u2_Display/n5306 ,\u2_Display/n5307 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c21 ),
    .fco(\u2_Display/lt166_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_24|u2_Display/lt166_23  (
    .a({\u2_Display/n5304 ,\u2_Display/n5305 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c23 ),
    .fco(\u2_Display/lt166_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_26|u2_Display/lt166_25  (
    .a({\u2_Display/n5302 ,\u2_Display/n5303 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c25 ),
    .fco(\u2_Display/lt166_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_28|u2_Display/lt166_27  (
    .a({\u2_Display/n5300 ,\u2_Display/n5301 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c27 ),
    .fco(\u2_Display/lt166_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_2|u2_Display/lt166_1  (
    .a({\u2_Display/n5326 ,\u2_Display/n5327 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c1 ),
    .fco(\u2_Display/lt166_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_30|u2_Display/lt166_29  (
    .a({\u2_Display/n5298 ,\u2_Display/n5299 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c29 ),
    .fco(\u2_Display/lt166_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_4|u2_Display/lt166_3  (
    .a({\u2_Display/n5324 ,\u2_Display/n5325 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c3 ),
    .fco(\u2_Display/lt166_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_6|u2_Display/lt166_5  (
    .a({\u2_Display/n5322 ,\u2_Display/n5323 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c5 ),
    .fco(\u2_Display/lt166_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_8|u2_Display/lt166_7  (
    .a({\u2_Display/n5320 ,\u2_Display/n5321 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c7 ),
    .fco(\u2_Display/lt166_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_cout|u2_Display/lt166_31  (
    .a({1'b0,\u2_Display/n5297 }),
    .b(2'b10),
    .fci(\u2_Display/lt166_c31 ),
    .f({\u2_Display/n5329 ,open_n89094}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_0|u2_Display/lt167_cin  (
    .a({\u2_Display/n5363 ,1'b0}),
    .b({1'b0,open_n89100}),
    .fco(\u2_Display/lt167_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_10|u2_Display/lt167_9  (
    .a({\u2_Display/n5353 ,\u2_Display/n5354 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c9 ),
    .fco(\u2_Display/lt167_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_12|u2_Display/lt167_11  (
    .a({\u2_Display/n5351 ,\u2_Display/n5352 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c11 ),
    .fco(\u2_Display/lt167_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_14|u2_Display/lt167_13  (
    .a({\u2_Display/n5349 ,\u2_Display/n5350 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c13 ),
    .fco(\u2_Display/lt167_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_16|u2_Display/lt167_15  (
    .a({\u2_Display/n5347 ,\u2_Display/n5348 }),
    .b(2'b10),
    .fci(\u2_Display/lt167_c15 ),
    .fco(\u2_Display/lt167_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_18|u2_Display/lt167_17  (
    .a({\u2_Display/n5345 ,\u2_Display/n5346 }),
    .b(2'b10),
    .fci(\u2_Display/lt167_c17 ),
    .fco(\u2_Display/lt167_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_20|u2_Display/lt167_19  (
    .a({\u2_Display/n5343 ,\u2_Display/n5344 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c19 ),
    .fco(\u2_Display/lt167_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_22|u2_Display/lt167_21  (
    .a({\u2_Display/n5341 ,\u2_Display/n5342 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c21 ),
    .fco(\u2_Display/lt167_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_24|u2_Display/lt167_23  (
    .a({\u2_Display/n5339 ,\u2_Display/n5340 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c23 ),
    .fco(\u2_Display/lt167_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_26|u2_Display/lt167_25  (
    .a({\u2_Display/n5337 ,\u2_Display/n5338 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c25 ),
    .fco(\u2_Display/lt167_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_28|u2_Display/lt167_27  (
    .a({\u2_Display/n5335 ,\u2_Display/n5336 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c27 ),
    .fco(\u2_Display/lt167_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_2|u2_Display/lt167_1  (
    .a({\u2_Display/n5361 ,\u2_Display/n5362 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c1 ),
    .fco(\u2_Display/lt167_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_30|u2_Display/lt167_29  (
    .a({\u2_Display/n5333 ,\u2_Display/n5334 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c29 ),
    .fco(\u2_Display/lt167_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_4|u2_Display/lt167_3  (
    .a({\u2_Display/n5359 ,\u2_Display/n5360 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c3 ),
    .fco(\u2_Display/lt167_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_6|u2_Display/lt167_5  (
    .a({\u2_Display/n5357 ,\u2_Display/n5358 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c5 ),
    .fco(\u2_Display/lt167_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_8|u2_Display/lt167_7  (
    .a({\u2_Display/n5355 ,\u2_Display/n5356 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c7 ),
    .fco(\u2_Display/lt167_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_cout|u2_Display/lt167_31  (
    .a({1'b0,\u2_Display/n5332 }),
    .b(2'b10),
    .fci(\u2_Display/lt167_c31 ),
    .f({\u2_Display/n5364 ,open_n89504}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_0|u2_Display/lt168_cin  (
    .a({\u2_Display/n5398 ,1'b0}),
    .b({1'b0,open_n89510}),
    .fco(\u2_Display/lt168_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_10|u2_Display/lt168_9  (
    .a({\u2_Display/n5388 ,\u2_Display/n5389 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c9 ),
    .fco(\u2_Display/lt168_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_12|u2_Display/lt168_11  (
    .a({\u2_Display/n5386 ,\u2_Display/n5387 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c11 ),
    .fco(\u2_Display/lt168_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_14|u2_Display/lt168_13  (
    .a({\u2_Display/n5384 ,\u2_Display/n5385 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c13 ),
    .fco(\u2_Display/lt168_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_16|u2_Display/lt168_15  (
    .a({\u2_Display/n5382 ,\u2_Display/n5383 }),
    .b(2'b01),
    .fci(\u2_Display/lt168_c15 ),
    .fco(\u2_Display/lt168_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_18|u2_Display/lt168_17  (
    .a({\u2_Display/n5380 ,\u2_Display/n5381 }),
    .b(2'b01),
    .fci(\u2_Display/lt168_c17 ),
    .fco(\u2_Display/lt168_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_20|u2_Display/lt168_19  (
    .a({\u2_Display/n5378 ,\u2_Display/n5379 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c19 ),
    .fco(\u2_Display/lt168_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_22|u2_Display/lt168_21  (
    .a({\u2_Display/n5376 ,\u2_Display/n5377 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c21 ),
    .fco(\u2_Display/lt168_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_24|u2_Display/lt168_23  (
    .a({\u2_Display/n5374 ,\u2_Display/n5375 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c23 ),
    .fco(\u2_Display/lt168_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_26|u2_Display/lt168_25  (
    .a({\u2_Display/n5372 ,\u2_Display/n5373 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c25 ),
    .fco(\u2_Display/lt168_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_28|u2_Display/lt168_27  (
    .a({\u2_Display/n5370 ,\u2_Display/n5371 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c27 ),
    .fco(\u2_Display/lt168_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_2|u2_Display/lt168_1  (
    .a({\u2_Display/n5396 ,\u2_Display/n5397 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c1 ),
    .fco(\u2_Display/lt168_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_30|u2_Display/lt168_29  (
    .a({\u2_Display/n5368 ,\u2_Display/n5369 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c29 ),
    .fco(\u2_Display/lt168_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_4|u2_Display/lt168_3  (
    .a({\u2_Display/n5394 ,\u2_Display/n5395 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c3 ),
    .fco(\u2_Display/lt168_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_6|u2_Display/lt168_5  (
    .a({\u2_Display/n5392 ,\u2_Display/n5393 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c5 ),
    .fco(\u2_Display/lt168_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_8|u2_Display/lt168_7  (
    .a({\u2_Display/n5390 ,\u2_Display/n5391 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c7 ),
    .fco(\u2_Display/lt168_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_cout|u2_Display/lt168_31  (
    .a({1'b0,\u2_Display/n5367 }),
    .b(2'b10),
    .fci(\u2_Display/lt168_c31 ),
    .f({\u2_Display/n5399 ,open_n89914}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_0|u2_Display/lt169_cin  (
    .a({\u2_Display/n5433 ,1'b0}),
    .b({1'b0,open_n89920}),
    .fco(\u2_Display/lt169_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_10|u2_Display/lt169_9  (
    .a({\u2_Display/n5423 ,\u2_Display/n5424 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c9 ),
    .fco(\u2_Display/lt169_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_12|u2_Display/lt169_11  (
    .a({\u2_Display/n5421 ,\u2_Display/n5422 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c11 ),
    .fco(\u2_Display/lt169_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_14|u2_Display/lt169_13  (
    .a({\u2_Display/n5419 ,\u2_Display/n5420 }),
    .b(2'b10),
    .fci(\u2_Display/lt169_c13 ),
    .fco(\u2_Display/lt169_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_16|u2_Display/lt169_15  (
    .a({\u2_Display/n5417 ,\u2_Display/n5418 }),
    .b(2'b10),
    .fci(\u2_Display/lt169_c15 ),
    .fco(\u2_Display/lt169_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_18|u2_Display/lt169_17  (
    .a({\u2_Display/n5415 ,\u2_Display/n5416 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c17 ),
    .fco(\u2_Display/lt169_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_20|u2_Display/lt169_19  (
    .a({\u2_Display/n5413 ,\u2_Display/n5414 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c19 ),
    .fco(\u2_Display/lt169_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_22|u2_Display/lt169_21  (
    .a({\u2_Display/n5411 ,\u2_Display/n5412 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c21 ),
    .fco(\u2_Display/lt169_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_24|u2_Display/lt169_23  (
    .a({\u2_Display/n5409 ,\u2_Display/n5410 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c23 ),
    .fco(\u2_Display/lt169_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_26|u2_Display/lt169_25  (
    .a({\u2_Display/n5407 ,\u2_Display/n5408 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c25 ),
    .fco(\u2_Display/lt169_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_28|u2_Display/lt169_27  (
    .a({\u2_Display/n5405 ,\u2_Display/n5406 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c27 ),
    .fco(\u2_Display/lt169_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_2|u2_Display/lt169_1  (
    .a({\u2_Display/n5431 ,\u2_Display/n5432 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c1 ),
    .fco(\u2_Display/lt169_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_30|u2_Display/lt169_29  (
    .a({\u2_Display/n5403 ,\u2_Display/n5404 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c29 ),
    .fco(\u2_Display/lt169_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_4|u2_Display/lt169_3  (
    .a({\u2_Display/n5429 ,\u2_Display/n5430 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c3 ),
    .fco(\u2_Display/lt169_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_6|u2_Display/lt169_5  (
    .a({\u2_Display/n5427 ,\u2_Display/n5428 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c5 ),
    .fco(\u2_Display/lt169_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_8|u2_Display/lt169_7  (
    .a({\u2_Display/n5425 ,\u2_Display/n5426 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c7 ),
    .fco(\u2_Display/lt169_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_cout|u2_Display/lt169_31  (
    .a({1'b0,\u2_Display/n5402 }),
    .b(2'b10),
    .fci(\u2_Display/lt169_c31 ),
    .f({\u2_Display/n5434 ,open_n90324}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_0|u2_Display/lt170_cin  (
    .a({\u2_Display/n5468 ,1'b0}),
    .b({1'b0,open_n90330}),
    .fco(\u2_Display/lt170_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_10|u2_Display/lt170_9  (
    .a({\u2_Display/n5458 ,\u2_Display/n5459 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c9 ),
    .fco(\u2_Display/lt170_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_12|u2_Display/lt170_11  (
    .a({\u2_Display/n5456 ,\u2_Display/n5457 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c11 ),
    .fco(\u2_Display/lt170_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_14|u2_Display/lt170_13  (
    .a({\u2_Display/n5454 ,\u2_Display/n5455 }),
    .b(2'b01),
    .fci(\u2_Display/lt170_c13 ),
    .fco(\u2_Display/lt170_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_16|u2_Display/lt170_15  (
    .a({\u2_Display/n5452 ,\u2_Display/n5453 }),
    .b(2'b01),
    .fci(\u2_Display/lt170_c15 ),
    .fco(\u2_Display/lt170_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_18|u2_Display/lt170_17  (
    .a({\u2_Display/n5450 ,\u2_Display/n5451 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c17 ),
    .fco(\u2_Display/lt170_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_20|u2_Display/lt170_19  (
    .a({\u2_Display/n5448 ,\u2_Display/n5449 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c19 ),
    .fco(\u2_Display/lt170_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_22|u2_Display/lt170_21  (
    .a({\u2_Display/n5446 ,\u2_Display/n5447 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c21 ),
    .fco(\u2_Display/lt170_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_24|u2_Display/lt170_23  (
    .a({\u2_Display/n5444 ,\u2_Display/n5445 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c23 ),
    .fco(\u2_Display/lt170_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_26|u2_Display/lt170_25  (
    .a({\u2_Display/n5442 ,\u2_Display/n5443 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c25 ),
    .fco(\u2_Display/lt170_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_28|u2_Display/lt170_27  (
    .a({\u2_Display/n5440 ,\u2_Display/n5441 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c27 ),
    .fco(\u2_Display/lt170_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_2|u2_Display/lt170_1  (
    .a({\u2_Display/n5466 ,\u2_Display/n5467 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c1 ),
    .fco(\u2_Display/lt170_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_30|u2_Display/lt170_29  (
    .a({\u2_Display/n5438 ,\u2_Display/n5439 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c29 ),
    .fco(\u2_Display/lt170_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_4|u2_Display/lt170_3  (
    .a({\u2_Display/n5464 ,\u2_Display/n5465 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c3 ),
    .fco(\u2_Display/lt170_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_6|u2_Display/lt170_5  (
    .a({\u2_Display/n5462 ,\u2_Display/n5463 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c5 ),
    .fco(\u2_Display/lt170_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_8|u2_Display/lt170_7  (
    .a({\u2_Display/n5460 ,\u2_Display/n5461 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c7 ),
    .fco(\u2_Display/lt170_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_cout|u2_Display/lt170_31  (
    .a({1'b0,\u2_Display/n5437 }),
    .b(2'b10),
    .fci(\u2_Display/lt170_c31 ),
    .f({\u2_Display/n5469 ,open_n90734}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_0|u2_Display/lt171_cin  (
    .a({\u2_Display/n5503 ,1'b0}),
    .b({1'b0,open_n90740}),
    .fco(\u2_Display/lt171_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_10|u2_Display/lt171_9  (
    .a({\u2_Display/n5493 ,\u2_Display/n5494 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c9 ),
    .fco(\u2_Display/lt171_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_12|u2_Display/lt171_11  (
    .a({\u2_Display/n5491 ,\u2_Display/n5492 }),
    .b(2'b10),
    .fci(\u2_Display/lt171_c11 ),
    .fco(\u2_Display/lt171_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_14|u2_Display/lt171_13  (
    .a({\u2_Display/n5489 ,\u2_Display/n5490 }),
    .b(2'b10),
    .fci(\u2_Display/lt171_c13 ),
    .fco(\u2_Display/lt171_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_16|u2_Display/lt171_15  (
    .a({\u2_Display/n5487 ,\u2_Display/n5488 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c15 ),
    .fco(\u2_Display/lt171_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_18|u2_Display/lt171_17  (
    .a({\u2_Display/n5485 ,\u2_Display/n5486 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c17 ),
    .fco(\u2_Display/lt171_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_20|u2_Display/lt171_19  (
    .a({\u2_Display/n5483 ,\u2_Display/n5484 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c19 ),
    .fco(\u2_Display/lt171_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_22|u2_Display/lt171_21  (
    .a({\u2_Display/n5481 ,\u2_Display/n5482 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c21 ),
    .fco(\u2_Display/lt171_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_24|u2_Display/lt171_23  (
    .a({\u2_Display/n5479 ,\u2_Display/n5480 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c23 ),
    .fco(\u2_Display/lt171_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_26|u2_Display/lt171_25  (
    .a({\u2_Display/n5477 ,\u2_Display/n5478 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c25 ),
    .fco(\u2_Display/lt171_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_28|u2_Display/lt171_27  (
    .a({\u2_Display/n5475 ,\u2_Display/n5476 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c27 ),
    .fco(\u2_Display/lt171_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_2|u2_Display/lt171_1  (
    .a({\u2_Display/n5501 ,\u2_Display/n5502 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c1 ),
    .fco(\u2_Display/lt171_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_30|u2_Display/lt171_29  (
    .a({\u2_Display/n5473 ,\u2_Display/n5474 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c29 ),
    .fco(\u2_Display/lt171_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_4|u2_Display/lt171_3  (
    .a({\u2_Display/n5499 ,\u2_Display/n5500 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c3 ),
    .fco(\u2_Display/lt171_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_6|u2_Display/lt171_5  (
    .a({\u2_Display/n5497 ,\u2_Display/n5498 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c5 ),
    .fco(\u2_Display/lt171_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_8|u2_Display/lt171_7  (
    .a({\u2_Display/n5495 ,\u2_Display/n5496 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c7 ),
    .fco(\u2_Display/lt171_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_cout|u2_Display/lt171_31  (
    .a({1'b0,\u2_Display/n5472 }),
    .b(2'b10),
    .fci(\u2_Display/lt171_c31 ),
    .f({\u2_Display/n5504 ,open_n91144}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_0|u2_Display/lt172_cin  (
    .a({\u2_Display/n5538 ,1'b0}),
    .b({1'b0,open_n91150}),
    .fco(\u2_Display/lt172_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_10|u2_Display/lt172_9  (
    .a({\u2_Display/n5528 ,\u2_Display/n5529 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c9 ),
    .fco(\u2_Display/lt172_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_12|u2_Display/lt172_11  (
    .a({\u2_Display/n5526 ,\u2_Display/n5527 }),
    .b(2'b01),
    .fci(\u2_Display/lt172_c11 ),
    .fco(\u2_Display/lt172_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_14|u2_Display/lt172_13  (
    .a({\u2_Display/n5524 ,\u2_Display/n5525 }),
    .b(2'b01),
    .fci(\u2_Display/lt172_c13 ),
    .fco(\u2_Display/lt172_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_16|u2_Display/lt172_15  (
    .a({\u2_Display/n5522 ,\u2_Display/n5523 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c15 ),
    .fco(\u2_Display/lt172_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_18|u2_Display/lt172_17  (
    .a({\u2_Display/n5520 ,\u2_Display/n5521 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c17 ),
    .fco(\u2_Display/lt172_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_20|u2_Display/lt172_19  (
    .a({\u2_Display/n5518 ,\u2_Display/n5519 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c19 ),
    .fco(\u2_Display/lt172_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_22|u2_Display/lt172_21  (
    .a({\u2_Display/n5516 ,\u2_Display/n5517 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c21 ),
    .fco(\u2_Display/lt172_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_24|u2_Display/lt172_23  (
    .a({\u2_Display/n5514 ,\u2_Display/n5515 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c23 ),
    .fco(\u2_Display/lt172_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_26|u2_Display/lt172_25  (
    .a({\u2_Display/n5512 ,\u2_Display/n5513 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c25 ),
    .fco(\u2_Display/lt172_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_28|u2_Display/lt172_27  (
    .a({\u2_Display/n5510 ,\u2_Display/n5511 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c27 ),
    .fco(\u2_Display/lt172_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_2|u2_Display/lt172_1  (
    .a({\u2_Display/n5536 ,\u2_Display/n5537 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c1 ),
    .fco(\u2_Display/lt172_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_30|u2_Display/lt172_29  (
    .a({\u2_Display/n5508 ,\u2_Display/n5509 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c29 ),
    .fco(\u2_Display/lt172_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_4|u2_Display/lt172_3  (
    .a({\u2_Display/n5534 ,\u2_Display/n5535 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c3 ),
    .fco(\u2_Display/lt172_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_6|u2_Display/lt172_5  (
    .a({\u2_Display/n5532 ,\u2_Display/n5533 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c5 ),
    .fco(\u2_Display/lt172_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_8|u2_Display/lt172_7  (
    .a({\u2_Display/n5530 ,\u2_Display/n5531 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c7 ),
    .fco(\u2_Display/lt172_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_cout|u2_Display/lt172_31  (
    .a({1'b0,\u2_Display/n5507 }),
    .b(2'b10),
    .fci(\u2_Display/lt172_c31 ),
    .f({\u2_Display/n5539 ,open_n91554}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_0|u2_Display/lt173_cin  (
    .a({\u2_Display/n5573 ,1'b0}),
    .b({1'b0,open_n91560}),
    .fco(\u2_Display/lt173_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_10|u2_Display/lt173_9  (
    .a({\u2_Display/n5563 ,\u2_Display/n5564 }),
    .b(2'b10),
    .fci(\u2_Display/lt173_c9 ),
    .fco(\u2_Display/lt173_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_12|u2_Display/lt173_11  (
    .a({\u2_Display/n5561 ,\u2_Display/n5562 }),
    .b(2'b10),
    .fci(\u2_Display/lt173_c11 ),
    .fco(\u2_Display/lt173_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_14|u2_Display/lt173_13  (
    .a({\u2_Display/n5559 ,\u2_Display/n5560 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c13 ),
    .fco(\u2_Display/lt173_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_16|u2_Display/lt173_15  (
    .a({\u2_Display/n5557 ,\u2_Display/n5558 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c15 ),
    .fco(\u2_Display/lt173_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_18|u2_Display/lt173_17  (
    .a({\u2_Display/n5555 ,\u2_Display/n5556 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c17 ),
    .fco(\u2_Display/lt173_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_20|u2_Display/lt173_19  (
    .a({\u2_Display/n5553 ,\u2_Display/n5554 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c19 ),
    .fco(\u2_Display/lt173_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_22|u2_Display/lt173_21  (
    .a({\u2_Display/n5551 ,\u2_Display/n5552 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c21 ),
    .fco(\u2_Display/lt173_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_24|u2_Display/lt173_23  (
    .a({\u2_Display/n5549 ,\u2_Display/n5550 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c23 ),
    .fco(\u2_Display/lt173_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_26|u2_Display/lt173_25  (
    .a({\u2_Display/n5547 ,\u2_Display/n5548 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c25 ),
    .fco(\u2_Display/lt173_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_28|u2_Display/lt173_27  (
    .a({\u2_Display/n5545 ,\u2_Display/n5546 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c27 ),
    .fco(\u2_Display/lt173_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_2|u2_Display/lt173_1  (
    .a({\u2_Display/n5571 ,\u2_Display/n5572 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c1 ),
    .fco(\u2_Display/lt173_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_30|u2_Display/lt173_29  (
    .a({\u2_Display/n5543 ,\u2_Display/n5544 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c29 ),
    .fco(\u2_Display/lt173_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_4|u2_Display/lt173_3  (
    .a({\u2_Display/n5569 ,\u2_Display/n5570 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c3 ),
    .fco(\u2_Display/lt173_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_6|u2_Display/lt173_5  (
    .a({\u2_Display/n5567 ,\u2_Display/n5568 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c5 ),
    .fco(\u2_Display/lt173_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_8|u2_Display/lt173_7  (
    .a({\u2_Display/n5565 ,\u2_Display/n5566 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c7 ),
    .fco(\u2_Display/lt173_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_cout|u2_Display/lt173_31  (
    .a({1'b0,\u2_Display/n5542 }),
    .b(2'b10),
    .fci(\u2_Display/lt173_c31 ),
    .f({\u2_Display/n5574 ,open_n91964}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_0|u2_Display/lt174_cin  (
    .a({\u2_Display/n5608 ,1'b0}),
    .b({1'b0,open_n91970}),
    .fco(\u2_Display/lt174_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_10|u2_Display/lt174_9  (
    .a({\u2_Display/n5598 ,\u2_Display/n5599 }),
    .b(2'b01),
    .fci(\u2_Display/lt174_c9 ),
    .fco(\u2_Display/lt174_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_12|u2_Display/lt174_11  (
    .a({\u2_Display/n5596 ,\u2_Display/n5597 }),
    .b(2'b01),
    .fci(\u2_Display/lt174_c11 ),
    .fco(\u2_Display/lt174_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_14|u2_Display/lt174_13  (
    .a({\u2_Display/n5594 ,\u2_Display/n5595 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c13 ),
    .fco(\u2_Display/lt174_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_16|u2_Display/lt174_15  (
    .a({\u2_Display/n5592 ,\u2_Display/n5593 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c15 ),
    .fco(\u2_Display/lt174_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_18|u2_Display/lt174_17  (
    .a({\u2_Display/n5590 ,\u2_Display/n5591 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c17 ),
    .fco(\u2_Display/lt174_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_20|u2_Display/lt174_19  (
    .a({\u2_Display/n5588 ,\u2_Display/n5589 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c19 ),
    .fco(\u2_Display/lt174_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_22|u2_Display/lt174_21  (
    .a({\u2_Display/n5586 ,\u2_Display/n5587 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c21 ),
    .fco(\u2_Display/lt174_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_24|u2_Display/lt174_23  (
    .a({\u2_Display/n5584 ,\u2_Display/n5585 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c23 ),
    .fco(\u2_Display/lt174_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_26|u2_Display/lt174_25  (
    .a({\u2_Display/n5582 ,\u2_Display/n5583 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c25 ),
    .fco(\u2_Display/lt174_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_28|u2_Display/lt174_27  (
    .a({\u2_Display/n5580 ,\u2_Display/n5581 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c27 ),
    .fco(\u2_Display/lt174_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_2|u2_Display/lt174_1  (
    .a({\u2_Display/n5606 ,\u2_Display/n5607 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c1 ),
    .fco(\u2_Display/lt174_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_30|u2_Display/lt174_29  (
    .a({\u2_Display/n5578 ,\u2_Display/n5579 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c29 ),
    .fco(\u2_Display/lt174_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_4|u2_Display/lt174_3  (
    .a({\u2_Display/n5604 ,\u2_Display/n5605 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c3 ),
    .fco(\u2_Display/lt174_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_6|u2_Display/lt174_5  (
    .a({\u2_Display/n5602 ,\u2_Display/n5603 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c5 ),
    .fco(\u2_Display/lt174_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_8|u2_Display/lt174_7  (
    .a({\u2_Display/n5600 ,\u2_Display/n5601 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c7 ),
    .fco(\u2_Display/lt174_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_cout|u2_Display/lt174_31  (
    .a({1'b0,\u2_Display/n5577 }),
    .b(2'b10),
    .fci(\u2_Display/lt174_c31 ),
    .f({\u2_Display/n5609 ,open_n92374}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_0|u2_Display/lt175_cin  (
    .a({\u2_Display/n5643 ,1'b0}),
    .b({1'b0,open_n92380}),
    .fco(\u2_Display/lt175_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_10|u2_Display/lt175_9  (
    .a({\u2_Display/n5633 ,\u2_Display/n5634 }),
    .b(2'b10),
    .fci(\u2_Display/lt175_c9 ),
    .fco(\u2_Display/lt175_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_12|u2_Display/lt175_11  (
    .a({\u2_Display/n5631 ,\u2_Display/n5632 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c11 ),
    .fco(\u2_Display/lt175_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_14|u2_Display/lt175_13  (
    .a({\u2_Display/n5629 ,\u2_Display/n5630 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c13 ),
    .fco(\u2_Display/lt175_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_16|u2_Display/lt175_15  (
    .a({\u2_Display/n5627 ,\u2_Display/n5628 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c15 ),
    .fco(\u2_Display/lt175_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_18|u2_Display/lt175_17  (
    .a({\u2_Display/n5625 ,\u2_Display/n5626 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c17 ),
    .fco(\u2_Display/lt175_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_20|u2_Display/lt175_19  (
    .a({\u2_Display/n5623 ,\u2_Display/n5624 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c19 ),
    .fco(\u2_Display/lt175_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_22|u2_Display/lt175_21  (
    .a({\u2_Display/n5621 ,\u2_Display/n5622 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c21 ),
    .fco(\u2_Display/lt175_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_24|u2_Display/lt175_23  (
    .a({\u2_Display/n5619 ,\u2_Display/n5620 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c23 ),
    .fco(\u2_Display/lt175_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_26|u2_Display/lt175_25  (
    .a({\u2_Display/n5617 ,\u2_Display/n5618 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c25 ),
    .fco(\u2_Display/lt175_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_28|u2_Display/lt175_27  (
    .a({\u2_Display/n5615 ,\u2_Display/n5616 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c27 ),
    .fco(\u2_Display/lt175_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_2|u2_Display/lt175_1  (
    .a({\u2_Display/n5641 ,\u2_Display/n5642 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c1 ),
    .fco(\u2_Display/lt175_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_30|u2_Display/lt175_29  (
    .a({\u2_Display/n5613 ,\u2_Display/n5614 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c29 ),
    .fco(\u2_Display/lt175_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_4|u2_Display/lt175_3  (
    .a({\u2_Display/n5639 ,\u2_Display/n5640 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c3 ),
    .fco(\u2_Display/lt175_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_6|u2_Display/lt175_5  (
    .a({\u2_Display/n5637 ,\u2_Display/n5638 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c5 ),
    .fco(\u2_Display/lt175_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_8|u2_Display/lt175_7  (
    .a({\u2_Display/n5635 ,\u2_Display/n5636 }),
    .b(2'b10),
    .fci(\u2_Display/lt175_c7 ),
    .fco(\u2_Display/lt175_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_cout|u2_Display/lt175_31  (
    .a({1'b0,\u2_Display/n5612 }),
    .b(2'b10),
    .fci(\u2_Display/lt175_c31 ),
    .f({\u2_Display/n5644 ,open_n92784}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_0|u2_Display/lt176_cin  (
    .a({\u2_Display/n5678 ,1'b0}),
    .b({1'b0,open_n92790}),
    .fco(\u2_Display/lt176_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_10|u2_Display/lt176_9  (
    .a({\u2_Display/n5668 ,\u2_Display/n5669 }),
    .b(2'b01),
    .fci(\u2_Display/lt176_c9 ),
    .fco(\u2_Display/lt176_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_12|u2_Display/lt176_11  (
    .a({\u2_Display/n5666 ,\u2_Display/n5667 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c11 ),
    .fco(\u2_Display/lt176_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_14|u2_Display/lt176_13  (
    .a({\u2_Display/n5664 ,\u2_Display/n5665 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c13 ),
    .fco(\u2_Display/lt176_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_16|u2_Display/lt176_15  (
    .a({\u2_Display/n5662 ,\u2_Display/n5663 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c15 ),
    .fco(\u2_Display/lt176_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_18|u2_Display/lt176_17  (
    .a({\u2_Display/n5660 ,\u2_Display/n5661 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c17 ),
    .fco(\u2_Display/lt176_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_20|u2_Display/lt176_19  (
    .a({\u2_Display/n5658 ,\u2_Display/n5659 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c19 ),
    .fco(\u2_Display/lt176_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_22|u2_Display/lt176_21  (
    .a({\u2_Display/n5656 ,\u2_Display/n5657 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c21 ),
    .fco(\u2_Display/lt176_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_24|u2_Display/lt176_23  (
    .a({\u2_Display/n5654 ,\u2_Display/n5655 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c23 ),
    .fco(\u2_Display/lt176_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_26|u2_Display/lt176_25  (
    .a({\u2_Display/n5652 ,\u2_Display/n5653 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c25 ),
    .fco(\u2_Display/lt176_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_28|u2_Display/lt176_27  (
    .a({\u2_Display/n5650 ,\u2_Display/n5651 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c27 ),
    .fco(\u2_Display/lt176_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_2|u2_Display/lt176_1  (
    .a({\u2_Display/n5676 ,\u2_Display/n5677 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c1 ),
    .fco(\u2_Display/lt176_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_30|u2_Display/lt176_29  (
    .a({\u2_Display/n5648 ,\u2_Display/n5649 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c29 ),
    .fco(\u2_Display/lt176_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_4|u2_Display/lt176_3  (
    .a({\u2_Display/n5674 ,\u2_Display/n5675 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c3 ),
    .fco(\u2_Display/lt176_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_6|u2_Display/lt176_5  (
    .a({\u2_Display/n5672 ,\u2_Display/n5673 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c5 ),
    .fco(\u2_Display/lt176_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_8|u2_Display/lt176_7  (
    .a({\u2_Display/n5670 ,\u2_Display/n5671 }),
    .b(2'b01),
    .fci(\u2_Display/lt176_c7 ),
    .fco(\u2_Display/lt176_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_cout|u2_Display/lt176_31  (
    .a({1'b0,\u2_Display/n5647 }),
    .b(2'b10),
    .fci(\u2_Display/lt176_c31 ),
    .f({\u2_Display/n5679 ,open_n93194}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_0|u2_Display/lt1_cin  (
    .a({\u2_Display/i [0],1'b0}),
    .b({lcd_xpos[0],open_n93200}),
    .fco(\u2_Display/lt1_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_10|u2_Display/lt1_9  (
    .a(\u2_Display/i [10:9]),
    .b(lcd_xpos[10:9]),
    .fci(\u2_Display/lt1_c9 ),
    .fco(\u2_Display/lt1_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_2|u2_Display/lt1_1  (
    .a(\u2_Display/i [2:1]),
    .b(lcd_xpos[2:1]),
    .fci(\u2_Display/lt1_c1 ),
    .fco(\u2_Display/lt1_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_4|u2_Display/lt1_3  (
    .a(\u2_Display/i [4:3]),
    .b(lcd_xpos[4:3]),
    .fci(\u2_Display/lt1_c3 ),
    .fco(\u2_Display/lt1_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_6|u2_Display/lt1_5  (
    .a(\u2_Display/i [6:5]),
    .b(lcd_xpos[6:5]),
    .fci(\u2_Display/lt1_c5 ),
    .fco(\u2_Display/lt1_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_8|u2_Display/lt1_7  (
    .a(\u2_Display/i [8:7]),
    .b(lcd_xpos[8:7]),
    .fci(\u2_Display/lt1_c7 ),
    .fco(\u2_Display/lt1_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_cout|u2_Display/lt1_11  (
    .a(2'b00),
    .b({1'b1,lcd_xpos[11]}),
    .fci(\u2_Display/lt1_c11 ),
    .f({\u2_Display/n45 ,open_n93364}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_0|u2_Display/lt22_cin  (
    .a({\u2_Display/counta [0],1'b0}),
    .b({1'b0,open_n93370}),
    .fco(\u2_Display/lt22_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_10|u2_Display/lt22_9  (
    .a(\u2_Display/counta [10:9]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c9 ),
    .fco(\u2_Display/lt22_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_12|u2_Display/lt22_11  (
    .a(\u2_Display/counta [12:11]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c11 ),
    .fco(\u2_Display/lt22_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_14|u2_Display/lt22_13  (
    .a(\u2_Display/counta [14:13]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c13 ),
    .fco(\u2_Display/lt22_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_16|u2_Display/lt22_15  (
    .a(\u2_Display/counta [16:15]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c15 ),
    .fco(\u2_Display/lt22_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_18|u2_Display/lt22_17  (
    .a(\u2_Display/counta [18:17]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c17 ),
    .fco(\u2_Display/lt22_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_20|u2_Display/lt22_19  (
    .a(\u2_Display/counta [20:19]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c19 ),
    .fco(\u2_Display/lt22_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_22|u2_Display/lt22_21  (
    .a(\u2_Display/counta [22:21]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c21 ),
    .fco(\u2_Display/lt22_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_24|u2_Display/lt22_23  (
    .a(\u2_Display/counta [24:23]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c23 ),
    .fco(\u2_Display/lt22_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_26|u2_Display/lt22_25  (
    .a(\u2_Display/counta [26:25]),
    .b(2'b01),
    .fci(\u2_Display/lt22_c25 ),
    .fco(\u2_Display/lt22_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_28|u2_Display/lt22_27  (
    .a(\u2_Display/counta [28:27]),
    .b(2'b11),
    .fci(\u2_Display/lt22_c27 ),
    .fco(\u2_Display/lt22_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_2|u2_Display/lt22_1  (
    .a(\u2_Display/counta [2:1]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c1 ),
    .fco(\u2_Display/lt22_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_30|u2_Display/lt22_29  (
    .a(\u2_Display/counta [30:29]),
    .b(2'b11),
    .fci(\u2_Display/lt22_c29 ),
    .fco(\u2_Display/lt22_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_4|u2_Display/lt22_3  (
    .a(\u2_Display/counta [4:3]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c3 ),
    .fco(\u2_Display/lt22_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_6|u2_Display/lt22_5  (
    .a(\u2_Display/counta [6:5]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c5 ),
    .fco(\u2_Display/lt22_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_8|u2_Display/lt22_7  (
    .a(\u2_Display/counta [8:7]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c7 ),
    .fco(\u2_Display/lt22_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_cout|u2_Display/lt22_31  (
    .a({1'b0,\u2_Display/counta [31]}),
    .b(2'b11),
    .fci(\u2_Display/lt22_c31 ),
    .f({\u2_Display/n417 ,open_n93774}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_0|u2_Display/lt23_cin  (
    .a({\u2_Display/n451 ,1'b0}),
    .b({1'b0,open_n93780}),
    .fco(\u2_Display/lt23_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_10|u2_Display/lt23_9  (
    .a({\u2_Display/n441 ,\u2_Display/n442 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c9 ),
    .fco(\u2_Display/lt23_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_12|u2_Display/lt23_11  (
    .a({\u2_Display/n439 ,\u2_Display/n440 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c11 ),
    .fco(\u2_Display/lt23_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_14|u2_Display/lt23_13  (
    .a({\u2_Display/n437 ,\u2_Display/n438 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c13 ),
    .fco(\u2_Display/lt23_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_16|u2_Display/lt23_15  (
    .a({\u2_Display/n435 ,\u2_Display/n436 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c15 ),
    .fco(\u2_Display/lt23_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_18|u2_Display/lt23_17  (
    .a({\u2_Display/n433 ,\u2_Display/n434 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c17 ),
    .fco(\u2_Display/lt23_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_20|u2_Display/lt23_19  (
    .a({\u2_Display/n431 ,\u2_Display/n432 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c19 ),
    .fco(\u2_Display/lt23_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_22|u2_Display/lt23_21  (
    .a({\u2_Display/n429 ,\u2_Display/n430 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c21 ),
    .fco(\u2_Display/lt23_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_24|u2_Display/lt23_23  (
    .a({\u2_Display/n427 ,\u2_Display/n428 }),
    .b(2'b10),
    .fci(\u2_Display/lt23_c23 ),
    .fco(\u2_Display/lt23_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_26|u2_Display/lt23_25  (
    .a({\u2_Display/n425 ,\u2_Display/n426 }),
    .b(2'b10),
    .fci(\u2_Display/lt23_c25 ),
    .fco(\u2_Display/lt23_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_28|u2_Display/lt23_27  (
    .a({\u2_Display/n423 ,\u2_Display/n424 }),
    .b(2'b11),
    .fci(\u2_Display/lt23_c27 ),
    .fco(\u2_Display/lt23_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_2|u2_Display/lt23_1  (
    .a({\u2_Display/n449 ,\u2_Display/n450 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c1 ),
    .fco(\u2_Display/lt23_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_30|u2_Display/lt23_29  (
    .a({\u2_Display/n421 ,\u2_Display/n422 }),
    .b(2'b11),
    .fci(\u2_Display/lt23_c29 ),
    .fco(\u2_Display/lt23_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_4|u2_Display/lt23_3  (
    .a({\u2_Display/n447 ,\u2_Display/n448 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c3 ),
    .fco(\u2_Display/lt23_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_6|u2_Display/lt23_5  (
    .a({\u2_Display/n445 ,\u2_Display/n446 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c5 ),
    .fco(\u2_Display/lt23_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_8|u2_Display/lt23_7  (
    .a({\u2_Display/n443 ,\u2_Display/n444 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c7 ),
    .fco(\u2_Display/lt23_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_cout|u2_Display/lt23_31  (
    .a({1'b0,\u2_Display/n420 }),
    .b(2'b10),
    .fci(\u2_Display/lt23_c31 ),
    .f({\u2_Display/n452 ,open_n94184}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_0|u2_Display/lt24_cin  (
    .a({\u2_Display/n486 ,1'b0}),
    .b({1'b0,open_n94190}),
    .fco(\u2_Display/lt24_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_10|u2_Display/lt24_9  (
    .a({\u2_Display/n476 ,\u2_Display/n477 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c9 ),
    .fco(\u2_Display/lt24_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_12|u2_Display/lt24_11  (
    .a({\u2_Display/n474 ,\u2_Display/n475 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c11 ),
    .fco(\u2_Display/lt24_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_14|u2_Display/lt24_13  (
    .a({\u2_Display/n472 ,\u2_Display/n473 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c13 ),
    .fco(\u2_Display/lt24_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_16|u2_Display/lt24_15  (
    .a({\u2_Display/n470 ,\u2_Display/n471 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c15 ),
    .fco(\u2_Display/lt24_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_18|u2_Display/lt24_17  (
    .a({\u2_Display/n468 ,\u2_Display/n469 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c17 ),
    .fco(\u2_Display/lt24_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_20|u2_Display/lt24_19  (
    .a({\u2_Display/n466 ,\u2_Display/n467 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c19 ),
    .fco(\u2_Display/lt24_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_22|u2_Display/lt24_21  (
    .a({\u2_Display/n464 ,\u2_Display/n465 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c21 ),
    .fco(\u2_Display/lt24_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_24|u2_Display/lt24_23  (
    .a({\u2_Display/n462 ,\u2_Display/n463 }),
    .b(2'b01),
    .fci(\u2_Display/lt24_c23 ),
    .fco(\u2_Display/lt24_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_26|u2_Display/lt24_25  (
    .a({\u2_Display/n460 ,\u2_Display/n461 }),
    .b(2'b11),
    .fci(\u2_Display/lt24_c25 ),
    .fco(\u2_Display/lt24_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_28|u2_Display/lt24_27  (
    .a({\u2_Display/n458 ,\u2_Display/n459 }),
    .b(2'b11),
    .fci(\u2_Display/lt24_c27 ),
    .fco(\u2_Display/lt24_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_2|u2_Display/lt24_1  (
    .a({\u2_Display/n484 ,\u2_Display/n485 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c1 ),
    .fco(\u2_Display/lt24_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_30|u2_Display/lt24_29  (
    .a({\u2_Display/n456 ,\u2_Display/n457 }),
    .b(2'b01),
    .fci(\u2_Display/lt24_c29 ),
    .fco(\u2_Display/lt24_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_4|u2_Display/lt24_3  (
    .a({\u2_Display/n482 ,\u2_Display/n483 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c3 ),
    .fco(\u2_Display/lt24_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_6|u2_Display/lt24_5  (
    .a({\u2_Display/n480 ,\u2_Display/n481 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c5 ),
    .fco(\u2_Display/lt24_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_8|u2_Display/lt24_7  (
    .a({\u2_Display/n478 ,\u2_Display/n479 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c7 ),
    .fco(\u2_Display/lt24_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_cout|u2_Display/lt24_31  (
    .a({1'b0,\u2_Display/n455 }),
    .b(2'b10),
    .fci(\u2_Display/lt24_c31 ),
    .f({\u2_Display/n487 ,open_n94594}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_0|u2_Display/lt25_cin  (
    .a({\u2_Display/n521 ,1'b0}),
    .b({1'b0,open_n94600}),
    .fco(\u2_Display/lt25_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_10|u2_Display/lt25_9  (
    .a({\u2_Display/n511 ,\u2_Display/n512 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c9 ),
    .fco(\u2_Display/lt25_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_12|u2_Display/lt25_11  (
    .a({\u2_Display/n509 ,\u2_Display/n510 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c11 ),
    .fco(\u2_Display/lt25_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_14|u2_Display/lt25_13  (
    .a({\u2_Display/n507 ,\u2_Display/n508 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c13 ),
    .fco(\u2_Display/lt25_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_16|u2_Display/lt25_15  (
    .a({\u2_Display/n505 ,\u2_Display/n506 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c15 ),
    .fco(\u2_Display/lt25_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_18|u2_Display/lt25_17  (
    .a({\u2_Display/n503 ,\u2_Display/n504 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c17 ),
    .fco(\u2_Display/lt25_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_20|u2_Display/lt25_19  (
    .a({\u2_Display/n501 ,\u2_Display/n502 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c19 ),
    .fco(\u2_Display/lt25_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_22|u2_Display/lt25_21  (
    .a({\u2_Display/n499 ,\u2_Display/n500 }),
    .b(2'b10),
    .fci(\u2_Display/lt25_c21 ),
    .fco(\u2_Display/lt25_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_24|u2_Display/lt25_23  (
    .a({\u2_Display/n497 ,\u2_Display/n498 }),
    .b(2'b10),
    .fci(\u2_Display/lt25_c23 ),
    .fco(\u2_Display/lt25_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_26|u2_Display/lt25_25  (
    .a({\u2_Display/n495 ,\u2_Display/n496 }),
    .b(2'b11),
    .fci(\u2_Display/lt25_c25 ),
    .fco(\u2_Display/lt25_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_28|u2_Display/lt25_27  (
    .a({\u2_Display/n493 ,\u2_Display/n494 }),
    .b(2'b11),
    .fci(\u2_Display/lt25_c27 ),
    .fco(\u2_Display/lt25_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_2|u2_Display/lt25_1  (
    .a({\u2_Display/n519 ,\u2_Display/n520 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c1 ),
    .fco(\u2_Display/lt25_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_30|u2_Display/lt25_29  (
    .a({\u2_Display/n491 ,\u2_Display/n492 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c29 ),
    .fco(\u2_Display/lt25_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_4|u2_Display/lt25_3  (
    .a({\u2_Display/n517 ,\u2_Display/n518 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c3 ),
    .fco(\u2_Display/lt25_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_6|u2_Display/lt25_5  (
    .a({\u2_Display/n515 ,\u2_Display/n516 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c5 ),
    .fco(\u2_Display/lt25_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_8|u2_Display/lt25_7  (
    .a({\u2_Display/n513 ,\u2_Display/n514 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c7 ),
    .fco(\u2_Display/lt25_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_cout|u2_Display/lt25_31  (
    .a({1'b0,\u2_Display/n490 }),
    .b(2'b10),
    .fci(\u2_Display/lt25_c31 ),
    .f({\u2_Display/n522 ,open_n95004}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_0|u2_Display/lt26_cin  (
    .a({\u2_Display/n556 ,1'b0}),
    .b({1'b0,open_n95010}),
    .fco(\u2_Display/lt26_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_10|u2_Display/lt26_9  (
    .a({\u2_Display/n546 ,\u2_Display/n547 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c9 ),
    .fco(\u2_Display/lt26_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_12|u2_Display/lt26_11  (
    .a({\u2_Display/n544 ,\u2_Display/n545 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c11 ),
    .fco(\u2_Display/lt26_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_14|u2_Display/lt26_13  (
    .a({\u2_Display/n542 ,\u2_Display/n543 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c13 ),
    .fco(\u2_Display/lt26_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_16|u2_Display/lt26_15  (
    .a({\u2_Display/n540 ,\u2_Display/n541 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c15 ),
    .fco(\u2_Display/lt26_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_18|u2_Display/lt26_17  (
    .a({\u2_Display/n538 ,\u2_Display/n539 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c17 ),
    .fco(\u2_Display/lt26_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_20|u2_Display/lt26_19  (
    .a({\u2_Display/n536 ,\u2_Display/n537 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c19 ),
    .fco(\u2_Display/lt26_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_22|u2_Display/lt26_21  (
    .a({\u2_Display/n534 ,\u2_Display/n535 }),
    .b(2'b01),
    .fci(\u2_Display/lt26_c21 ),
    .fco(\u2_Display/lt26_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_24|u2_Display/lt26_23  (
    .a({\u2_Display/n532 ,\u2_Display/n533 }),
    .b(2'b11),
    .fci(\u2_Display/lt26_c23 ),
    .fco(\u2_Display/lt26_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_26|u2_Display/lt26_25  (
    .a({\u2_Display/n530 ,\u2_Display/n531 }),
    .b(2'b11),
    .fci(\u2_Display/lt26_c25 ),
    .fco(\u2_Display/lt26_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_28|u2_Display/lt26_27  (
    .a({\u2_Display/n528 ,\u2_Display/n529 }),
    .b(2'b01),
    .fci(\u2_Display/lt26_c27 ),
    .fco(\u2_Display/lt26_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_2|u2_Display/lt26_1  (
    .a({\u2_Display/n554 ,\u2_Display/n555 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c1 ),
    .fco(\u2_Display/lt26_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_30|u2_Display/lt26_29  (
    .a({\u2_Display/n526 ,\u2_Display/n527 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c29 ),
    .fco(\u2_Display/lt26_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_4|u2_Display/lt26_3  (
    .a({\u2_Display/n552 ,\u2_Display/n553 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c3 ),
    .fco(\u2_Display/lt26_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_6|u2_Display/lt26_5  (
    .a({\u2_Display/n550 ,\u2_Display/n551 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c5 ),
    .fco(\u2_Display/lt26_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_8|u2_Display/lt26_7  (
    .a({\u2_Display/n548 ,\u2_Display/n549 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c7 ),
    .fco(\u2_Display/lt26_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_cout|u2_Display/lt26_31  (
    .a({1'b0,\u2_Display/n525 }),
    .b(2'b10),
    .fci(\u2_Display/lt26_c31 ),
    .f({\u2_Display/n557 ,open_n95414}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_0|u2_Display/lt27_cin  (
    .a({\u2_Display/n591 ,1'b0}),
    .b({1'b0,open_n95420}),
    .fco(\u2_Display/lt27_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_10|u2_Display/lt27_9  (
    .a({\u2_Display/n581 ,\u2_Display/n582 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c9 ),
    .fco(\u2_Display/lt27_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_12|u2_Display/lt27_11  (
    .a({\u2_Display/n579 ,\u2_Display/n580 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c11 ),
    .fco(\u2_Display/lt27_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_14|u2_Display/lt27_13  (
    .a({\u2_Display/n577 ,\u2_Display/n578 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c13 ),
    .fco(\u2_Display/lt27_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_16|u2_Display/lt27_15  (
    .a({\u2_Display/n575 ,\u2_Display/n576 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c15 ),
    .fco(\u2_Display/lt27_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_18|u2_Display/lt27_17  (
    .a({\u2_Display/n573 ,\u2_Display/n574 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c17 ),
    .fco(\u2_Display/lt27_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_20|u2_Display/lt27_19  (
    .a({\u2_Display/n571 ,\u2_Display/n572 }),
    .b(2'b10),
    .fci(\u2_Display/lt27_c19 ),
    .fco(\u2_Display/lt27_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_22|u2_Display/lt27_21  (
    .a({\u2_Display/n569 ,\u2_Display/n570 }),
    .b(2'b10),
    .fci(\u2_Display/lt27_c21 ),
    .fco(\u2_Display/lt27_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_24|u2_Display/lt27_23  (
    .a({\u2_Display/n567 ,\u2_Display/n568 }),
    .b(2'b11),
    .fci(\u2_Display/lt27_c23 ),
    .fco(\u2_Display/lt27_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_26|u2_Display/lt27_25  (
    .a({\u2_Display/n565 ,\u2_Display/n566 }),
    .b(2'b11),
    .fci(\u2_Display/lt27_c25 ),
    .fco(\u2_Display/lt27_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_28|u2_Display/lt27_27  (
    .a({\u2_Display/n563 ,\u2_Display/n564 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c27 ),
    .fco(\u2_Display/lt27_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_2|u2_Display/lt27_1  (
    .a({\u2_Display/n589 ,\u2_Display/n590 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c1 ),
    .fco(\u2_Display/lt27_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_30|u2_Display/lt27_29  (
    .a({\u2_Display/n561 ,\u2_Display/n562 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c29 ),
    .fco(\u2_Display/lt27_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_4|u2_Display/lt27_3  (
    .a({\u2_Display/n587 ,\u2_Display/n588 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c3 ),
    .fco(\u2_Display/lt27_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_6|u2_Display/lt27_5  (
    .a({\u2_Display/n585 ,\u2_Display/n586 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c5 ),
    .fco(\u2_Display/lt27_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_8|u2_Display/lt27_7  (
    .a({\u2_Display/n583 ,\u2_Display/n584 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c7 ),
    .fco(\u2_Display/lt27_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_cout|u2_Display/lt27_31  (
    .a({1'b0,\u2_Display/n560 }),
    .b(2'b10),
    .fci(\u2_Display/lt27_c31 ),
    .f({\u2_Display/n592 ,open_n95824}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_0|u2_Display/lt28_cin  (
    .a({\u2_Display/n626 ,1'b0}),
    .b({1'b0,open_n95830}),
    .fco(\u2_Display/lt28_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_10|u2_Display/lt28_9  (
    .a({\u2_Display/n616 ,\u2_Display/n617 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c9 ),
    .fco(\u2_Display/lt28_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_12|u2_Display/lt28_11  (
    .a({\u2_Display/n614 ,\u2_Display/n615 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c11 ),
    .fco(\u2_Display/lt28_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_14|u2_Display/lt28_13  (
    .a({\u2_Display/n612 ,\u2_Display/n613 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c13 ),
    .fco(\u2_Display/lt28_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_16|u2_Display/lt28_15  (
    .a({\u2_Display/n610 ,\u2_Display/n611 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c15 ),
    .fco(\u2_Display/lt28_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_18|u2_Display/lt28_17  (
    .a({\u2_Display/n608 ,\u2_Display/n609 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c17 ),
    .fco(\u2_Display/lt28_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_20|u2_Display/lt28_19  (
    .a({\u2_Display/n606 ,\u2_Display/n607 }),
    .b(2'b01),
    .fci(\u2_Display/lt28_c19 ),
    .fco(\u2_Display/lt28_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_22|u2_Display/lt28_21  (
    .a({\u2_Display/n604 ,\u2_Display/n605 }),
    .b(2'b11),
    .fci(\u2_Display/lt28_c21 ),
    .fco(\u2_Display/lt28_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_24|u2_Display/lt28_23  (
    .a({\u2_Display/n602 ,\u2_Display/n603 }),
    .b(2'b11),
    .fci(\u2_Display/lt28_c23 ),
    .fco(\u2_Display/lt28_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_26|u2_Display/lt28_25  (
    .a({\u2_Display/n600 ,\u2_Display/n601 }),
    .b(2'b01),
    .fci(\u2_Display/lt28_c25 ),
    .fco(\u2_Display/lt28_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_28|u2_Display/lt28_27  (
    .a({\u2_Display/n598 ,\u2_Display/n599 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c27 ),
    .fco(\u2_Display/lt28_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_2|u2_Display/lt28_1  (
    .a({\u2_Display/n624 ,\u2_Display/n625 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c1 ),
    .fco(\u2_Display/lt28_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_30|u2_Display/lt28_29  (
    .a({\u2_Display/n596 ,\u2_Display/n597 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c29 ),
    .fco(\u2_Display/lt28_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_4|u2_Display/lt28_3  (
    .a({\u2_Display/n622 ,\u2_Display/n623 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c3 ),
    .fco(\u2_Display/lt28_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_6|u2_Display/lt28_5  (
    .a({\u2_Display/n620 ,\u2_Display/n621 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c5 ),
    .fco(\u2_Display/lt28_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_8|u2_Display/lt28_7  (
    .a({\u2_Display/n618 ,\u2_Display/n619 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c7 ),
    .fco(\u2_Display/lt28_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_cout|u2_Display/lt28_31  (
    .a({1'b0,\u2_Display/n595 }),
    .b(2'b10),
    .fci(\u2_Display/lt28_c31 ),
    .f({\u2_Display/n627 ,open_n96234}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_0|u2_Display/lt29_cin  (
    .a({\u2_Display/n661 ,1'b0}),
    .b({1'b0,open_n96240}),
    .fco(\u2_Display/lt29_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_10|u2_Display/lt29_9  (
    .a({\u2_Display/n651 ,\u2_Display/n652 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c9 ),
    .fco(\u2_Display/lt29_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_12|u2_Display/lt29_11  (
    .a({\u2_Display/n649 ,\u2_Display/n650 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c11 ),
    .fco(\u2_Display/lt29_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_14|u2_Display/lt29_13  (
    .a({\u2_Display/n647 ,\u2_Display/n648 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c13 ),
    .fco(\u2_Display/lt29_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_16|u2_Display/lt29_15  (
    .a({\u2_Display/n645 ,\u2_Display/n646 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c15 ),
    .fco(\u2_Display/lt29_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_18|u2_Display/lt29_17  (
    .a({\u2_Display/n643 ,\u2_Display/n644 }),
    .b(2'b10),
    .fci(\u2_Display/lt29_c17 ),
    .fco(\u2_Display/lt29_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_20|u2_Display/lt29_19  (
    .a({\u2_Display/n641 ,\u2_Display/n642 }),
    .b(2'b10),
    .fci(\u2_Display/lt29_c19 ),
    .fco(\u2_Display/lt29_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_22|u2_Display/lt29_21  (
    .a({\u2_Display/n639 ,\u2_Display/n640 }),
    .b(2'b11),
    .fci(\u2_Display/lt29_c21 ),
    .fco(\u2_Display/lt29_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_24|u2_Display/lt29_23  (
    .a({\u2_Display/n637 ,\u2_Display/n638 }),
    .b(2'b11),
    .fci(\u2_Display/lt29_c23 ),
    .fco(\u2_Display/lt29_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_26|u2_Display/lt29_25  (
    .a({\u2_Display/n635 ,\u2_Display/n636 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c25 ),
    .fco(\u2_Display/lt29_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_28|u2_Display/lt29_27  (
    .a({\u2_Display/n633 ,\u2_Display/n634 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c27 ),
    .fco(\u2_Display/lt29_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_2|u2_Display/lt29_1  (
    .a({\u2_Display/n659 ,\u2_Display/n660 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c1 ),
    .fco(\u2_Display/lt29_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_30|u2_Display/lt29_29  (
    .a({\u2_Display/n631 ,\u2_Display/n632 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c29 ),
    .fco(\u2_Display/lt29_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_4|u2_Display/lt29_3  (
    .a({\u2_Display/n657 ,\u2_Display/n658 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c3 ),
    .fco(\u2_Display/lt29_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_6|u2_Display/lt29_5  (
    .a({\u2_Display/n655 ,\u2_Display/n656 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c5 ),
    .fco(\u2_Display/lt29_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_8|u2_Display/lt29_7  (
    .a({\u2_Display/n653 ,\u2_Display/n654 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c7 ),
    .fco(\u2_Display/lt29_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_cout|u2_Display/lt29_31  (
    .a({1'b0,\u2_Display/n630 }),
    .b(2'b10),
    .fci(\u2_Display/lt29_c31 ),
    .f({\u2_Display/n662 ,open_n96644}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_0|u2_Display/lt2_2_cin  (
    .a({lcd_ypos[0],1'b0}),
    .b({\u2_Display/j [0],open_n96650}),
    .fco(\u2_Display/lt2_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_10|u2_Display/lt2_2_9  (
    .a(lcd_ypos[10:9]),
    .b({1'b1,\u2_Display/j [9]}),
    .fci(\u2_Display/lt2_2_c9 ),
    .fco(\u2_Display/lt2_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_2|u2_Display/lt2_2_1  (
    .a(lcd_ypos[2:1]),
    .b(\u2_Display/j [2:1]),
    .fci(\u2_Display/lt2_2_c1 ),
    .fco(\u2_Display/lt2_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_4|u2_Display/lt2_2_3  (
    .a(lcd_ypos[4:3]),
    .b(\u2_Display/j [4:3]),
    .fci(\u2_Display/lt2_2_c3 ),
    .fco(\u2_Display/lt2_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_6|u2_Display/lt2_2_5  (
    .a(lcd_ypos[6:5]),
    .b(\u2_Display/j [6:5]),
    .fci(\u2_Display/lt2_2_c5 ),
    .fco(\u2_Display/lt2_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_8|u2_Display/lt2_2_7  (
    .a(lcd_ypos[8:7]),
    .b(\u2_Display/j [8:7]),
    .fci(\u2_Display/lt2_2_c7 ),
    .fco(\u2_Display/lt2_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_cout|u2_Display/lt2_2_11  (
    .a({1'b0,lcd_ypos[11]}),
    .b(2'b10),
    .fci(\u2_Display/lt2_2_c11 ),
    .f({\u2_Display/n48 ,open_n96814}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_0|u2_Display/lt30_cin  (
    .a({\u2_Display/n696 ,1'b0}),
    .b({1'b0,open_n96820}),
    .fco(\u2_Display/lt30_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_10|u2_Display/lt30_9  (
    .a({\u2_Display/n686 ,\u2_Display/n687 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c9 ),
    .fco(\u2_Display/lt30_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_12|u2_Display/lt30_11  (
    .a({\u2_Display/n684 ,\u2_Display/n685 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c11 ),
    .fco(\u2_Display/lt30_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_14|u2_Display/lt30_13  (
    .a({\u2_Display/n682 ,\u2_Display/n683 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c13 ),
    .fco(\u2_Display/lt30_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_16|u2_Display/lt30_15  (
    .a({\u2_Display/n680 ,\u2_Display/n681 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c15 ),
    .fco(\u2_Display/lt30_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_18|u2_Display/lt30_17  (
    .a({\u2_Display/n678 ,\u2_Display/n679 }),
    .b(2'b01),
    .fci(\u2_Display/lt30_c17 ),
    .fco(\u2_Display/lt30_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_20|u2_Display/lt30_19  (
    .a({\u2_Display/n676 ,\u2_Display/n677 }),
    .b(2'b11),
    .fci(\u2_Display/lt30_c19 ),
    .fco(\u2_Display/lt30_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_22|u2_Display/lt30_21  (
    .a({\u2_Display/n674 ,\u2_Display/n675 }),
    .b(2'b11),
    .fci(\u2_Display/lt30_c21 ),
    .fco(\u2_Display/lt30_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_24|u2_Display/lt30_23  (
    .a({\u2_Display/n672 ,\u2_Display/n673 }),
    .b(2'b01),
    .fci(\u2_Display/lt30_c23 ),
    .fco(\u2_Display/lt30_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_26|u2_Display/lt30_25  (
    .a({\u2_Display/n670 ,\u2_Display/n671 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c25 ),
    .fco(\u2_Display/lt30_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_28|u2_Display/lt30_27  (
    .a({\u2_Display/n668 ,\u2_Display/n669 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c27 ),
    .fco(\u2_Display/lt30_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_2|u2_Display/lt30_1  (
    .a({\u2_Display/n694 ,\u2_Display/n695 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c1 ),
    .fco(\u2_Display/lt30_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_30|u2_Display/lt30_29  (
    .a({\u2_Display/n666 ,\u2_Display/n667 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c29 ),
    .fco(\u2_Display/lt30_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_4|u2_Display/lt30_3  (
    .a({\u2_Display/n692 ,\u2_Display/n693 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c3 ),
    .fco(\u2_Display/lt30_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_6|u2_Display/lt30_5  (
    .a({\u2_Display/n690 ,\u2_Display/n691 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c5 ),
    .fco(\u2_Display/lt30_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_8|u2_Display/lt30_7  (
    .a({\u2_Display/n688 ,\u2_Display/n689 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c7 ),
    .fco(\u2_Display/lt30_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_cout|u2_Display/lt30_31  (
    .a({1'b0,\u2_Display/n665 }),
    .b(2'b10),
    .fci(\u2_Display/lt30_c31 ),
    .f({\u2_Display/n697 ,open_n97224}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_0|u2_Display/lt31_cin  (
    .a({\u2_Display/n731 ,1'b0}),
    .b({1'b0,open_n97230}),
    .fco(\u2_Display/lt31_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_10|u2_Display/lt31_9  (
    .a({\u2_Display/n721 ,\u2_Display/n722 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c9 ),
    .fco(\u2_Display/lt31_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_12|u2_Display/lt31_11  (
    .a({\u2_Display/n719 ,\u2_Display/n720 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c11 ),
    .fco(\u2_Display/lt31_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_14|u2_Display/lt31_13  (
    .a({\u2_Display/n717 ,\u2_Display/n718 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c13 ),
    .fco(\u2_Display/lt31_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_16|u2_Display/lt31_15  (
    .a({\u2_Display/n715 ,\u2_Display/n716 }),
    .b(2'b10),
    .fci(\u2_Display/lt31_c15 ),
    .fco(\u2_Display/lt31_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_18|u2_Display/lt31_17  (
    .a({\u2_Display/n713 ,\u2_Display/n714 }),
    .b(2'b10),
    .fci(\u2_Display/lt31_c17 ),
    .fco(\u2_Display/lt31_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_20|u2_Display/lt31_19  (
    .a({\u2_Display/n711 ,\u2_Display/n712 }),
    .b(2'b11),
    .fci(\u2_Display/lt31_c19 ),
    .fco(\u2_Display/lt31_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_22|u2_Display/lt31_21  (
    .a({\u2_Display/n709 ,\u2_Display/n710 }),
    .b(2'b11),
    .fci(\u2_Display/lt31_c21 ),
    .fco(\u2_Display/lt31_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_24|u2_Display/lt31_23  (
    .a({\u2_Display/n707 ,\u2_Display/n708 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c23 ),
    .fco(\u2_Display/lt31_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_26|u2_Display/lt31_25  (
    .a({\u2_Display/n705 ,\u2_Display/n706 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c25 ),
    .fco(\u2_Display/lt31_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_28|u2_Display/lt31_27  (
    .a({\u2_Display/n703 ,\u2_Display/n704 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c27 ),
    .fco(\u2_Display/lt31_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_2|u2_Display/lt31_1  (
    .a({\u2_Display/n729 ,\u2_Display/n730 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c1 ),
    .fco(\u2_Display/lt31_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_30|u2_Display/lt31_29  (
    .a({\u2_Display/n701 ,\u2_Display/n702 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c29 ),
    .fco(\u2_Display/lt31_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_4|u2_Display/lt31_3  (
    .a({\u2_Display/n727 ,\u2_Display/n728 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c3 ),
    .fco(\u2_Display/lt31_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_6|u2_Display/lt31_5  (
    .a({\u2_Display/n725 ,\u2_Display/n726 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c5 ),
    .fco(\u2_Display/lt31_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_8|u2_Display/lt31_7  (
    .a({\u2_Display/n723 ,\u2_Display/n724 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c7 ),
    .fco(\u2_Display/lt31_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_cout|u2_Display/lt31_31  (
    .a({1'b0,\u2_Display/n700 }),
    .b(2'b10),
    .fci(\u2_Display/lt31_c31 ),
    .f({\u2_Display/n732 ,open_n97634}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_0|u2_Display/lt32_cin  (
    .a({\u2_Display/n766 ,1'b0}),
    .b({1'b0,open_n97640}),
    .fco(\u2_Display/lt32_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_10|u2_Display/lt32_9  (
    .a({\u2_Display/n756 ,\u2_Display/n757 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c9 ),
    .fco(\u2_Display/lt32_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_12|u2_Display/lt32_11  (
    .a({\u2_Display/n754 ,\u2_Display/n755 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c11 ),
    .fco(\u2_Display/lt32_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_14|u2_Display/lt32_13  (
    .a({\u2_Display/n752 ,\u2_Display/n753 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c13 ),
    .fco(\u2_Display/lt32_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_16|u2_Display/lt32_15  (
    .a({\u2_Display/n750 ,\u2_Display/n751 }),
    .b(2'b01),
    .fci(\u2_Display/lt32_c15 ),
    .fco(\u2_Display/lt32_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_18|u2_Display/lt32_17  (
    .a({\u2_Display/n748 ,\u2_Display/n749 }),
    .b(2'b11),
    .fci(\u2_Display/lt32_c17 ),
    .fco(\u2_Display/lt32_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_20|u2_Display/lt32_19  (
    .a({\u2_Display/n746 ,\u2_Display/n747 }),
    .b(2'b11),
    .fci(\u2_Display/lt32_c19 ),
    .fco(\u2_Display/lt32_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_22|u2_Display/lt32_21  (
    .a({\u2_Display/n744 ,\u2_Display/n745 }),
    .b(2'b01),
    .fci(\u2_Display/lt32_c21 ),
    .fco(\u2_Display/lt32_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_24|u2_Display/lt32_23  (
    .a({\u2_Display/n742 ,\u2_Display/n743 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c23 ),
    .fco(\u2_Display/lt32_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_26|u2_Display/lt32_25  (
    .a({\u2_Display/n740 ,\u2_Display/n741 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c25 ),
    .fco(\u2_Display/lt32_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_28|u2_Display/lt32_27  (
    .a({\u2_Display/n738 ,\u2_Display/n739 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c27 ),
    .fco(\u2_Display/lt32_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_2|u2_Display/lt32_1  (
    .a({\u2_Display/n764 ,\u2_Display/n765 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c1 ),
    .fco(\u2_Display/lt32_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_30|u2_Display/lt32_29  (
    .a({\u2_Display/n736 ,\u2_Display/n737 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c29 ),
    .fco(\u2_Display/lt32_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_4|u2_Display/lt32_3  (
    .a({\u2_Display/n762 ,\u2_Display/n763 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c3 ),
    .fco(\u2_Display/lt32_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_6|u2_Display/lt32_5  (
    .a({\u2_Display/n760 ,\u2_Display/n761 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c5 ),
    .fco(\u2_Display/lt32_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_8|u2_Display/lt32_7  (
    .a({\u2_Display/n758 ,\u2_Display/n759 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c7 ),
    .fco(\u2_Display/lt32_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_cout|u2_Display/lt32_31  (
    .a({1'b0,\u2_Display/n735 }),
    .b(2'b10),
    .fci(\u2_Display/lt32_c31 ),
    .f({\u2_Display/n767 ,open_n98044}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_0|u2_Display/lt33_cin  (
    .a({\u2_Display/n801 ,1'b0}),
    .b({1'b0,open_n98050}),
    .fco(\u2_Display/lt33_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_10|u2_Display/lt33_9  (
    .a({\u2_Display/n791 ,\u2_Display/n792 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c9 ),
    .fco(\u2_Display/lt33_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_12|u2_Display/lt33_11  (
    .a({\u2_Display/n789 ,\u2_Display/n790 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c11 ),
    .fco(\u2_Display/lt33_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_14|u2_Display/lt33_13  (
    .a({\u2_Display/n787 ,\u2_Display/n788 }),
    .b(2'b10),
    .fci(\u2_Display/lt33_c13 ),
    .fco(\u2_Display/lt33_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_16|u2_Display/lt33_15  (
    .a({\u2_Display/n785 ,\u2_Display/n786 }),
    .b(2'b10),
    .fci(\u2_Display/lt33_c15 ),
    .fco(\u2_Display/lt33_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_18|u2_Display/lt33_17  (
    .a({\u2_Display/n783 ,\u2_Display/n784 }),
    .b(2'b11),
    .fci(\u2_Display/lt33_c17 ),
    .fco(\u2_Display/lt33_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_20|u2_Display/lt33_19  (
    .a({\u2_Display/n781 ,\u2_Display/n782 }),
    .b(2'b11),
    .fci(\u2_Display/lt33_c19 ),
    .fco(\u2_Display/lt33_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_22|u2_Display/lt33_21  (
    .a({\u2_Display/n779 ,\u2_Display/n780 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c21 ),
    .fco(\u2_Display/lt33_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_24|u2_Display/lt33_23  (
    .a({\u2_Display/n777 ,\u2_Display/n778 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c23 ),
    .fco(\u2_Display/lt33_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_26|u2_Display/lt33_25  (
    .a({\u2_Display/n775 ,\u2_Display/n776 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c25 ),
    .fco(\u2_Display/lt33_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_28|u2_Display/lt33_27  (
    .a({\u2_Display/n773 ,\u2_Display/n774 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c27 ),
    .fco(\u2_Display/lt33_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_2|u2_Display/lt33_1  (
    .a({\u2_Display/n799 ,\u2_Display/n800 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c1 ),
    .fco(\u2_Display/lt33_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_30|u2_Display/lt33_29  (
    .a({\u2_Display/n771 ,\u2_Display/n772 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c29 ),
    .fco(\u2_Display/lt33_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_4|u2_Display/lt33_3  (
    .a({\u2_Display/n797 ,\u2_Display/n798 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c3 ),
    .fco(\u2_Display/lt33_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_6|u2_Display/lt33_5  (
    .a({\u2_Display/n795 ,\u2_Display/n796 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c5 ),
    .fco(\u2_Display/lt33_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_8|u2_Display/lt33_7  (
    .a({\u2_Display/n793 ,\u2_Display/n794 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c7 ),
    .fco(\u2_Display/lt33_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_cout|u2_Display/lt33_31  (
    .a({1'b0,\u2_Display/n770 }),
    .b(2'b10),
    .fci(\u2_Display/lt33_c31 ),
    .f({\u2_Display/n802 ,open_n98454}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_0|u2_Display/lt34_cin  (
    .a({\u2_Display/n836 ,1'b0}),
    .b({1'b0,open_n98460}),
    .fco(\u2_Display/lt34_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_10|u2_Display/lt34_9  (
    .a({\u2_Display/n826 ,\u2_Display/n827 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c9 ),
    .fco(\u2_Display/lt34_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_12|u2_Display/lt34_11  (
    .a({\u2_Display/n824 ,\u2_Display/n825 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c11 ),
    .fco(\u2_Display/lt34_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_14|u2_Display/lt34_13  (
    .a({\u2_Display/n822 ,\u2_Display/n823 }),
    .b(2'b01),
    .fci(\u2_Display/lt34_c13 ),
    .fco(\u2_Display/lt34_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_16|u2_Display/lt34_15  (
    .a({\u2_Display/n820 ,\u2_Display/n821 }),
    .b(2'b11),
    .fci(\u2_Display/lt34_c15 ),
    .fco(\u2_Display/lt34_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_18|u2_Display/lt34_17  (
    .a({\u2_Display/n818 ,\u2_Display/n819 }),
    .b(2'b11),
    .fci(\u2_Display/lt34_c17 ),
    .fco(\u2_Display/lt34_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_20|u2_Display/lt34_19  (
    .a({\u2_Display/n816 ,\u2_Display/n817 }),
    .b(2'b01),
    .fci(\u2_Display/lt34_c19 ),
    .fco(\u2_Display/lt34_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_22|u2_Display/lt34_21  (
    .a({\u2_Display/n814 ,\u2_Display/n815 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c21 ),
    .fco(\u2_Display/lt34_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_24|u2_Display/lt34_23  (
    .a({\u2_Display/n812 ,\u2_Display/n813 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c23 ),
    .fco(\u2_Display/lt34_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_26|u2_Display/lt34_25  (
    .a({\u2_Display/n810 ,\u2_Display/n811 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c25 ),
    .fco(\u2_Display/lt34_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_28|u2_Display/lt34_27  (
    .a({\u2_Display/n808 ,\u2_Display/n809 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c27 ),
    .fco(\u2_Display/lt34_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_2|u2_Display/lt34_1  (
    .a({\u2_Display/n834 ,\u2_Display/n835 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c1 ),
    .fco(\u2_Display/lt34_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_30|u2_Display/lt34_29  (
    .a({\u2_Display/n806 ,\u2_Display/n807 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c29 ),
    .fco(\u2_Display/lt34_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_4|u2_Display/lt34_3  (
    .a({\u2_Display/n832 ,\u2_Display/n833 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c3 ),
    .fco(\u2_Display/lt34_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_6|u2_Display/lt34_5  (
    .a({\u2_Display/n830 ,\u2_Display/n831 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c5 ),
    .fco(\u2_Display/lt34_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_8|u2_Display/lt34_7  (
    .a({\u2_Display/n828 ,\u2_Display/n829 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c7 ),
    .fco(\u2_Display/lt34_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_cout|u2_Display/lt34_31  (
    .a({1'b0,\u2_Display/n805 }),
    .b(2'b10),
    .fci(\u2_Display/lt34_c31 ),
    .f({\u2_Display/n837 ,open_n98864}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_0|u2_Display/lt35_cin  (
    .a({\u2_Display/n871 ,1'b0}),
    .b({1'b0,open_n98870}),
    .fco(\u2_Display/lt35_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_10|u2_Display/lt35_9  (
    .a({\u2_Display/n861 ,\u2_Display/n862 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c9 ),
    .fco(\u2_Display/lt35_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_12|u2_Display/lt35_11  (
    .a({\u2_Display/n859 ,\u2_Display/n860 }),
    .b(2'b10),
    .fci(\u2_Display/lt35_c11 ),
    .fco(\u2_Display/lt35_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_14|u2_Display/lt35_13  (
    .a({\u2_Display/n857 ,\u2_Display/n858 }),
    .b(2'b10),
    .fci(\u2_Display/lt35_c13 ),
    .fco(\u2_Display/lt35_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_16|u2_Display/lt35_15  (
    .a({\u2_Display/n855 ,\u2_Display/n856 }),
    .b(2'b11),
    .fci(\u2_Display/lt35_c15 ),
    .fco(\u2_Display/lt35_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_18|u2_Display/lt35_17  (
    .a({\u2_Display/n853 ,\u2_Display/n854 }),
    .b(2'b11),
    .fci(\u2_Display/lt35_c17 ),
    .fco(\u2_Display/lt35_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_20|u2_Display/lt35_19  (
    .a({\u2_Display/n851 ,\u2_Display/n852 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c19 ),
    .fco(\u2_Display/lt35_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_22|u2_Display/lt35_21  (
    .a({\u2_Display/n849 ,\u2_Display/n850 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c21 ),
    .fco(\u2_Display/lt35_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_24|u2_Display/lt35_23  (
    .a({\u2_Display/n847 ,\u2_Display/n848 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c23 ),
    .fco(\u2_Display/lt35_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_26|u2_Display/lt35_25  (
    .a({\u2_Display/n845 ,\u2_Display/n846 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c25 ),
    .fco(\u2_Display/lt35_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_28|u2_Display/lt35_27  (
    .a({\u2_Display/n843 ,\u2_Display/n844 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c27 ),
    .fco(\u2_Display/lt35_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_2|u2_Display/lt35_1  (
    .a({\u2_Display/n869 ,\u2_Display/n870 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c1 ),
    .fco(\u2_Display/lt35_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_30|u2_Display/lt35_29  (
    .a({\u2_Display/n841 ,\u2_Display/n842 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c29 ),
    .fco(\u2_Display/lt35_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_4|u2_Display/lt35_3  (
    .a({\u2_Display/n867 ,\u2_Display/n868 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c3 ),
    .fco(\u2_Display/lt35_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_6|u2_Display/lt35_5  (
    .a({\u2_Display/n865 ,\u2_Display/n866 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c5 ),
    .fco(\u2_Display/lt35_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_8|u2_Display/lt35_7  (
    .a({\u2_Display/n863 ,\u2_Display/n864 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c7 ),
    .fco(\u2_Display/lt35_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_cout|u2_Display/lt35_31  (
    .a({1'b0,\u2_Display/n840 }),
    .b(2'b10),
    .fci(\u2_Display/lt35_c31 ),
    .f({\u2_Display/n872 ,open_n99274}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_0|u2_Display/lt36_cin  (
    .a({\u2_Display/n906 ,1'b0}),
    .b({1'b0,open_n99280}),
    .fco(\u2_Display/lt36_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_10|u2_Display/lt36_9  (
    .a({\u2_Display/n896 ,\u2_Display/n897 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c9 ),
    .fco(\u2_Display/lt36_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_12|u2_Display/lt36_11  (
    .a({\u2_Display/n894 ,\u2_Display/n895 }),
    .b(2'b01),
    .fci(\u2_Display/lt36_c11 ),
    .fco(\u2_Display/lt36_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_14|u2_Display/lt36_13  (
    .a({\u2_Display/n892 ,\u2_Display/n893 }),
    .b(2'b11),
    .fci(\u2_Display/lt36_c13 ),
    .fco(\u2_Display/lt36_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_16|u2_Display/lt36_15  (
    .a({\u2_Display/n890 ,\u2_Display/n891 }),
    .b(2'b11),
    .fci(\u2_Display/lt36_c15 ),
    .fco(\u2_Display/lt36_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_18|u2_Display/lt36_17  (
    .a({\u2_Display/n888 ,\u2_Display/n889 }),
    .b(2'b01),
    .fci(\u2_Display/lt36_c17 ),
    .fco(\u2_Display/lt36_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_20|u2_Display/lt36_19  (
    .a({\u2_Display/n886 ,\u2_Display/n887 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c19 ),
    .fco(\u2_Display/lt36_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_22|u2_Display/lt36_21  (
    .a({\u2_Display/n884 ,\u2_Display/n885 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c21 ),
    .fco(\u2_Display/lt36_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_24|u2_Display/lt36_23  (
    .a({\u2_Display/n882 ,\u2_Display/n883 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c23 ),
    .fco(\u2_Display/lt36_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_26|u2_Display/lt36_25  (
    .a({\u2_Display/n880 ,\u2_Display/n881 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c25 ),
    .fco(\u2_Display/lt36_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_28|u2_Display/lt36_27  (
    .a({\u2_Display/n878 ,\u2_Display/n879 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c27 ),
    .fco(\u2_Display/lt36_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_2|u2_Display/lt36_1  (
    .a({\u2_Display/n904 ,\u2_Display/n905 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c1 ),
    .fco(\u2_Display/lt36_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_30|u2_Display/lt36_29  (
    .a({\u2_Display/n876 ,\u2_Display/n877 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c29 ),
    .fco(\u2_Display/lt36_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_4|u2_Display/lt36_3  (
    .a({\u2_Display/n902 ,\u2_Display/n903 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c3 ),
    .fco(\u2_Display/lt36_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_6|u2_Display/lt36_5  (
    .a({\u2_Display/n900 ,\u2_Display/n901 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c5 ),
    .fco(\u2_Display/lt36_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_8|u2_Display/lt36_7  (
    .a({\u2_Display/n898 ,\u2_Display/n899 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c7 ),
    .fco(\u2_Display/lt36_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_cout|u2_Display/lt36_31  (
    .a({1'b0,\u2_Display/n875 }),
    .b(2'b10),
    .fci(\u2_Display/lt36_c31 ),
    .f({\u2_Display/n907 ,open_n99684}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_0|u2_Display/lt37_cin  (
    .a({\u2_Display/n941 ,1'b0}),
    .b({1'b0,open_n99690}),
    .fco(\u2_Display/lt37_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_10|u2_Display/lt37_9  (
    .a({\u2_Display/n931 ,\u2_Display/n932 }),
    .b(2'b10),
    .fci(\u2_Display/lt37_c9 ),
    .fco(\u2_Display/lt37_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_12|u2_Display/lt37_11  (
    .a({\u2_Display/n929 ,\u2_Display/n930 }),
    .b(2'b10),
    .fci(\u2_Display/lt37_c11 ),
    .fco(\u2_Display/lt37_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_14|u2_Display/lt37_13  (
    .a({\u2_Display/n927 ,\u2_Display/n928 }),
    .b(2'b11),
    .fci(\u2_Display/lt37_c13 ),
    .fco(\u2_Display/lt37_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_16|u2_Display/lt37_15  (
    .a({\u2_Display/n925 ,\u2_Display/n926 }),
    .b(2'b11),
    .fci(\u2_Display/lt37_c15 ),
    .fco(\u2_Display/lt37_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_18|u2_Display/lt37_17  (
    .a({\u2_Display/n923 ,\u2_Display/n924 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c17 ),
    .fco(\u2_Display/lt37_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_20|u2_Display/lt37_19  (
    .a({\u2_Display/n921 ,\u2_Display/n922 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c19 ),
    .fco(\u2_Display/lt37_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_22|u2_Display/lt37_21  (
    .a({\u2_Display/n919 ,\u2_Display/n920 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c21 ),
    .fco(\u2_Display/lt37_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_24|u2_Display/lt37_23  (
    .a({\u2_Display/n917 ,\u2_Display/n918 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c23 ),
    .fco(\u2_Display/lt37_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_26|u2_Display/lt37_25  (
    .a({\u2_Display/n915 ,\u2_Display/n916 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c25 ),
    .fco(\u2_Display/lt37_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_28|u2_Display/lt37_27  (
    .a({\u2_Display/n913 ,\u2_Display/n914 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c27 ),
    .fco(\u2_Display/lt37_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_2|u2_Display/lt37_1  (
    .a({\u2_Display/n939 ,\u2_Display/n940 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c1 ),
    .fco(\u2_Display/lt37_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_30|u2_Display/lt37_29  (
    .a({\u2_Display/n911 ,\u2_Display/n912 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c29 ),
    .fco(\u2_Display/lt37_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_4|u2_Display/lt37_3  (
    .a({\u2_Display/n937 ,\u2_Display/n938 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c3 ),
    .fco(\u2_Display/lt37_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_6|u2_Display/lt37_5  (
    .a({\u2_Display/n935 ,\u2_Display/n936 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c5 ),
    .fco(\u2_Display/lt37_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_8|u2_Display/lt37_7  (
    .a({\u2_Display/n933 ,\u2_Display/n934 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c7 ),
    .fco(\u2_Display/lt37_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_cout|u2_Display/lt37_31  (
    .a({1'b0,\u2_Display/n910 }),
    .b(2'b10),
    .fci(\u2_Display/lt37_c31 ),
    .f({\u2_Display/n942 ,open_n100094}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_0|u2_Display/lt38_cin  (
    .a({\u2_Display/n976 ,1'b0}),
    .b({1'b0,open_n100100}),
    .fco(\u2_Display/lt38_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_10|u2_Display/lt38_9  (
    .a({\u2_Display/n966 ,\u2_Display/n967 }),
    .b(2'b01),
    .fci(\u2_Display/lt38_c9 ),
    .fco(\u2_Display/lt38_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_12|u2_Display/lt38_11  (
    .a({\u2_Display/n964 ,\u2_Display/n965 }),
    .b(2'b11),
    .fci(\u2_Display/lt38_c11 ),
    .fco(\u2_Display/lt38_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_14|u2_Display/lt38_13  (
    .a({\u2_Display/n962 ,\u2_Display/n963 }),
    .b(2'b11),
    .fci(\u2_Display/lt38_c13 ),
    .fco(\u2_Display/lt38_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_16|u2_Display/lt38_15  (
    .a({\u2_Display/n960 ,\u2_Display/n961 }),
    .b(2'b01),
    .fci(\u2_Display/lt38_c15 ),
    .fco(\u2_Display/lt38_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_18|u2_Display/lt38_17  (
    .a({\u2_Display/n958 ,\u2_Display/n959 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c17 ),
    .fco(\u2_Display/lt38_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_20|u2_Display/lt38_19  (
    .a({\u2_Display/n956 ,\u2_Display/n957 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c19 ),
    .fco(\u2_Display/lt38_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_22|u2_Display/lt38_21  (
    .a({\u2_Display/n954 ,\u2_Display/n955 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c21 ),
    .fco(\u2_Display/lt38_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_24|u2_Display/lt38_23  (
    .a({\u2_Display/n952 ,\u2_Display/n953 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c23 ),
    .fco(\u2_Display/lt38_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_26|u2_Display/lt38_25  (
    .a({\u2_Display/n950 ,\u2_Display/n951 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c25 ),
    .fco(\u2_Display/lt38_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_28|u2_Display/lt38_27  (
    .a({\u2_Display/n948 ,\u2_Display/n949 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c27 ),
    .fco(\u2_Display/lt38_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_2|u2_Display/lt38_1  (
    .a({\u2_Display/n974 ,\u2_Display/n975 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c1 ),
    .fco(\u2_Display/lt38_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_30|u2_Display/lt38_29  (
    .a({\u2_Display/n946 ,\u2_Display/n947 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c29 ),
    .fco(\u2_Display/lt38_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_4|u2_Display/lt38_3  (
    .a({\u2_Display/n972 ,\u2_Display/n973 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c3 ),
    .fco(\u2_Display/lt38_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_6|u2_Display/lt38_5  (
    .a({\u2_Display/n970 ,\u2_Display/n971 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c5 ),
    .fco(\u2_Display/lt38_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_8|u2_Display/lt38_7  (
    .a({\u2_Display/n968 ,\u2_Display/n969 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c7 ),
    .fco(\u2_Display/lt38_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_cout|u2_Display/lt38_31  (
    .a({1'b0,\u2_Display/n945 }),
    .b(2'b10),
    .fci(\u2_Display/lt38_c31 ),
    .f({\u2_Display/n977 ,open_n100504}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_0|u2_Display/lt39_cin  (
    .a({\u2_Display/n1011 ,1'b0}),
    .b({1'b0,open_n100510}),
    .fco(\u2_Display/lt39_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_10|u2_Display/lt39_9  (
    .a({\u2_Display/n1001 ,\u2_Display/n1002 }),
    .b(2'b10),
    .fci(\u2_Display/lt39_c9 ),
    .fco(\u2_Display/lt39_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_12|u2_Display/lt39_11  (
    .a({\u2_Display/n999 ,\u2_Display/n1000 }),
    .b(2'b11),
    .fci(\u2_Display/lt39_c11 ),
    .fco(\u2_Display/lt39_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_14|u2_Display/lt39_13  (
    .a({\u2_Display/n997 ,\u2_Display/n998 }),
    .b(2'b11),
    .fci(\u2_Display/lt39_c13 ),
    .fco(\u2_Display/lt39_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_16|u2_Display/lt39_15  (
    .a({\u2_Display/n995 ,\u2_Display/n996 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c15 ),
    .fco(\u2_Display/lt39_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_18|u2_Display/lt39_17  (
    .a({\u2_Display/n993 ,\u2_Display/n994 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c17 ),
    .fco(\u2_Display/lt39_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_20|u2_Display/lt39_19  (
    .a({\u2_Display/n991 ,\u2_Display/n992 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c19 ),
    .fco(\u2_Display/lt39_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_22|u2_Display/lt39_21  (
    .a({\u2_Display/n989 ,\u2_Display/n990 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c21 ),
    .fco(\u2_Display/lt39_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_24|u2_Display/lt39_23  (
    .a({\u2_Display/n987 ,\u2_Display/n988 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c23 ),
    .fco(\u2_Display/lt39_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_26|u2_Display/lt39_25  (
    .a({\u2_Display/n985 ,\u2_Display/n986 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c25 ),
    .fco(\u2_Display/lt39_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_28|u2_Display/lt39_27  (
    .a({\u2_Display/n983 ,\u2_Display/n984 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c27 ),
    .fco(\u2_Display/lt39_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_2|u2_Display/lt39_1  (
    .a({\u2_Display/n1009 ,\u2_Display/n1010 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c1 ),
    .fco(\u2_Display/lt39_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_30|u2_Display/lt39_29  (
    .a({\u2_Display/n981 ,\u2_Display/n982 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c29 ),
    .fco(\u2_Display/lt39_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_4|u2_Display/lt39_3  (
    .a({\u2_Display/n1007 ,\u2_Display/n1008 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c3 ),
    .fco(\u2_Display/lt39_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_6|u2_Display/lt39_5  (
    .a({\u2_Display/n1005 ,\u2_Display/n1006 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c5 ),
    .fco(\u2_Display/lt39_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_8|u2_Display/lt39_7  (
    .a({\u2_Display/n1003 ,\u2_Display/n1004 }),
    .b(2'b10),
    .fci(\u2_Display/lt39_c7 ),
    .fco(\u2_Display/lt39_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_cout|u2_Display/lt39_31  (
    .a({1'b0,\u2_Display/n980 }),
    .b(2'b10),
    .fci(\u2_Display/lt39_c31 ),
    .f({\u2_Display/n1012 ,open_n100914}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_0|u2_Display/lt3_cin  (
    .a({\u2_Display/j [0],1'b0}),
    .b({lcd_ypos[0],open_n100920}),
    .fco(\u2_Display/lt3_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_10|u2_Display/lt3_9  (
    .a({1'b0,\u2_Display/j [9]}),
    .b(lcd_ypos[10:9]),
    .fci(\u2_Display/lt3_c9 ),
    .fco(\u2_Display/lt3_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_2|u2_Display/lt3_1  (
    .a(\u2_Display/j [2:1]),
    .b(lcd_ypos[2:1]),
    .fci(\u2_Display/lt3_c1 ),
    .fco(\u2_Display/lt3_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_4|u2_Display/lt3_3  (
    .a(\u2_Display/j [4:3]),
    .b(lcd_ypos[4:3]),
    .fci(\u2_Display/lt3_c3 ),
    .fco(\u2_Display/lt3_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_6|u2_Display/lt3_5  (
    .a(\u2_Display/j [6:5]),
    .b(lcd_ypos[6:5]),
    .fci(\u2_Display/lt3_c5 ),
    .fco(\u2_Display/lt3_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_8|u2_Display/lt3_7  (
    .a(\u2_Display/j [8:7]),
    .b(lcd_ypos[8:7]),
    .fci(\u2_Display/lt3_c7 ),
    .fco(\u2_Display/lt3_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_cout|u2_Display/lt3_11  (
    .a(2'b00),
    .b({1'b1,lcd_ypos[11]}),
    .fci(\u2_Display/lt3_c11 ),
    .f({\u2_Display/n50 ,open_n101084}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_0|u2_Display/lt40_cin  (
    .a({\u2_Display/n1046 ,1'b0}),
    .b({1'b0,open_n101090}),
    .fco(\u2_Display/lt40_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_10|u2_Display/lt40_9  (
    .a({\u2_Display/n1036 ,\u2_Display/n1037 }),
    .b(2'b11),
    .fci(\u2_Display/lt40_c9 ),
    .fco(\u2_Display/lt40_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_12|u2_Display/lt40_11  (
    .a({\u2_Display/n1034 ,\u2_Display/n1035 }),
    .b(2'b11),
    .fci(\u2_Display/lt40_c11 ),
    .fco(\u2_Display/lt40_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_14|u2_Display/lt40_13  (
    .a({\u2_Display/n1032 ,\u2_Display/n1033 }),
    .b(2'b01),
    .fci(\u2_Display/lt40_c13 ),
    .fco(\u2_Display/lt40_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_16|u2_Display/lt40_15  (
    .a({\u2_Display/n1030 ,\u2_Display/n1031 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c15 ),
    .fco(\u2_Display/lt40_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_18|u2_Display/lt40_17  (
    .a({\u2_Display/n1028 ,\u2_Display/n1029 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c17 ),
    .fco(\u2_Display/lt40_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_20|u2_Display/lt40_19  (
    .a({\u2_Display/n1026 ,\u2_Display/n1027 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c19 ),
    .fco(\u2_Display/lt40_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_22|u2_Display/lt40_21  (
    .a({\u2_Display/n1024 ,\u2_Display/n1025 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c21 ),
    .fco(\u2_Display/lt40_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_24|u2_Display/lt40_23  (
    .a({\u2_Display/n1022 ,\u2_Display/n1023 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c23 ),
    .fco(\u2_Display/lt40_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_26|u2_Display/lt40_25  (
    .a({\u2_Display/n1020 ,\u2_Display/n1021 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c25 ),
    .fco(\u2_Display/lt40_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_28|u2_Display/lt40_27  (
    .a({\u2_Display/n1018 ,\u2_Display/n1019 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c27 ),
    .fco(\u2_Display/lt40_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_2|u2_Display/lt40_1  (
    .a({\u2_Display/n1044 ,\u2_Display/n1045 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c1 ),
    .fco(\u2_Display/lt40_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_30|u2_Display/lt40_29  (
    .a({\u2_Display/n1016 ,\u2_Display/n1017 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c29 ),
    .fco(\u2_Display/lt40_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_4|u2_Display/lt40_3  (
    .a({\u2_Display/n1042 ,\u2_Display/n1043 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c3 ),
    .fco(\u2_Display/lt40_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_6|u2_Display/lt40_5  (
    .a({\u2_Display/n1040 ,\u2_Display/n1041 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c5 ),
    .fco(\u2_Display/lt40_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_8|u2_Display/lt40_7  (
    .a({\u2_Display/n1038 ,\u2_Display/n1039 }),
    .b(2'b01),
    .fci(\u2_Display/lt40_c7 ),
    .fco(\u2_Display/lt40_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_cout|u2_Display/lt40_31  (
    .a({1'b0,\u2_Display/n1015 }),
    .b(2'b10),
    .fci(\u2_Display/lt40_c31 ),
    .f({\u2_Display/n1047 ,open_n101494}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_0|u2_Display/lt41_cin  (
    .a({\u2_Display/n1081 ,1'b0}),
    .b({1'b0,open_n101500}),
    .fco(\u2_Display/lt41_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_10|u2_Display/lt41_9  (
    .a({\u2_Display/n1071 ,\u2_Display/n1072 }),
    .b(2'b11),
    .fci(\u2_Display/lt41_c9 ),
    .fco(\u2_Display/lt41_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_12|u2_Display/lt41_11  (
    .a({\u2_Display/n1069 ,\u2_Display/n1070 }),
    .b(2'b11),
    .fci(\u2_Display/lt41_c11 ),
    .fco(\u2_Display/lt41_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_14|u2_Display/lt41_13  (
    .a({\u2_Display/n1067 ,\u2_Display/n1068 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c13 ),
    .fco(\u2_Display/lt41_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_16|u2_Display/lt41_15  (
    .a({\u2_Display/n1065 ,\u2_Display/n1066 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c15 ),
    .fco(\u2_Display/lt41_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_18|u2_Display/lt41_17  (
    .a({\u2_Display/n1063 ,\u2_Display/n1064 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c17 ),
    .fco(\u2_Display/lt41_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_20|u2_Display/lt41_19  (
    .a({\u2_Display/n1061 ,\u2_Display/n1062 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c19 ),
    .fco(\u2_Display/lt41_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_22|u2_Display/lt41_21  (
    .a({\u2_Display/n1059 ,\u2_Display/n1060 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c21 ),
    .fco(\u2_Display/lt41_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_24|u2_Display/lt41_23  (
    .a({\u2_Display/n1057 ,\u2_Display/n1058 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c23 ),
    .fco(\u2_Display/lt41_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_26|u2_Display/lt41_25  (
    .a({\u2_Display/n1055 ,\u2_Display/n1056 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c25 ),
    .fco(\u2_Display/lt41_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_28|u2_Display/lt41_27  (
    .a({\u2_Display/n1053 ,\u2_Display/n1054 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c27 ),
    .fco(\u2_Display/lt41_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_2|u2_Display/lt41_1  (
    .a({\u2_Display/n1079 ,\u2_Display/n1080 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c1 ),
    .fco(\u2_Display/lt41_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_30|u2_Display/lt41_29  (
    .a({\u2_Display/n1051 ,\u2_Display/n1052 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c29 ),
    .fco(\u2_Display/lt41_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_4|u2_Display/lt41_3  (
    .a({\u2_Display/n1077 ,\u2_Display/n1078 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c3 ),
    .fco(\u2_Display/lt41_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_6|u2_Display/lt41_5  (
    .a({\u2_Display/n1075 ,\u2_Display/n1076 }),
    .b(2'b10),
    .fci(\u2_Display/lt41_c5 ),
    .fco(\u2_Display/lt41_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_8|u2_Display/lt41_7  (
    .a({\u2_Display/n1073 ,\u2_Display/n1074 }),
    .b(2'b10),
    .fci(\u2_Display/lt41_c7 ),
    .fco(\u2_Display/lt41_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_cout|u2_Display/lt41_31  (
    .a({1'b0,\u2_Display/n1050 }),
    .b(2'b10),
    .fci(\u2_Display/lt41_c31 ),
    .f({\u2_Display/n1082 ,open_n101904}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_0|u2_Display/lt42_cin  (
    .a({\u2_Display/n1116 ,1'b0}),
    .b({1'b0,open_n101910}),
    .fco(\u2_Display/lt42_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_10|u2_Display/lt42_9  (
    .a({\u2_Display/n1106 ,\u2_Display/n1107 }),
    .b(2'b11),
    .fci(\u2_Display/lt42_c9 ),
    .fco(\u2_Display/lt42_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_12|u2_Display/lt42_11  (
    .a({\u2_Display/n1104 ,\u2_Display/n1105 }),
    .b(2'b01),
    .fci(\u2_Display/lt42_c11 ),
    .fco(\u2_Display/lt42_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_14|u2_Display/lt42_13  (
    .a({\u2_Display/n1102 ,\u2_Display/n1103 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c13 ),
    .fco(\u2_Display/lt42_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_16|u2_Display/lt42_15  (
    .a({\u2_Display/n1100 ,\u2_Display/n1101 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c15 ),
    .fco(\u2_Display/lt42_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_18|u2_Display/lt42_17  (
    .a({\u2_Display/n1098 ,\u2_Display/n1099 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c17 ),
    .fco(\u2_Display/lt42_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_20|u2_Display/lt42_19  (
    .a({\u2_Display/n1096 ,\u2_Display/n1097 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c19 ),
    .fco(\u2_Display/lt42_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_22|u2_Display/lt42_21  (
    .a({\u2_Display/n1094 ,\u2_Display/n1095 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c21 ),
    .fco(\u2_Display/lt42_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_24|u2_Display/lt42_23  (
    .a({\u2_Display/n1092 ,\u2_Display/n1093 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c23 ),
    .fco(\u2_Display/lt42_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_26|u2_Display/lt42_25  (
    .a({\u2_Display/n1090 ,\u2_Display/n1091 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c25 ),
    .fco(\u2_Display/lt42_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_28|u2_Display/lt42_27  (
    .a({\u2_Display/n1088 ,\u2_Display/n1089 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c27 ),
    .fco(\u2_Display/lt42_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_2|u2_Display/lt42_1  (
    .a({\u2_Display/n1114 ,\u2_Display/n1115 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c1 ),
    .fco(\u2_Display/lt42_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_30|u2_Display/lt42_29  (
    .a({\u2_Display/n1086 ,\u2_Display/n1087 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c29 ),
    .fco(\u2_Display/lt42_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_4|u2_Display/lt42_3  (
    .a({\u2_Display/n1112 ,\u2_Display/n1113 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c3 ),
    .fco(\u2_Display/lt42_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_6|u2_Display/lt42_5  (
    .a({\u2_Display/n1110 ,\u2_Display/n1111 }),
    .b(2'b01),
    .fci(\u2_Display/lt42_c5 ),
    .fco(\u2_Display/lt42_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_8|u2_Display/lt42_7  (
    .a({\u2_Display/n1108 ,\u2_Display/n1109 }),
    .b(2'b11),
    .fci(\u2_Display/lt42_c7 ),
    .fco(\u2_Display/lt42_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_cout|u2_Display/lt42_31  (
    .a({1'b0,\u2_Display/n1085 }),
    .b(2'b10),
    .fci(\u2_Display/lt42_c31 ),
    .f({\u2_Display/n1117 ,open_n102314}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_0|u2_Display/lt43_cin  (
    .a({\u2_Display/n1151 ,1'b0}),
    .b({1'b0,open_n102320}),
    .fco(\u2_Display/lt43_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_10|u2_Display/lt43_9  (
    .a({\u2_Display/n1141 ,\u2_Display/n1142 }),
    .b(2'b11),
    .fci(\u2_Display/lt43_c9 ),
    .fco(\u2_Display/lt43_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_12|u2_Display/lt43_11  (
    .a({\u2_Display/n1139 ,\u2_Display/n1140 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c11 ),
    .fco(\u2_Display/lt43_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_14|u2_Display/lt43_13  (
    .a({\u2_Display/n1137 ,\u2_Display/n1138 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c13 ),
    .fco(\u2_Display/lt43_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_16|u2_Display/lt43_15  (
    .a({\u2_Display/n1135 ,\u2_Display/n1136 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c15 ),
    .fco(\u2_Display/lt43_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_18|u2_Display/lt43_17  (
    .a({\u2_Display/n1133 ,\u2_Display/n1134 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c17 ),
    .fco(\u2_Display/lt43_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_20|u2_Display/lt43_19  (
    .a({\u2_Display/n1131 ,\u2_Display/n1132 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c19 ),
    .fco(\u2_Display/lt43_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_22|u2_Display/lt43_21  (
    .a({\u2_Display/n1129 ,\u2_Display/n1130 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c21 ),
    .fco(\u2_Display/lt43_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_24|u2_Display/lt43_23  (
    .a({\u2_Display/n1127 ,\u2_Display/n1128 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c23 ),
    .fco(\u2_Display/lt43_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_26|u2_Display/lt43_25  (
    .a({\u2_Display/n1125 ,\u2_Display/n1126 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c25 ),
    .fco(\u2_Display/lt43_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_28|u2_Display/lt43_27  (
    .a({\u2_Display/n1123 ,\u2_Display/n1124 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c27 ),
    .fco(\u2_Display/lt43_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_2|u2_Display/lt43_1  (
    .a({\u2_Display/n1149 ,\u2_Display/n1150 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c1 ),
    .fco(\u2_Display/lt43_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_30|u2_Display/lt43_29  (
    .a({\u2_Display/n1121 ,\u2_Display/n1122 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c29 ),
    .fco(\u2_Display/lt43_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_4|u2_Display/lt43_3  (
    .a({\u2_Display/n1147 ,\u2_Display/n1148 }),
    .b(2'b10),
    .fci(\u2_Display/lt43_c3 ),
    .fco(\u2_Display/lt43_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_6|u2_Display/lt43_5  (
    .a({\u2_Display/n1145 ,\u2_Display/n1146 }),
    .b(2'b10),
    .fci(\u2_Display/lt43_c5 ),
    .fco(\u2_Display/lt43_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_8|u2_Display/lt43_7  (
    .a({\u2_Display/n1143 ,\u2_Display/n1144 }),
    .b(2'b11),
    .fci(\u2_Display/lt43_c7 ),
    .fco(\u2_Display/lt43_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_cout|u2_Display/lt43_31  (
    .a({1'b0,\u2_Display/n1120 }),
    .b(2'b10),
    .fci(\u2_Display/lt43_c31 ),
    .f({\u2_Display/n1152 ,open_n102724}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_0|u2_Display/lt44_cin  (
    .a({\u2_Display/n1186 ,1'b0}),
    .b({1'b0,open_n102730}),
    .fco(\u2_Display/lt44_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_10|u2_Display/lt44_9  (
    .a({\u2_Display/n1176 ,\u2_Display/n1177 }),
    .b(2'b01),
    .fci(\u2_Display/lt44_c9 ),
    .fco(\u2_Display/lt44_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_12|u2_Display/lt44_11  (
    .a({\u2_Display/n1174 ,\u2_Display/n1175 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c11 ),
    .fco(\u2_Display/lt44_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_14|u2_Display/lt44_13  (
    .a({\u2_Display/n1172 ,\u2_Display/n1173 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c13 ),
    .fco(\u2_Display/lt44_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_16|u2_Display/lt44_15  (
    .a({\u2_Display/n1170 ,\u2_Display/n1171 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c15 ),
    .fco(\u2_Display/lt44_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_18|u2_Display/lt44_17  (
    .a({\u2_Display/n1168 ,\u2_Display/n1169 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c17 ),
    .fco(\u2_Display/lt44_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_20|u2_Display/lt44_19  (
    .a({\u2_Display/n1166 ,\u2_Display/n1167 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c19 ),
    .fco(\u2_Display/lt44_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_22|u2_Display/lt44_21  (
    .a({\u2_Display/n1164 ,\u2_Display/n1165 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c21 ),
    .fco(\u2_Display/lt44_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_24|u2_Display/lt44_23  (
    .a({\u2_Display/n1162 ,\u2_Display/n1163 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c23 ),
    .fco(\u2_Display/lt44_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_26|u2_Display/lt44_25  (
    .a({\u2_Display/n1160 ,\u2_Display/n1161 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c25 ),
    .fco(\u2_Display/lt44_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_28|u2_Display/lt44_27  (
    .a({\u2_Display/n1158 ,\u2_Display/n1159 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c27 ),
    .fco(\u2_Display/lt44_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_2|u2_Display/lt44_1  (
    .a({\u2_Display/n1184 ,\u2_Display/n1185 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c1 ),
    .fco(\u2_Display/lt44_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_30|u2_Display/lt44_29  (
    .a({\u2_Display/n1156 ,\u2_Display/n1157 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c29 ),
    .fco(\u2_Display/lt44_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_4|u2_Display/lt44_3  (
    .a({\u2_Display/n1182 ,\u2_Display/n1183 }),
    .b(2'b01),
    .fci(\u2_Display/lt44_c3 ),
    .fco(\u2_Display/lt44_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_6|u2_Display/lt44_5  (
    .a({\u2_Display/n1180 ,\u2_Display/n1181 }),
    .b(2'b11),
    .fci(\u2_Display/lt44_c5 ),
    .fco(\u2_Display/lt44_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_8|u2_Display/lt44_7  (
    .a({\u2_Display/n1178 ,\u2_Display/n1179 }),
    .b(2'b11),
    .fci(\u2_Display/lt44_c7 ),
    .fco(\u2_Display/lt44_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_cout|u2_Display/lt44_31  (
    .a({1'b0,\u2_Display/n1155 }),
    .b(2'b10),
    .fci(\u2_Display/lt44_c31 ),
    .f({\u2_Display/n1187 ,open_n103134}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_0|u2_Display/lt4_2_cin  (
    .a({lcd_xpos[0],1'b0}),
    .b({\u2_Display/i [0],open_n103140}),
    .fco(\u2_Display/lt4_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_10|u2_Display/lt4_2_9  (
    .a(lcd_xpos[10:9]),
    .b(\u2_Display/n94 [3:2]),
    .fci(\u2_Display/lt4_2_c9 ),
    .fco(\u2_Display/lt4_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_2|u2_Display/lt4_2_1  (
    .a(lcd_xpos[2:1]),
    .b(\u2_Display/i [2:1]),
    .fci(\u2_Display/lt4_2_c1 ),
    .fco(\u2_Display/lt4_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_4|u2_Display/lt4_2_3  (
    .a(lcd_xpos[4:3]),
    .b(\u2_Display/i [4:3]),
    .fci(\u2_Display/lt4_2_c3 ),
    .fco(\u2_Display/lt4_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_6|u2_Display/lt4_2_5  (
    .a(lcd_xpos[6:5]),
    .b(\u2_Display/i [6:5]),
    .fci(\u2_Display/lt4_2_c5 ),
    .fco(\u2_Display/lt4_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_8|u2_Display/lt4_2_7  (
    .a(lcd_xpos[8:7]),
    .b(\u2_Display/n94 [1:0]),
    .fci(\u2_Display/lt4_2_c7 ),
    .fco(\u2_Display/lt4_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_cout|u2_Display/lt4_2_11  (
    .a({1'b0,lcd_xpos[11]}),
    .b({1'b1,\u2_Display/add4_2_co }),
    .fci(\u2_Display/lt4_2_c11 ),
    .f({\u2_Display/n95 ,open_n103304}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_0|u2_Display/lt55_cin  (
    .a({\u2_Display/counta [0],1'b0}),
    .b({1'b0,open_n103310}),
    .fco(\u2_Display/lt55_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_10|u2_Display/lt55_9  (
    .a(\u2_Display/counta [10:9]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c9 ),
    .fco(\u2_Display/lt55_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_12|u2_Display/lt55_11  (
    .a(\u2_Display/counta [12:11]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c11 ),
    .fco(\u2_Display/lt55_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_14|u2_Display/lt55_13  (
    .a(\u2_Display/counta [14:13]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c13 ),
    .fco(\u2_Display/lt55_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_16|u2_Display/lt55_15  (
    .a(\u2_Display/counta [16:15]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c15 ),
    .fco(\u2_Display/lt55_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_18|u2_Display/lt55_17  (
    .a(\u2_Display/counta [18:17]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c17 ),
    .fco(\u2_Display/lt55_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_20|u2_Display/lt55_19  (
    .a(\u2_Display/counta [20:19]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c19 ),
    .fco(\u2_Display/lt55_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_22|u2_Display/lt55_21  (
    .a(\u2_Display/counta [22:21]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c21 ),
    .fco(\u2_Display/lt55_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_24|u2_Display/lt55_23  (
    .a(\u2_Display/counta [24:23]),
    .b(2'b10),
    .fci(\u2_Display/lt55_c23 ),
    .fco(\u2_Display/lt55_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_26|u2_Display/lt55_25  (
    .a(\u2_Display/counta [26:25]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c25 ),
    .fco(\u2_Display/lt55_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_28|u2_Display/lt55_27  (
    .a(\u2_Display/counta [28:27]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c27 ),
    .fco(\u2_Display/lt55_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_2|u2_Display/lt55_1  (
    .a(\u2_Display/counta [2:1]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c1 ),
    .fco(\u2_Display/lt55_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_30|u2_Display/lt55_29  (
    .a(\u2_Display/counta [30:29]),
    .b(2'b11),
    .fci(\u2_Display/lt55_c29 ),
    .fco(\u2_Display/lt55_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_4|u2_Display/lt55_3  (
    .a(\u2_Display/counta [4:3]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c3 ),
    .fco(\u2_Display/lt55_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_6|u2_Display/lt55_5  (
    .a(\u2_Display/counta [6:5]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c5 ),
    .fco(\u2_Display/lt55_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_8|u2_Display/lt55_7  (
    .a(\u2_Display/counta [8:7]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c7 ),
    .fco(\u2_Display/lt55_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_cout|u2_Display/lt55_31  (
    .a({1'b0,\u2_Display/counta [31]}),
    .b(2'b11),
    .fci(\u2_Display/lt55_c31 ),
    .f({\u2_Display/n1540 ,open_n103714}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_0|u2_Display/lt56_cin  (
    .a({\u2_Display/n1574 ,1'b0}),
    .b({1'b0,open_n103720}),
    .fco(\u2_Display/lt56_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_10|u2_Display/lt56_9  (
    .a({\u2_Display/n1564 ,\u2_Display/n1565 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c9 ),
    .fco(\u2_Display/lt56_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_12|u2_Display/lt56_11  (
    .a({\u2_Display/n1562 ,\u2_Display/n1563 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c11 ),
    .fco(\u2_Display/lt56_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_14|u2_Display/lt56_13  (
    .a({\u2_Display/n1560 ,\u2_Display/n1561 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c13 ),
    .fco(\u2_Display/lt56_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_16|u2_Display/lt56_15  (
    .a({\u2_Display/n1558 ,\u2_Display/n1559 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c15 ),
    .fco(\u2_Display/lt56_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_18|u2_Display/lt56_17  (
    .a({\u2_Display/n1556 ,\u2_Display/n1557 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c17 ),
    .fco(\u2_Display/lt56_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_20|u2_Display/lt56_19  (
    .a({\u2_Display/n1554 ,\u2_Display/n1555 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c19 ),
    .fco(\u2_Display/lt56_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_22|u2_Display/lt56_21  (
    .a({\u2_Display/n1552 ,\u2_Display/n1553 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c21 ),
    .fco(\u2_Display/lt56_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_24|u2_Display/lt56_23  (
    .a({\u2_Display/n1550 ,\u2_Display/n1551 }),
    .b(2'b01),
    .fci(\u2_Display/lt56_c23 ),
    .fco(\u2_Display/lt56_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_26|u2_Display/lt56_25  (
    .a({\u2_Display/n1548 ,\u2_Display/n1549 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c25 ),
    .fco(\u2_Display/lt56_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_28|u2_Display/lt56_27  (
    .a({\u2_Display/n1546 ,\u2_Display/n1547 }),
    .b(2'b10),
    .fci(\u2_Display/lt56_c27 ),
    .fco(\u2_Display/lt56_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_2|u2_Display/lt56_1  (
    .a({\u2_Display/n1572 ,\u2_Display/n1573 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c1 ),
    .fco(\u2_Display/lt56_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_30|u2_Display/lt56_29  (
    .a({\u2_Display/n1544 ,\u2_Display/n1545 }),
    .b(2'b11),
    .fci(\u2_Display/lt56_c29 ),
    .fco(\u2_Display/lt56_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_4|u2_Display/lt56_3  (
    .a({\u2_Display/n1570 ,\u2_Display/n1571 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c3 ),
    .fco(\u2_Display/lt56_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_6|u2_Display/lt56_5  (
    .a({\u2_Display/n1568 ,\u2_Display/n1569 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c5 ),
    .fco(\u2_Display/lt56_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_8|u2_Display/lt56_7  (
    .a({\u2_Display/n1566 ,\u2_Display/n1567 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c7 ),
    .fco(\u2_Display/lt56_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_cout|u2_Display/lt56_31  (
    .a({1'b0,\u2_Display/n1543 }),
    .b(2'b10),
    .fci(\u2_Display/lt56_c31 ),
    .f({\u2_Display/n1575 ,open_n104124}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_0|u2_Display/lt57_cin  (
    .a({\u2_Display/n1609 ,1'b0}),
    .b({1'b0,open_n104130}),
    .fco(\u2_Display/lt57_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_10|u2_Display/lt57_9  (
    .a({\u2_Display/n1599 ,\u2_Display/n1600 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c9 ),
    .fco(\u2_Display/lt57_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_12|u2_Display/lt57_11  (
    .a({\u2_Display/n1597 ,\u2_Display/n1598 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c11 ),
    .fco(\u2_Display/lt57_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_14|u2_Display/lt57_13  (
    .a({\u2_Display/n1595 ,\u2_Display/n1596 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c13 ),
    .fco(\u2_Display/lt57_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_16|u2_Display/lt57_15  (
    .a({\u2_Display/n1593 ,\u2_Display/n1594 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c15 ),
    .fco(\u2_Display/lt57_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_18|u2_Display/lt57_17  (
    .a({\u2_Display/n1591 ,\u2_Display/n1592 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c17 ),
    .fco(\u2_Display/lt57_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_20|u2_Display/lt57_19  (
    .a({\u2_Display/n1589 ,\u2_Display/n1590 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c19 ),
    .fco(\u2_Display/lt57_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_22|u2_Display/lt57_21  (
    .a({\u2_Display/n1587 ,\u2_Display/n1588 }),
    .b(2'b10),
    .fci(\u2_Display/lt57_c21 ),
    .fco(\u2_Display/lt57_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_24|u2_Display/lt57_23  (
    .a({\u2_Display/n1585 ,\u2_Display/n1586 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c23 ),
    .fco(\u2_Display/lt57_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_26|u2_Display/lt57_25  (
    .a({\u2_Display/n1583 ,\u2_Display/n1584 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c25 ),
    .fco(\u2_Display/lt57_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_28|u2_Display/lt57_27  (
    .a({\u2_Display/n1581 ,\u2_Display/n1582 }),
    .b(2'b11),
    .fci(\u2_Display/lt57_c27 ),
    .fco(\u2_Display/lt57_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_2|u2_Display/lt57_1  (
    .a({\u2_Display/n1607 ,\u2_Display/n1608 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c1 ),
    .fco(\u2_Display/lt57_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_30|u2_Display/lt57_29  (
    .a({\u2_Display/n1579 ,\u2_Display/n1580 }),
    .b(2'b01),
    .fci(\u2_Display/lt57_c29 ),
    .fco(\u2_Display/lt57_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_4|u2_Display/lt57_3  (
    .a({\u2_Display/n1605 ,\u2_Display/n1606 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c3 ),
    .fco(\u2_Display/lt57_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_6|u2_Display/lt57_5  (
    .a({\u2_Display/n1603 ,\u2_Display/n1604 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c5 ),
    .fco(\u2_Display/lt57_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_8|u2_Display/lt57_7  (
    .a({\u2_Display/n1601 ,\u2_Display/n1602 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c7 ),
    .fco(\u2_Display/lt57_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_cout|u2_Display/lt57_31  (
    .a({1'b0,\u2_Display/n1578 }),
    .b(2'b10),
    .fci(\u2_Display/lt57_c31 ),
    .f({\u2_Display/n1610 ,open_n104534}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_0|u2_Display/lt58_cin  (
    .a({\u2_Display/n1644 ,1'b0}),
    .b({1'b0,open_n104540}),
    .fco(\u2_Display/lt58_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_10|u2_Display/lt58_9  (
    .a({\u2_Display/n1634 ,\u2_Display/n1635 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c9 ),
    .fco(\u2_Display/lt58_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_12|u2_Display/lt58_11  (
    .a({\u2_Display/n1632 ,\u2_Display/n1633 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c11 ),
    .fco(\u2_Display/lt58_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_14|u2_Display/lt58_13  (
    .a({\u2_Display/n1630 ,\u2_Display/n1631 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c13 ),
    .fco(\u2_Display/lt58_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_16|u2_Display/lt58_15  (
    .a({\u2_Display/n1628 ,\u2_Display/n1629 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c15 ),
    .fco(\u2_Display/lt58_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_18|u2_Display/lt58_17  (
    .a({\u2_Display/n1626 ,\u2_Display/n1627 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c17 ),
    .fco(\u2_Display/lt58_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_20|u2_Display/lt58_19  (
    .a({\u2_Display/n1624 ,\u2_Display/n1625 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c19 ),
    .fco(\u2_Display/lt58_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_22|u2_Display/lt58_21  (
    .a({\u2_Display/n1622 ,\u2_Display/n1623 }),
    .b(2'b01),
    .fci(\u2_Display/lt58_c21 ),
    .fco(\u2_Display/lt58_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_24|u2_Display/lt58_23  (
    .a({\u2_Display/n1620 ,\u2_Display/n1621 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c23 ),
    .fco(\u2_Display/lt58_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_26|u2_Display/lt58_25  (
    .a({\u2_Display/n1618 ,\u2_Display/n1619 }),
    .b(2'b10),
    .fci(\u2_Display/lt58_c25 ),
    .fco(\u2_Display/lt58_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_28|u2_Display/lt58_27  (
    .a({\u2_Display/n1616 ,\u2_Display/n1617 }),
    .b(2'b11),
    .fci(\u2_Display/lt58_c27 ),
    .fco(\u2_Display/lt58_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_2|u2_Display/lt58_1  (
    .a({\u2_Display/n1642 ,\u2_Display/n1643 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c1 ),
    .fco(\u2_Display/lt58_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_30|u2_Display/lt58_29  (
    .a({\u2_Display/n1614 ,\u2_Display/n1615 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c29 ),
    .fco(\u2_Display/lt58_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_4|u2_Display/lt58_3  (
    .a({\u2_Display/n1640 ,\u2_Display/n1641 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c3 ),
    .fco(\u2_Display/lt58_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_6|u2_Display/lt58_5  (
    .a({\u2_Display/n1638 ,\u2_Display/n1639 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c5 ),
    .fco(\u2_Display/lt58_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_8|u2_Display/lt58_7  (
    .a({\u2_Display/n1636 ,\u2_Display/n1637 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c7 ),
    .fco(\u2_Display/lt58_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_cout|u2_Display/lt58_31  (
    .a({1'b0,\u2_Display/n1613 }),
    .b(2'b10),
    .fci(\u2_Display/lt58_c31 ),
    .f({\u2_Display/n1645 ,open_n104944}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_0|u2_Display/lt59_cin  (
    .a({\u2_Display/n1679 ,1'b0}),
    .b({1'b0,open_n104950}),
    .fco(\u2_Display/lt59_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_10|u2_Display/lt59_9  (
    .a({\u2_Display/n1669 ,\u2_Display/n1670 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c9 ),
    .fco(\u2_Display/lt59_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_12|u2_Display/lt59_11  (
    .a({\u2_Display/n1667 ,\u2_Display/n1668 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c11 ),
    .fco(\u2_Display/lt59_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_14|u2_Display/lt59_13  (
    .a({\u2_Display/n1665 ,\u2_Display/n1666 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c13 ),
    .fco(\u2_Display/lt59_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_16|u2_Display/lt59_15  (
    .a({\u2_Display/n1663 ,\u2_Display/n1664 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c15 ),
    .fco(\u2_Display/lt59_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_18|u2_Display/lt59_17  (
    .a({\u2_Display/n1661 ,\u2_Display/n1662 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c17 ),
    .fco(\u2_Display/lt59_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_20|u2_Display/lt59_19  (
    .a({\u2_Display/n1659 ,\u2_Display/n1660 }),
    .b(2'b10),
    .fci(\u2_Display/lt59_c19 ),
    .fco(\u2_Display/lt59_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_22|u2_Display/lt59_21  (
    .a({\u2_Display/n1657 ,\u2_Display/n1658 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c21 ),
    .fco(\u2_Display/lt59_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_24|u2_Display/lt59_23  (
    .a({\u2_Display/n1655 ,\u2_Display/n1656 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c23 ),
    .fco(\u2_Display/lt59_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_26|u2_Display/lt59_25  (
    .a({\u2_Display/n1653 ,\u2_Display/n1654 }),
    .b(2'b11),
    .fci(\u2_Display/lt59_c25 ),
    .fco(\u2_Display/lt59_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_28|u2_Display/lt59_27  (
    .a({\u2_Display/n1651 ,\u2_Display/n1652 }),
    .b(2'b01),
    .fci(\u2_Display/lt59_c27 ),
    .fco(\u2_Display/lt59_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_2|u2_Display/lt59_1  (
    .a({\u2_Display/n1677 ,\u2_Display/n1678 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c1 ),
    .fco(\u2_Display/lt59_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_30|u2_Display/lt59_29  (
    .a({\u2_Display/n1649 ,\u2_Display/n1650 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c29 ),
    .fco(\u2_Display/lt59_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_4|u2_Display/lt59_3  (
    .a({\u2_Display/n1675 ,\u2_Display/n1676 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c3 ),
    .fco(\u2_Display/lt59_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_6|u2_Display/lt59_5  (
    .a({\u2_Display/n1673 ,\u2_Display/n1674 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c5 ),
    .fco(\u2_Display/lt59_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_8|u2_Display/lt59_7  (
    .a({\u2_Display/n1671 ,\u2_Display/n1672 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c7 ),
    .fco(\u2_Display/lt59_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_cout|u2_Display/lt59_31  (
    .a({1'b0,\u2_Display/n1648 }),
    .b(2'b10),
    .fci(\u2_Display/lt59_c31 ),
    .f({\u2_Display/n1680 ,open_n105354}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_0|u2_Display/lt5_2_cin  (
    .a({\u2_Display/n96 [0],1'b0}),
    .b({lcd_xpos[0],open_n105360}),
    .fco(\u2_Display/lt5_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_10|u2_Display/lt5_2_9  (
    .a(\u2_Display/n96 [10:9]),
    .b(lcd_xpos[10:9]),
    .fci(\u2_Display/lt5_2_c9 ),
    .fco(\u2_Display/lt5_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_12|u2_Display/lt5_2_11  (
    .a({\u2_Display/n96 [31],\u2_Display/n96 [31]}),
    .b({1'b0,lcd_xpos[11]}),
    .fci(\u2_Display/lt5_2_c11 ),
    .fco(\u2_Display/lt5_2_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_2|u2_Display/lt5_2_1  (
    .a(\u2_Display/n96 [2:1]),
    .b(lcd_xpos[2:1]),
    .fci(\u2_Display/lt5_2_c1 ),
    .fco(\u2_Display/lt5_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_4|u2_Display/lt5_2_3  (
    .a(\u2_Display/n96 [4:3]),
    .b(lcd_xpos[4:3]),
    .fci(\u2_Display/lt5_2_c3 ),
    .fco(\u2_Display/lt5_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_6|u2_Display/lt5_2_5  (
    .a(\u2_Display/n96 [6:5]),
    .b(lcd_xpos[6:5]),
    .fci(\u2_Display/lt5_2_c5 ),
    .fco(\u2_Display/lt5_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_8|u2_Display/lt5_2_7  (
    .a(\u2_Display/n96 [8:7]),
    .b(lcd_xpos[8:7]),
    .fci(\u2_Display/lt5_2_c7 ),
    .fco(\u2_Display/lt5_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_cout_al_u5061  (
    .a({open_n105530,1'b0}),
    .b({open_n105531,1'b1}),
    .fci(\u2_Display/lt5_2_c13 ),
    .f({open_n105550,\u2_Display/n97 }));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_0|u2_Display/lt60_cin  (
    .a({\u2_Display/n1714 ,1'b0}),
    .b({1'b0,open_n105556}),
    .fco(\u2_Display/lt60_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_10|u2_Display/lt60_9  (
    .a({\u2_Display/n1704 ,\u2_Display/n1705 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c9 ),
    .fco(\u2_Display/lt60_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_12|u2_Display/lt60_11  (
    .a({\u2_Display/n1702 ,\u2_Display/n1703 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c11 ),
    .fco(\u2_Display/lt60_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_14|u2_Display/lt60_13  (
    .a({\u2_Display/n1700 ,\u2_Display/n1701 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c13 ),
    .fco(\u2_Display/lt60_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_16|u2_Display/lt60_15  (
    .a({\u2_Display/n1698 ,\u2_Display/n1699 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c15 ),
    .fco(\u2_Display/lt60_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_18|u2_Display/lt60_17  (
    .a({\u2_Display/n1696 ,\u2_Display/n1697 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c17 ),
    .fco(\u2_Display/lt60_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_20|u2_Display/lt60_19  (
    .a({\u2_Display/n1694 ,\u2_Display/n1695 }),
    .b(2'b01),
    .fci(\u2_Display/lt60_c19 ),
    .fco(\u2_Display/lt60_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_22|u2_Display/lt60_21  (
    .a({\u2_Display/n1692 ,\u2_Display/n1693 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c21 ),
    .fco(\u2_Display/lt60_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_24|u2_Display/lt60_23  (
    .a({\u2_Display/n1690 ,\u2_Display/n1691 }),
    .b(2'b10),
    .fci(\u2_Display/lt60_c23 ),
    .fco(\u2_Display/lt60_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_26|u2_Display/lt60_25  (
    .a({\u2_Display/n1688 ,\u2_Display/n1689 }),
    .b(2'b11),
    .fci(\u2_Display/lt60_c25 ),
    .fco(\u2_Display/lt60_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_28|u2_Display/lt60_27  (
    .a({\u2_Display/n1686 ,\u2_Display/n1687 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c27 ),
    .fco(\u2_Display/lt60_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_2|u2_Display/lt60_1  (
    .a({\u2_Display/n1712 ,\u2_Display/n1713 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c1 ),
    .fco(\u2_Display/lt60_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_30|u2_Display/lt60_29  (
    .a({\u2_Display/n1684 ,\u2_Display/n1685 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c29 ),
    .fco(\u2_Display/lt60_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_4|u2_Display/lt60_3  (
    .a({\u2_Display/n1710 ,\u2_Display/n1711 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c3 ),
    .fco(\u2_Display/lt60_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_6|u2_Display/lt60_5  (
    .a({\u2_Display/n1708 ,\u2_Display/n1709 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c5 ),
    .fco(\u2_Display/lt60_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_8|u2_Display/lt60_7  (
    .a({\u2_Display/n1706 ,\u2_Display/n1707 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c7 ),
    .fco(\u2_Display/lt60_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_cout|u2_Display/lt60_31  (
    .a({1'b0,\u2_Display/n1683 }),
    .b(2'b10),
    .fci(\u2_Display/lt60_c31 ),
    .f({\u2_Display/n1715 ,open_n105960}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_0|u2_Display/lt61_cin  (
    .a({\u2_Display/n1749 ,1'b0}),
    .b({1'b0,open_n105966}),
    .fco(\u2_Display/lt61_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_10|u2_Display/lt61_9  (
    .a({\u2_Display/n1739 ,\u2_Display/n1740 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c9 ),
    .fco(\u2_Display/lt61_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_12|u2_Display/lt61_11  (
    .a({\u2_Display/n1737 ,\u2_Display/n1738 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c11 ),
    .fco(\u2_Display/lt61_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_14|u2_Display/lt61_13  (
    .a({\u2_Display/n1735 ,\u2_Display/n1736 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c13 ),
    .fco(\u2_Display/lt61_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_16|u2_Display/lt61_15  (
    .a({\u2_Display/n1733 ,\u2_Display/n1734 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c15 ),
    .fco(\u2_Display/lt61_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_18|u2_Display/lt61_17  (
    .a({\u2_Display/n1731 ,\u2_Display/n1732 }),
    .b(2'b10),
    .fci(\u2_Display/lt61_c17 ),
    .fco(\u2_Display/lt61_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_20|u2_Display/lt61_19  (
    .a({\u2_Display/n1729 ,\u2_Display/n1730 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c19 ),
    .fco(\u2_Display/lt61_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_22|u2_Display/lt61_21  (
    .a({\u2_Display/n1727 ,\u2_Display/n1728 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c21 ),
    .fco(\u2_Display/lt61_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_24|u2_Display/lt61_23  (
    .a({\u2_Display/n1725 ,\u2_Display/n1726 }),
    .b(2'b11),
    .fci(\u2_Display/lt61_c23 ),
    .fco(\u2_Display/lt61_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_26|u2_Display/lt61_25  (
    .a({\u2_Display/n1723 ,\u2_Display/n1724 }),
    .b(2'b01),
    .fci(\u2_Display/lt61_c25 ),
    .fco(\u2_Display/lt61_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_28|u2_Display/lt61_27  (
    .a({\u2_Display/n1721 ,\u2_Display/n1722 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c27 ),
    .fco(\u2_Display/lt61_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_2|u2_Display/lt61_1  (
    .a({\u2_Display/n1747 ,\u2_Display/n1748 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c1 ),
    .fco(\u2_Display/lt61_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_30|u2_Display/lt61_29  (
    .a({\u2_Display/n1719 ,\u2_Display/n1720 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c29 ),
    .fco(\u2_Display/lt61_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_4|u2_Display/lt61_3  (
    .a({\u2_Display/n1745 ,\u2_Display/n1746 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c3 ),
    .fco(\u2_Display/lt61_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_6|u2_Display/lt61_5  (
    .a({\u2_Display/n1743 ,\u2_Display/n1744 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c5 ),
    .fco(\u2_Display/lt61_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_8|u2_Display/lt61_7  (
    .a({\u2_Display/n1741 ,\u2_Display/n1742 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c7 ),
    .fco(\u2_Display/lt61_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_cout|u2_Display/lt61_31  (
    .a({1'b0,\u2_Display/n1718 }),
    .b(2'b10),
    .fci(\u2_Display/lt61_c31 ),
    .f({\u2_Display/n1750 ,open_n106370}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_0|u2_Display/lt62_cin  (
    .a({\u2_Display/n1784 ,1'b0}),
    .b({1'b0,open_n106376}),
    .fco(\u2_Display/lt62_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_10|u2_Display/lt62_9  (
    .a({\u2_Display/n1774 ,\u2_Display/n1775 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c9 ),
    .fco(\u2_Display/lt62_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_12|u2_Display/lt62_11  (
    .a({\u2_Display/n1772 ,\u2_Display/n1773 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c11 ),
    .fco(\u2_Display/lt62_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_14|u2_Display/lt62_13  (
    .a({\u2_Display/n1770 ,\u2_Display/n1771 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c13 ),
    .fco(\u2_Display/lt62_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_16|u2_Display/lt62_15  (
    .a({\u2_Display/n1768 ,\u2_Display/n1769 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c15 ),
    .fco(\u2_Display/lt62_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_18|u2_Display/lt62_17  (
    .a({\u2_Display/n1766 ,\u2_Display/n1767 }),
    .b(2'b01),
    .fci(\u2_Display/lt62_c17 ),
    .fco(\u2_Display/lt62_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_20|u2_Display/lt62_19  (
    .a({\u2_Display/n1764 ,\u2_Display/n1765 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c19 ),
    .fco(\u2_Display/lt62_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_22|u2_Display/lt62_21  (
    .a({\u2_Display/n1762 ,\u2_Display/n1763 }),
    .b(2'b10),
    .fci(\u2_Display/lt62_c21 ),
    .fco(\u2_Display/lt62_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_24|u2_Display/lt62_23  (
    .a({\u2_Display/n1760 ,\u2_Display/n1761 }),
    .b(2'b11),
    .fci(\u2_Display/lt62_c23 ),
    .fco(\u2_Display/lt62_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_26|u2_Display/lt62_25  (
    .a({\u2_Display/n1758 ,\u2_Display/n1759 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c25 ),
    .fco(\u2_Display/lt62_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_28|u2_Display/lt62_27  (
    .a({\u2_Display/n1756 ,\u2_Display/n1757 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c27 ),
    .fco(\u2_Display/lt62_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_2|u2_Display/lt62_1  (
    .a({\u2_Display/n1782 ,\u2_Display/n1783 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c1 ),
    .fco(\u2_Display/lt62_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_30|u2_Display/lt62_29  (
    .a({\u2_Display/n1754 ,\u2_Display/n1755 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c29 ),
    .fco(\u2_Display/lt62_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_4|u2_Display/lt62_3  (
    .a({\u2_Display/n1780 ,\u2_Display/n1781 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c3 ),
    .fco(\u2_Display/lt62_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_6|u2_Display/lt62_5  (
    .a({\u2_Display/n1778 ,\u2_Display/n1779 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c5 ),
    .fco(\u2_Display/lt62_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_8|u2_Display/lt62_7  (
    .a({\u2_Display/n1776 ,\u2_Display/n1777 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c7 ),
    .fco(\u2_Display/lt62_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_cout|u2_Display/lt62_31  (
    .a({1'b0,\u2_Display/n1753 }),
    .b(2'b10),
    .fci(\u2_Display/lt62_c31 ),
    .f({\u2_Display/n1785 ,open_n106780}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_0|u2_Display/lt63_cin  (
    .a({\u2_Display/n1819 ,1'b0}),
    .b({1'b0,open_n106786}),
    .fco(\u2_Display/lt63_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_10|u2_Display/lt63_9  (
    .a({\u2_Display/n1809 ,\u2_Display/n1810 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c9 ),
    .fco(\u2_Display/lt63_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_12|u2_Display/lt63_11  (
    .a({\u2_Display/n1807 ,\u2_Display/n1808 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c11 ),
    .fco(\u2_Display/lt63_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_14|u2_Display/lt63_13  (
    .a({\u2_Display/n1805 ,\u2_Display/n1806 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c13 ),
    .fco(\u2_Display/lt63_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_16|u2_Display/lt63_15  (
    .a({\u2_Display/n1803 ,\u2_Display/n1804 }),
    .b(2'b10),
    .fci(\u2_Display/lt63_c15 ),
    .fco(\u2_Display/lt63_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_18|u2_Display/lt63_17  (
    .a({\u2_Display/n1801 ,\u2_Display/n1802 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c17 ),
    .fco(\u2_Display/lt63_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_20|u2_Display/lt63_19  (
    .a({\u2_Display/n1799 ,\u2_Display/n1800 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c19 ),
    .fco(\u2_Display/lt63_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_22|u2_Display/lt63_21  (
    .a({\u2_Display/n1797 ,\u2_Display/n1798 }),
    .b(2'b11),
    .fci(\u2_Display/lt63_c21 ),
    .fco(\u2_Display/lt63_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_24|u2_Display/lt63_23  (
    .a({\u2_Display/n1795 ,\u2_Display/n1796 }),
    .b(2'b01),
    .fci(\u2_Display/lt63_c23 ),
    .fco(\u2_Display/lt63_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_26|u2_Display/lt63_25  (
    .a({\u2_Display/n1793 ,\u2_Display/n1794 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c25 ),
    .fco(\u2_Display/lt63_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_28|u2_Display/lt63_27  (
    .a({\u2_Display/n1791 ,\u2_Display/n1792 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c27 ),
    .fco(\u2_Display/lt63_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_2|u2_Display/lt63_1  (
    .a({\u2_Display/n1817 ,\u2_Display/n1818 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c1 ),
    .fco(\u2_Display/lt63_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_30|u2_Display/lt63_29  (
    .a({\u2_Display/n1789 ,\u2_Display/n1790 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c29 ),
    .fco(\u2_Display/lt63_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_4|u2_Display/lt63_3  (
    .a({\u2_Display/n1815 ,\u2_Display/n1816 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c3 ),
    .fco(\u2_Display/lt63_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_6|u2_Display/lt63_5  (
    .a({\u2_Display/n1813 ,\u2_Display/n1814 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c5 ),
    .fco(\u2_Display/lt63_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_8|u2_Display/lt63_7  (
    .a({\u2_Display/n1811 ,\u2_Display/n1812 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c7 ),
    .fco(\u2_Display/lt63_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_cout|u2_Display/lt63_31  (
    .a({1'b0,\u2_Display/n1788 }),
    .b(2'b10),
    .fci(\u2_Display/lt63_c31 ),
    .f({\u2_Display/n1820 ,open_n107190}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_0|u2_Display/lt64_cin  (
    .a({\u2_Display/n1854 ,1'b0}),
    .b({1'b0,open_n107196}),
    .fco(\u2_Display/lt64_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_10|u2_Display/lt64_9  (
    .a({\u2_Display/n1844 ,\u2_Display/n1845 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c9 ),
    .fco(\u2_Display/lt64_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_12|u2_Display/lt64_11  (
    .a({\u2_Display/n1842 ,\u2_Display/n1843 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c11 ),
    .fco(\u2_Display/lt64_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_14|u2_Display/lt64_13  (
    .a({\u2_Display/n1840 ,\u2_Display/n1841 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c13 ),
    .fco(\u2_Display/lt64_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_16|u2_Display/lt64_15  (
    .a({\u2_Display/n1838 ,\u2_Display/n1839 }),
    .b(2'b01),
    .fci(\u2_Display/lt64_c15 ),
    .fco(\u2_Display/lt64_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_18|u2_Display/lt64_17  (
    .a({\u2_Display/n1836 ,\u2_Display/n1837 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c17 ),
    .fco(\u2_Display/lt64_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_20|u2_Display/lt64_19  (
    .a({\u2_Display/n1834 ,\u2_Display/n1835 }),
    .b(2'b10),
    .fci(\u2_Display/lt64_c19 ),
    .fco(\u2_Display/lt64_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_22|u2_Display/lt64_21  (
    .a({\u2_Display/n1832 ,\u2_Display/n1833 }),
    .b(2'b11),
    .fci(\u2_Display/lt64_c21 ),
    .fco(\u2_Display/lt64_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_24|u2_Display/lt64_23  (
    .a({\u2_Display/n1830 ,\u2_Display/n1831 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c23 ),
    .fco(\u2_Display/lt64_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_26|u2_Display/lt64_25  (
    .a({\u2_Display/n1828 ,\u2_Display/n1829 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c25 ),
    .fco(\u2_Display/lt64_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_28|u2_Display/lt64_27  (
    .a({\u2_Display/n1826 ,\u2_Display/n1827 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c27 ),
    .fco(\u2_Display/lt64_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_2|u2_Display/lt64_1  (
    .a({\u2_Display/n1852 ,\u2_Display/n1853 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c1 ),
    .fco(\u2_Display/lt64_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_30|u2_Display/lt64_29  (
    .a({\u2_Display/n1824 ,\u2_Display/n1825 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c29 ),
    .fco(\u2_Display/lt64_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_4|u2_Display/lt64_3  (
    .a({\u2_Display/n1850 ,\u2_Display/n1851 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c3 ),
    .fco(\u2_Display/lt64_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_6|u2_Display/lt64_5  (
    .a({\u2_Display/n1848 ,\u2_Display/n1849 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c5 ),
    .fco(\u2_Display/lt64_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_8|u2_Display/lt64_7  (
    .a({\u2_Display/n1846 ,\u2_Display/n1847 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c7 ),
    .fco(\u2_Display/lt64_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_cout|u2_Display/lt64_31  (
    .a({1'b0,\u2_Display/n1823 }),
    .b(2'b10),
    .fci(\u2_Display/lt64_c31 ),
    .f({\u2_Display/n1855 ,open_n107600}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_0|u2_Display/lt65_cin  (
    .a({\u2_Display/n1889 ,1'b0}),
    .b({1'b0,open_n107606}),
    .fco(\u2_Display/lt65_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_10|u2_Display/lt65_9  (
    .a({\u2_Display/n1879 ,\u2_Display/n1880 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c9 ),
    .fco(\u2_Display/lt65_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_12|u2_Display/lt65_11  (
    .a({\u2_Display/n1877 ,\u2_Display/n1878 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c11 ),
    .fco(\u2_Display/lt65_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_14|u2_Display/lt65_13  (
    .a({\u2_Display/n1875 ,\u2_Display/n1876 }),
    .b(2'b10),
    .fci(\u2_Display/lt65_c13 ),
    .fco(\u2_Display/lt65_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_16|u2_Display/lt65_15  (
    .a({\u2_Display/n1873 ,\u2_Display/n1874 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c15 ),
    .fco(\u2_Display/lt65_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_18|u2_Display/lt65_17  (
    .a({\u2_Display/n1871 ,\u2_Display/n1872 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c17 ),
    .fco(\u2_Display/lt65_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_20|u2_Display/lt65_19  (
    .a({\u2_Display/n1869 ,\u2_Display/n1870 }),
    .b(2'b11),
    .fci(\u2_Display/lt65_c19 ),
    .fco(\u2_Display/lt65_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_22|u2_Display/lt65_21  (
    .a({\u2_Display/n1867 ,\u2_Display/n1868 }),
    .b(2'b01),
    .fci(\u2_Display/lt65_c21 ),
    .fco(\u2_Display/lt65_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_24|u2_Display/lt65_23  (
    .a({\u2_Display/n1865 ,\u2_Display/n1866 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c23 ),
    .fco(\u2_Display/lt65_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_26|u2_Display/lt65_25  (
    .a({\u2_Display/n1863 ,\u2_Display/n1864 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c25 ),
    .fco(\u2_Display/lt65_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_28|u2_Display/lt65_27  (
    .a({\u2_Display/n1861 ,\u2_Display/n1862 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c27 ),
    .fco(\u2_Display/lt65_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_2|u2_Display/lt65_1  (
    .a({\u2_Display/n1887 ,\u2_Display/n1888 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c1 ),
    .fco(\u2_Display/lt65_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_30|u2_Display/lt65_29  (
    .a({\u2_Display/n1859 ,\u2_Display/n1860 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c29 ),
    .fco(\u2_Display/lt65_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_4|u2_Display/lt65_3  (
    .a({\u2_Display/n1885 ,\u2_Display/n1886 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c3 ),
    .fco(\u2_Display/lt65_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_6|u2_Display/lt65_5  (
    .a({\u2_Display/n1883 ,\u2_Display/n1884 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c5 ),
    .fco(\u2_Display/lt65_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_8|u2_Display/lt65_7  (
    .a({\u2_Display/n1881 ,\u2_Display/n1882 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c7 ),
    .fco(\u2_Display/lt65_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_cout|u2_Display/lt65_31  (
    .a({1'b0,\u2_Display/n1858 }),
    .b(2'b10),
    .fci(\u2_Display/lt65_c31 ),
    .f({\u2_Display/n1890 ,open_n108010}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_0|u2_Display/lt66_cin  (
    .a({\u2_Display/n1924 ,1'b0}),
    .b({1'b0,open_n108016}),
    .fco(\u2_Display/lt66_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_10|u2_Display/lt66_9  (
    .a({\u2_Display/n1914 ,\u2_Display/n1915 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c9 ),
    .fco(\u2_Display/lt66_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_12|u2_Display/lt66_11  (
    .a({\u2_Display/n1912 ,\u2_Display/n1913 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c11 ),
    .fco(\u2_Display/lt66_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_14|u2_Display/lt66_13  (
    .a({\u2_Display/n1910 ,\u2_Display/n1911 }),
    .b(2'b01),
    .fci(\u2_Display/lt66_c13 ),
    .fco(\u2_Display/lt66_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_16|u2_Display/lt66_15  (
    .a({\u2_Display/n1908 ,\u2_Display/n1909 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c15 ),
    .fco(\u2_Display/lt66_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_18|u2_Display/lt66_17  (
    .a({\u2_Display/n1906 ,\u2_Display/n1907 }),
    .b(2'b10),
    .fci(\u2_Display/lt66_c17 ),
    .fco(\u2_Display/lt66_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_20|u2_Display/lt66_19  (
    .a({\u2_Display/n1904 ,\u2_Display/n1905 }),
    .b(2'b11),
    .fci(\u2_Display/lt66_c19 ),
    .fco(\u2_Display/lt66_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_22|u2_Display/lt66_21  (
    .a({\u2_Display/n1902 ,\u2_Display/n1903 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c21 ),
    .fco(\u2_Display/lt66_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_24|u2_Display/lt66_23  (
    .a({\u2_Display/n1900 ,\u2_Display/n1901 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c23 ),
    .fco(\u2_Display/lt66_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_26|u2_Display/lt66_25  (
    .a({\u2_Display/n1898 ,\u2_Display/n1899 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c25 ),
    .fco(\u2_Display/lt66_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_28|u2_Display/lt66_27  (
    .a({\u2_Display/n1896 ,\u2_Display/n1897 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c27 ),
    .fco(\u2_Display/lt66_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_2|u2_Display/lt66_1  (
    .a({\u2_Display/n1922 ,\u2_Display/n1923 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c1 ),
    .fco(\u2_Display/lt66_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_30|u2_Display/lt66_29  (
    .a({\u2_Display/n1894 ,\u2_Display/n1895 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c29 ),
    .fco(\u2_Display/lt66_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_4|u2_Display/lt66_3  (
    .a({\u2_Display/n1920 ,\u2_Display/n1921 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c3 ),
    .fco(\u2_Display/lt66_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_6|u2_Display/lt66_5  (
    .a({\u2_Display/n1918 ,\u2_Display/n1919 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c5 ),
    .fco(\u2_Display/lt66_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_8|u2_Display/lt66_7  (
    .a({\u2_Display/n1916 ,\u2_Display/n1917 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c7 ),
    .fco(\u2_Display/lt66_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_cout|u2_Display/lt66_31  (
    .a({1'b0,\u2_Display/n1893 }),
    .b(2'b10),
    .fci(\u2_Display/lt66_c31 ),
    .f({\u2_Display/n1925 ,open_n108420}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_0|u2_Display/lt67_cin  (
    .a({\u2_Display/n1959 ,1'b0}),
    .b({1'b0,open_n108426}),
    .fco(\u2_Display/lt67_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_10|u2_Display/lt67_9  (
    .a({\u2_Display/n1949 ,\u2_Display/n1950 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c9 ),
    .fco(\u2_Display/lt67_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_12|u2_Display/lt67_11  (
    .a({\u2_Display/n1947 ,\u2_Display/n1948 }),
    .b(2'b10),
    .fci(\u2_Display/lt67_c11 ),
    .fco(\u2_Display/lt67_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_14|u2_Display/lt67_13  (
    .a({\u2_Display/n1945 ,\u2_Display/n1946 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c13 ),
    .fco(\u2_Display/lt67_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_16|u2_Display/lt67_15  (
    .a({\u2_Display/n1943 ,\u2_Display/n1944 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c15 ),
    .fco(\u2_Display/lt67_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_18|u2_Display/lt67_17  (
    .a({\u2_Display/n1941 ,\u2_Display/n1942 }),
    .b(2'b11),
    .fci(\u2_Display/lt67_c17 ),
    .fco(\u2_Display/lt67_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_20|u2_Display/lt67_19  (
    .a({\u2_Display/n1939 ,\u2_Display/n1940 }),
    .b(2'b01),
    .fci(\u2_Display/lt67_c19 ),
    .fco(\u2_Display/lt67_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_22|u2_Display/lt67_21  (
    .a({\u2_Display/n1937 ,\u2_Display/n1938 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c21 ),
    .fco(\u2_Display/lt67_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_24|u2_Display/lt67_23  (
    .a({\u2_Display/n1935 ,\u2_Display/n1936 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c23 ),
    .fco(\u2_Display/lt67_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_26|u2_Display/lt67_25  (
    .a({\u2_Display/n1933 ,\u2_Display/n1934 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c25 ),
    .fco(\u2_Display/lt67_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_28|u2_Display/lt67_27  (
    .a({\u2_Display/n1931 ,\u2_Display/n1932 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c27 ),
    .fco(\u2_Display/lt67_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_2|u2_Display/lt67_1  (
    .a({\u2_Display/n1957 ,\u2_Display/n1958 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c1 ),
    .fco(\u2_Display/lt67_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_30|u2_Display/lt67_29  (
    .a({\u2_Display/n1929 ,\u2_Display/n1930 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c29 ),
    .fco(\u2_Display/lt67_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_4|u2_Display/lt67_3  (
    .a({\u2_Display/n1955 ,\u2_Display/n1956 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c3 ),
    .fco(\u2_Display/lt67_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_6|u2_Display/lt67_5  (
    .a({\u2_Display/n1953 ,\u2_Display/n1954 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c5 ),
    .fco(\u2_Display/lt67_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_8|u2_Display/lt67_7  (
    .a({\u2_Display/n1951 ,\u2_Display/n1952 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c7 ),
    .fco(\u2_Display/lt67_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_cout|u2_Display/lt67_31  (
    .a({1'b0,\u2_Display/n1928 }),
    .b(2'b10),
    .fci(\u2_Display/lt67_c31 ),
    .f({\u2_Display/n1960 ,open_n108830}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_0|u2_Display/lt68_cin  (
    .a({\u2_Display/n1994 ,1'b0}),
    .b({1'b0,open_n108836}),
    .fco(\u2_Display/lt68_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_10|u2_Display/lt68_9  (
    .a({\u2_Display/n1984 ,\u2_Display/n1985 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c9 ),
    .fco(\u2_Display/lt68_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_12|u2_Display/lt68_11  (
    .a({\u2_Display/n1982 ,\u2_Display/n1983 }),
    .b(2'b01),
    .fci(\u2_Display/lt68_c11 ),
    .fco(\u2_Display/lt68_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_14|u2_Display/lt68_13  (
    .a({\u2_Display/n1980 ,\u2_Display/n1981 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c13 ),
    .fco(\u2_Display/lt68_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_16|u2_Display/lt68_15  (
    .a({\u2_Display/n1978 ,\u2_Display/n1979 }),
    .b(2'b10),
    .fci(\u2_Display/lt68_c15 ),
    .fco(\u2_Display/lt68_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_18|u2_Display/lt68_17  (
    .a({\u2_Display/n1976 ,\u2_Display/n1977 }),
    .b(2'b11),
    .fci(\u2_Display/lt68_c17 ),
    .fco(\u2_Display/lt68_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_20|u2_Display/lt68_19  (
    .a({\u2_Display/n1974 ,\u2_Display/n1975 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c19 ),
    .fco(\u2_Display/lt68_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_22|u2_Display/lt68_21  (
    .a({\u2_Display/n1972 ,\u2_Display/n1973 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c21 ),
    .fco(\u2_Display/lt68_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_24|u2_Display/lt68_23  (
    .a({\u2_Display/n1970 ,\u2_Display/n1971 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c23 ),
    .fco(\u2_Display/lt68_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_26|u2_Display/lt68_25  (
    .a({\u2_Display/n1968 ,\u2_Display/n1969 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c25 ),
    .fco(\u2_Display/lt68_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_28|u2_Display/lt68_27  (
    .a({\u2_Display/n1966 ,\u2_Display/n1967 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c27 ),
    .fco(\u2_Display/lt68_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_2|u2_Display/lt68_1  (
    .a({\u2_Display/n1992 ,\u2_Display/n1993 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c1 ),
    .fco(\u2_Display/lt68_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_30|u2_Display/lt68_29  (
    .a({\u2_Display/n1964 ,\u2_Display/n1965 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c29 ),
    .fco(\u2_Display/lt68_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_4|u2_Display/lt68_3  (
    .a({\u2_Display/n1990 ,\u2_Display/n1991 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c3 ),
    .fco(\u2_Display/lt68_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_6|u2_Display/lt68_5  (
    .a({\u2_Display/n1988 ,\u2_Display/n1989 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c5 ),
    .fco(\u2_Display/lt68_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_8|u2_Display/lt68_7  (
    .a({\u2_Display/n1986 ,\u2_Display/n1987 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c7 ),
    .fco(\u2_Display/lt68_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_cout|u2_Display/lt68_31  (
    .a({1'b0,\u2_Display/n1963 }),
    .b(2'b10),
    .fci(\u2_Display/lt68_c31 ),
    .f({\u2_Display/n1995 ,open_n109240}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_0|u2_Display/lt69_cin  (
    .a({\u2_Display/n2029 ,1'b0}),
    .b({1'b0,open_n109246}),
    .fco(\u2_Display/lt69_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_10|u2_Display/lt69_9  (
    .a({\u2_Display/n2019 ,\u2_Display/n2020 }),
    .b(2'b10),
    .fci(\u2_Display/lt69_c9 ),
    .fco(\u2_Display/lt69_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_12|u2_Display/lt69_11  (
    .a({\u2_Display/n2017 ,\u2_Display/n2018 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c11 ),
    .fco(\u2_Display/lt69_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_14|u2_Display/lt69_13  (
    .a({\u2_Display/n2015 ,\u2_Display/n2016 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c13 ),
    .fco(\u2_Display/lt69_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_16|u2_Display/lt69_15  (
    .a({\u2_Display/n2013 ,\u2_Display/n2014 }),
    .b(2'b11),
    .fci(\u2_Display/lt69_c15 ),
    .fco(\u2_Display/lt69_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_18|u2_Display/lt69_17  (
    .a({\u2_Display/n2011 ,\u2_Display/n2012 }),
    .b(2'b01),
    .fci(\u2_Display/lt69_c17 ),
    .fco(\u2_Display/lt69_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_20|u2_Display/lt69_19  (
    .a({\u2_Display/n2009 ,\u2_Display/n2010 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c19 ),
    .fco(\u2_Display/lt69_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_22|u2_Display/lt69_21  (
    .a({\u2_Display/n2007 ,\u2_Display/n2008 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c21 ),
    .fco(\u2_Display/lt69_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_24|u2_Display/lt69_23  (
    .a({\u2_Display/n2005 ,\u2_Display/n2006 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c23 ),
    .fco(\u2_Display/lt69_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_26|u2_Display/lt69_25  (
    .a({\u2_Display/n2003 ,\u2_Display/n2004 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c25 ),
    .fco(\u2_Display/lt69_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_28|u2_Display/lt69_27  (
    .a({\u2_Display/n2001 ,\u2_Display/n2002 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c27 ),
    .fco(\u2_Display/lt69_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_2|u2_Display/lt69_1  (
    .a({\u2_Display/n2027 ,\u2_Display/n2028 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c1 ),
    .fco(\u2_Display/lt69_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_30|u2_Display/lt69_29  (
    .a({\u2_Display/n1999 ,\u2_Display/n2000 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c29 ),
    .fco(\u2_Display/lt69_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_4|u2_Display/lt69_3  (
    .a({\u2_Display/n2025 ,\u2_Display/n2026 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c3 ),
    .fco(\u2_Display/lt69_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_6|u2_Display/lt69_5  (
    .a({\u2_Display/n2023 ,\u2_Display/n2024 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c5 ),
    .fco(\u2_Display/lt69_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_8|u2_Display/lt69_7  (
    .a({\u2_Display/n2021 ,\u2_Display/n2022 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c7 ),
    .fco(\u2_Display/lt69_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_cout|u2_Display/lt69_31  (
    .a({1'b0,\u2_Display/n1998 }),
    .b(2'b10),
    .fci(\u2_Display/lt69_c31 ),
    .f({\u2_Display/n2030 ,open_n109650}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_0|u2_Display/lt6_2_cin  (
    .a({lcd_ypos[0],1'b0}),
    .b({\u2_Display/j [0],open_n109656}),
    .fco(\u2_Display/lt6_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_10|u2_Display/lt6_2_9  (
    .a(lcd_ypos[10:9]),
    .b({\u2_Display/j [9],\u2_Display/n99 [0]}),
    .fci(\u2_Display/lt6_2_c9 ),
    .fco(\u2_Display/lt6_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_2|u2_Display/lt6_2_1  (
    .a(lcd_ypos[2:1]),
    .b(\u2_Display/j [2:1]),
    .fci(\u2_Display/lt6_2_c1 ),
    .fco(\u2_Display/lt6_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_4|u2_Display/lt6_2_3  (
    .a(lcd_ypos[4:3]),
    .b(\u2_Display/j [4:3]),
    .fci(\u2_Display/lt6_2_c3 ),
    .fco(\u2_Display/lt6_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_6|u2_Display/lt6_2_5  (
    .a(lcd_ypos[6:5]),
    .b(\u2_Display/j [6:5]),
    .fci(\u2_Display/lt6_2_c5 ),
    .fco(\u2_Display/lt6_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_8|u2_Display/lt6_2_7  (
    .a(lcd_ypos[8:7]),
    .b(\u2_Display/j [8:7]),
    .fci(\u2_Display/lt6_2_c7 ),
    .fco(\u2_Display/lt6_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_cout|u2_Display/lt6_2_11  (
    .a({1'b0,lcd_ypos[11]}),
    .b(2'b10),
    .fci(\u2_Display/lt6_2_c11 ),
    .f({\u2_Display/n100 ,open_n109820}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_0|u2_Display/lt70_cin  (
    .a({\u2_Display/n2064 ,1'b0}),
    .b({1'b0,open_n109826}),
    .fco(\u2_Display/lt70_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_10|u2_Display/lt70_9  (
    .a({\u2_Display/n2054 ,\u2_Display/n2055 }),
    .b(2'b01),
    .fci(\u2_Display/lt70_c9 ),
    .fco(\u2_Display/lt70_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_12|u2_Display/lt70_11  (
    .a({\u2_Display/n2052 ,\u2_Display/n2053 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c11 ),
    .fco(\u2_Display/lt70_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_14|u2_Display/lt70_13  (
    .a({\u2_Display/n2050 ,\u2_Display/n2051 }),
    .b(2'b10),
    .fci(\u2_Display/lt70_c13 ),
    .fco(\u2_Display/lt70_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_16|u2_Display/lt70_15  (
    .a({\u2_Display/n2048 ,\u2_Display/n2049 }),
    .b(2'b11),
    .fci(\u2_Display/lt70_c15 ),
    .fco(\u2_Display/lt70_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_18|u2_Display/lt70_17  (
    .a({\u2_Display/n2046 ,\u2_Display/n2047 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c17 ),
    .fco(\u2_Display/lt70_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_20|u2_Display/lt70_19  (
    .a({\u2_Display/n2044 ,\u2_Display/n2045 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c19 ),
    .fco(\u2_Display/lt70_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_22|u2_Display/lt70_21  (
    .a({\u2_Display/n2042 ,\u2_Display/n2043 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c21 ),
    .fco(\u2_Display/lt70_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_24|u2_Display/lt70_23  (
    .a({\u2_Display/n2040 ,\u2_Display/n2041 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c23 ),
    .fco(\u2_Display/lt70_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_26|u2_Display/lt70_25  (
    .a({\u2_Display/n2038 ,\u2_Display/n2039 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c25 ),
    .fco(\u2_Display/lt70_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_28|u2_Display/lt70_27  (
    .a({\u2_Display/n2036 ,\u2_Display/n2037 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c27 ),
    .fco(\u2_Display/lt70_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_2|u2_Display/lt70_1  (
    .a({\u2_Display/n2062 ,\u2_Display/n2063 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c1 ),
    .fco(\u2_Display/lt70_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_30|u2_Display/lt70_29  (
    .a({\u2_Display/n2034 ,\u2_Display/n2035 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c29 ),
    .fco(\u2_Display/lt70_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_4|u2_Display/lt70_3  (
    .a({\u2_Display/n2060 ,\u2_Display/n2061 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c3 ),
    .fco(\u2_Display/lt70_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_6|u2_Display/lt70_5  (
    .a({\u2_Display/n2058 ,\u2_Display/n2059 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c5 ),
    .fco(\u2_Display/lt70_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_8|u2_Display/lt70_7  (
    .a({\u2_Display/n2056 ,\u2_Display/n2057 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c7 ),
    .fco(\u2_Display/lt70_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_cout|u2_Display/lt70_31  (
    .a({1'b0,\u2_Display/n2033 }),
    .b(2'b10),
    .fci(\u2_Display/lt70_c31 ),
    .f({\u2_Display/n2065 ,open_n110230}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_0|u2_Display/lt71_cin  (
    .a({\u2_Display/n2099 ,1'b0}),
    .b({1'b0,open_n110236}),
    .fco(\u2_Display/lt71_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_10|u2_Display/lt71_9  (
    .a({\u2_Display/n2089 ,\u2_Display/n2090 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c9 ),
    .fco(\u2_Display/lt71_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_12|u2_Display/lt71_11  (
    .a({\u2_Display/n2087 ,\u2_Display/n2088 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c11 ),
    .fco(\u2_Display/lt71_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_14|u2_Display/lt71_13  (
    .a({\u2_Display/n2085 ,\u2_Display/n2086 }),
    .b(2'b11),
    .fci(\u2_Display/lt71_c13 ),
    .fco(\u2_Display/lt71_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_16|u2_Display/lt71_15  (
    .a({\u2_Display/n2083 ,\u2_Display/n2084 }),
    .b(2'b01),
    .fci(\u2_Display/lt71_c15 ),
    .fco(\u2_Display/lt71_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_18|u2_Display/lt71_17  (
    .a({\u2_Display/n2081 ,\u2_Display/n2082 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c17 ),
    .fco(\u2_Display/lt71_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_20|u2_Display/lt71_19  (
    .a({\u2_Display/n2079 ,\u2_Display/n2080 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c19 ),
    .fco(\u2_Display/lt71_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_22|u2_Display/lt71_21  (
    .a({\u2_Display/n2077 ,\u2_Display/n2078 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c21 ),
    .fco(\u2_Display/lt71_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_24|u2_Display/lt71_23  (
    .a({\u2_Display/n2075 ,\u2_Display/n2076 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c23 ),
    .fco(\u2_Display/lt71_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_26|u2_Display/lt71_25  (
    .a({\u2_Display/n2073 ,\u2_Display/n2074 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c25 ),
    .fco(\u2_Display/lt71_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_28|u2_Display/lt71_27  (
    .a({\u2_Display/n2071 ,\u2_Display/n2072 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c27 ),
    .fco(\u2_Display/lt71_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_2|u2_Display/lt71_1  (
    .a({\u2_Display/n2097 ,\u2_Display/n2098 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c1 ),
    .fco(\u2_Display/lt71_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_30|u2_Display/lt71_29  (
    .a({\u2_Display/n2069 ,\u2_Display/n2070 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c29 ),
    .fco(\u2_Display/lt71_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_4|u2_Display/lt71_3  (
    .a({\u2_Display/n2095 ,\u2_Display/n2096 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c3 ),
    .fco(\u2_Display/lt71_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_6|u2_Display/lt71_5  (
    .a({\u2_Display/n2093 ,\u2_Display/n2094 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c5 ),
    .fco(\u2_Display/lt71_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_8|u2_Display/lt71_7  (
    .a({\u2_Display/n2091 ,\u2_Display/n2092 }),
    .b(2'b10),
    .fci(\u2_Display/lt71_c7 ),
    .fco(\u2_Display/lt71_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_cout|u2_Display/lt71_31  (
    .a({1'b0,\u2_Display/n2068 }),
    .b(2'b10),
    .fci(\u2_Display/lt71_c31 ),
    .f({\u2_Display/n2100 ,open_n110640}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_0|u2_Display/lt72_cin  (
    .a({\u2_Display/n2134 ,1'b0}),
    .b({1'b0,open_n110646}),
    .fco(\u2_Display/lt72_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_10|u2_Display/lt72_9  (
    .a({\u2_Display/n2124 ,\u2_Display/n2125 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c9 ),
    .fco(\u2_Display/lt72_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_12|u2_Display/lt72_11  (
    .a({\u2_Display/n2122 ,\u2_Display/n2123 }),
    .b(2'b10),
    .fci(\u2_Display/lt72_c11 ),
    .fco(\u2_Display/lt72_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_14|u2_Display/lt72_13  (
    .a({\u2_Display/n2120 ,\u2_Display/n2121 }),
    .b(2'b11),
    .fci(\u2_Display/lt72_c13 ),
    .fco(\u2_Display/lt72_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_16|u2_Display/lt72_15  (
    .a({\u2_Display/n2118 ,\u2_Display/n2119 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c15 ),
    .fco(\u2_Display/lt72_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_18|u2_Display/lt72_17  (
    .a({\u2_Display/n2116 ,\u2_Display/n2117 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c17 ),
    .fco(\u2_Display/lt72_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_20|u2_Display/lt72_19  (
    .a({\u2_Display/n2114 ,\u2_Display/n2115 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c19 ),
    .fco(\u2_Display/lt72_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_22|u2_Display/lt72_21  (
    .a({\u2_Display/n2112 ,\u2_Display/n2113 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c21 ),
    .fco(\u2_Display/lt72_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_24|u2_Display/lt72_23  (
    .a({\u2_Display/n2110 ,\u2_Display/n2111 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c23 ),
    .fco(\u2_Display/lt72_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_26|u2_Display/lt72_25  (
    .a({\u2_Display/n2108 ,\u2_Display/n2109 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c25 ),
    .fco(\u2_Display/lt72_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_28|u2_Display/lt72_27  (
    .a({\u2_Display/n2106 ,\u2_Display/n2107 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c27 ),
    .fco(\u2_Display/lt72_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_2|u2_Display/lt72_1  (
    .a({\u2_Display/n2132 ,\u2_Display/n2133 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c1 ),
    .fco(\u2_Display/lt72_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_30|u2_Display/lt72_29  (
    .a({\u2_Display/n2104 ,\u2_Display/n2105 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c29 ),
    .fco(\u2_Display/lt72_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_4|u2_Display/lt72_3  (
    .a({\u2_Display/n2130 ,\u2_Display/n2131 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c3 ),
    .fco(\u2_Display/lt72_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_6|u2_Display/lt72_5  (
    .a({\u2_Display/n2128 ,\u2_Display/n2129 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c5 ),
    .fco(\u2_Display/lt72_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_8|u2_Display/lt72_7  (
    .a({\u2_Display/n2126 ,\u2_Display/n2127 }),
    .b(2'b01),
    .fci(\u2_Display/lt72_c7 ),
    .fco(\u2_Display/lt72_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_cout|u2_Display/lt72_31  (
    .a({1'b0,\u2_Display/n2103 }),
    .b(2'b10),
    .fci(\u2_Display/lt72_c31 ),
    .f({\u2_Display/n2135 ,open_n111050}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_0|u2_Display/lt73_cin  (
    .a({\u2_Display/n2169 ,1'b0}),
    .b({1'b0,open_n111056}),
    .fco(\u2_Display/lt73_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_10|u2_Display/lt73_9  (
    .a({\u2_Display/n2159 ,\u2_Display/n2160 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c9 ),
    .fco(\u2_Display/lt73_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_12|u2_Display/lt73_11  (
    .a({\u2_Display/n2157 ,\u2_Display/n2158 }),
    .b(2'b11),
    .fci(\u2_Display/lt73_c11 ),
    .fco(\u2_Display/lt73_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_14|u2_Display/lt73_13  (
    .a({\u2_Display/n2155 ,\u2_Display/n2156 }),
    .b(2'b01),
    .fci(\u2_Display/lt73_c13 ),
    .fco(\u2_Display/lt73_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_16|u2_Display/lt73_15  (
    .a({\u2_Display/n2153 ,\u2_Display/n2154 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c15 ),
    .fco(\u2_Display/lt73_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_18|u2_Display/lt73_17  (
    .a({\u2_Display/n2151 ,\u2_Display/n2152 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c17 ),
    .fco(\u2_Display/lt73_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_20|u2_Display/lt73_19  (
    .a({\u2_Display/n2149 ,\u2_Display/n2150 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c19 ),
    .fco(\u2_Display/lt73_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_22|u2_Display/lt73_21  (
    .a({\u2_Display/n2147 ,\u2_Display/n2148 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c21 ),
    .fco(\u2_Display/lt73_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_24|u2_Display/lt73_23  (
    .a({\u2_Display/n2145 ,\u2_Display/n2146 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c23 ),
    .fco(\u2_Display/lt73_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_26|u2_Display/lt73_25  (
    .a({\u2_Display/n2143 ,\u2_Display/n2144 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c25 ),
    .fco(\u2_Display/lt73_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_28|u2_Display/lt73_27  (
    .a({\u2_Display/n2141 ,\u2_Display/n2142 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c27 ),
    .fco(\u2_Display/lt73_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_2|u2_Display/lt73_1  (
    .a({\u2_Display/n2167 ,\u2_Display/n2168 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c1 ),
    .fco(\u2_Display/lt73_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_30|u2_Display/lt73_29  (
    .a({\u2_Display/n2139 ,\u2_Display/n2140 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c29 ),
    .fco(\u2_Display/lt73_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_4|u2_Display/lt73_3  (
    .a({\u2_Display/n2165 ,\u2_Display/n2166 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c3 ),
    .fco(\u2_Display/lt73_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_6|u2_Display/lt73_5  (
    .a({\u2_Display/n2163 ,\u2_Display/n2164 }),
    .b(2'b10),
    .fci(\u2_Display/lt73_c5 ),
    .fco(\u2_Display/lt73_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_8|u2_Display/lt73_7  (
    .a({\u2_Display/n2161 ,\u2_Display/n2162 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c7 ),
    .fco(\u2_Display/lt73_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_cout|u2_Display/lt73_31  (
    .a({1'b0,\u2_Display/n2138 }),
    .b(2'b10),
    .fci(\u2_Display/lt73_c31 ),
    .f({\u2_Display/n2170 ,open_n111460}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_0|u2_Display/lt74_cin  (
    .a({\u2_Display/n2204 ,1'b0}),
    .b({1'b0,open_n111466}),
    .fco(\u2_Display/lt74_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_10|u2_Display/lt74_9  (
    .a({\u2_Display/n2194 ,\u2_Display/n2195 }),
    .b(2'b10),
    .fci(\u2_Display/lt74_c9 ),
    .fco(\u2_Display/lt74_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_12|u2_Display/lt74_11  (
    .a({\u2_Display/n2192 ,\u2_Display/n2193 }),
    .b(2'b11),
    .fci(\u2_Display/lt74_c11 ),
    .fco(\u2_Display/lt74_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_14|u2_Display/lt74_13  (
    .a({\u2_Display/n2190 ,\u2_Display/n2191 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c13 ),
    .fco(\u2_Display/lt74_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_16|u2_Display/lt74_15  (
    .a({\u2_Display/n2188 ,\u2_Display/n2189 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c15 ),
    .fco(\u2_Display/lt74_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_18|u2_Display/lt74_17  (
    .a({\u2_Display/n2186 ,\u2_Display/n2187 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c17 ),
    .fco(\u2_Display/lt74_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_20|u2_Display/lt74_19  (
    .a({\u2_Display/n2184 ,\u2_Display/n2185 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c19 ),
    .fco(\u2_Display/lt74_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_22|u2_Display/lt74_21  (
    .a({\u2_Display/n2182 ,\u2_Display/n2183 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c21 ),
    .fco(\u2_Display/lt74_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_24|u2_Display/lt74_23  (
    .a({\u2_Display/n2180 ,\u2_Display/n2181 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c23 ),
    .fco(\u2_Display/lt74_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_26|u2_Display/lt74_25  (
    .a({\u2_Display/n2178 ,\u2_Display/n2179 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c25 ),
    .fco(\u2_Display/lt74_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_28|u2_Display/lt74_27  (
    .a({\u2_Display/n2176 ,\u2_Display/n2177 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c27 ),
    .fco(\u2_Display/lt74_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_2|u2_Display/lt74_1  (
    .a({\u2_Display/n2202 ,\u2_Display/n2203 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c1 ),
    .fco(\u2_Display/lt74_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_30|u2_Display/lt74_29  (
    .a({\u2_Display/n2174 ,\u2_Display/n2175 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c29 ),
    .fco(\u2_Display/lt74_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_4|u2_Display/lt74_3  (
    .a({\u2_Display/n2200 ,\u2_Display/n2201 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c3 ),
    .fco(\u2_Display/lt74_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_6|u2_Display/lt74_5  (
    .a({\u2_Display/n2198 ,\u2_Display/n2199 }),
    .b(2'b01),
    .fci(\u2_Display/lt74_c5 ),
    .fco(\u2_Display/lt74_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_8|u2_Display/lt74_7  (
    .a({\u2_Display/n2196 ,\u2_Display/n2197 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c7 ),
    .fco(\u2_Display/lt74_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_cout|u2_Display/lt74_31  (
    .a({1'b0,\u2_Display/n2173 }),
    .b(2'b10),
    .fci(\u2_Display/lt74_c31 ),
    .f({\u2_Display/n2205 ,open_n111870}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_0|u2_Display/lt75_cin  (
    .a({\u2_Display/n2239 ,1'b0}),
    .b({1'b0,open_n111876}),
    .fco(\u2_Display/lt75_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_10|u2_Display/lt75_9  (
    .a({\u2_Display/n2229 ,\u2_Display/n2230 }),
    .b(2'b11),
    .fci(\u2_Display/lt75_c9 ),
    .fco(\u2_Display/lt75_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_12|u2_Display/lt75_11  (
    .a({\u2_Display/n2227 ,\u2_Display/n2228 }),
    .b(2'b01),
    .fci(\u2_Display/lt75_c11 ),
    .fco(\u2_Display/lt75_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_14|u2_Display/lt75_13  (
    .a({\u2_Display/n2225 ,\u2_Display/n2226 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c13 ),
    .fco(\u2_Display/lt75_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_16|u2_Display/lt75_15  (
    .a({\u2_Display/n2223 ,\u2_Display/n2224 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c15 ),
    .fco(\u2_Display/lt75_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_18|u2_Display/lt75_17  (
    .a({\u2_Display/n2221 ,\u2_Display/n2222 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c17 ),
    .fco(\u2_Display/lt75_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_20|u2_Display/lt75_19  (
    .a({\u2_Display/n2219 ,\u2_Display/n2220 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c19 ),
    .fco(\u2_Display/lt75_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_22|u2_Display/lt75_21  (
    .a({\u2_Display/n2217 ,\u2_Display/n2218 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c21 ),
    .fco(\u2_Display/lt75_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_24|u2_Display/lt75_23  (
    .a({\u2_Display/n2215 ,\u2_Display/n2216 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c23 ),
    .fco(\u2_Display/lt75_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_26|u2_Display/lt75_25  (
    .a({\u2_Display/n2213 ,\u2_Display/n2214 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c25 ),
    .fco(\u2_Display/lt75_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_28|u2_Display/lt75_27  (
    .a({\u2_Display/n2211 ,\u2_Display/n2212 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c27 ),
    .fco(\u2_Display/lt75_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_2|u2_Display/lt75_1  (
    .a({\u2_Display/n2237 ,\u2_Display/n2238 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c1 ),
    .fco(\u2_Display/lt75_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_30|u2_Display/lt75_29  (
    .a({\u2_Display/n2209 ,\u2_Display/n2210 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c29 ),
    .fco(\u2_Display/lt75_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_4|u2_Display/lt75_3  (
    .a({\u2_Display/n2235 ,\u2_Display/n2236 }),
    .b(2'b10),
    .fci(\u2_Display/lt75_c3 ),
    .fco(\u2_Display/lt75_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_6|u2_Display/lt75_5  (
    .a({\u2_Display/n2233 ,\u2_Display/n2234 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c5 ),
    .fco(\u2_Display/lt75_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_8|u2_Display/lt75_7  (
    .a({\u2_Display/n2231 ,\u2_Display/n2232 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c7 ),
    .fco(\u2_Display/lt75_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_cout|u2_Display/lt75_31  (
    .a({1'b0,\u2_Display/n2208 }),
    .b(2'b10),
    .fci(\u2_Display/lt75_c31 ),
    .f({\u2_Display/n2240 ,open_n112280}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_0|u2_Display/lt76_cin  (
    .a({\u2_Display/n2274 ,1'b0}),
    .b({1'b0,open_n112286}),
    .fco(\u2_Display/lt76_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_10|u2_Display/lt76_9  (
    .a({\u2_Display/n2264 ,\u2_Display/n2265 }),
    .b(2'b11),
    .fci(\u2_Display/lt76_c9 ),
    .fco(\u2_Display/lt76_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_12|u2_Display/lt76_11  (
    .a({\u2_Display/n2262 ,\u2_Display/n2263 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c11 ),
    .fco(\u2_Display/lt76_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_14|u2_Display/lt76_13  (
    .a({\u2_Display/n2260 ,\u2_Display/n2261 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c13 ),
    .fco(\u2_Display/lt76_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_16|u2_Display/lt76_15  (
    .a({\u2_Display/n2258 ,\u2_Display/n2259 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c15 ),
    .fco(\u2_Display/lt76_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_18|u2_Display/lt76_17  (
    .a({\u2_Display/n2256 ,\u2_Display/n2257 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c17 ),
    .fco(\u2_Display/lt76_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_20|u2_Display/lt76_19  (
    .a({\u2_Display/n2254 ,\u2_Display/n2255 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c19 ),
    .fco(\u2_Display/lt76_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_22|u2_Display/lt76_21  (
    .a({\u2_Display/n2252 ,\u2_Display/n2253 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c21 ),
    .fco(\u2_Display/lt76_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_24|u2_Display/lt76_23  (
    .a({\u2_Display/n2250 ,\u2_Display/n2251 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c23 ),
    .fco(\u2_Display/lt76_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_26|u2_Display/lt76_25  (
    .a({\u2_Display/n2248 ,\u2_Display/n2249 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c25 ),
    .fco(\u2_Display/lt76_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_28|u2_Display/lt76_27  (
    .a({\u2_Display/n2246 ,\u2_Display/n2247 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c27 ),
    .fco(\u2_Display/lt76_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_2|u2_Display/lt76_1  (
    .a({\u2_Display/n2272 ,\u2_Display/n2273 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c1 ),
    .fco(\u2_Display/lt76_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_30|u2_Display/lt76_29  (
    .a({\u2_Display/n2244 ,\u2_Display/n2245 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c29 ),
    .fco(\u2_Display/lt76_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_4|u2_Display/lt76_3  (
    .a({\u2_Display/n2270 ,\u2_Display/n2271 }),
    .b(2'b01),
    .fci(\u2_Display/lt76_c3 ),
    .fco(\u2_Display/lt76_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_6|u2_Display/lt76_5  (
    .a({\u2_Display/n2268 ,\u2_Display/n2269 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c5 ),
    .fco(\u2_Display/lt76_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_8|u2_Display/lt76_7  (
    .a({\u2_Display/n2266 ,\u2_Display/n2267 }),
    .b(2'b10),
    .fci(\u2_Display/lt76_c7 ),
    .fco(\u2_Display/lt76_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_cout|u2_Display/lt76_31  (
    .a({1'b0,\u2_Display/n2243 }),
    .b(2'b10),
    .fci(\u2_Display/lt76_c31 ),
    .f({\u2_Display/n2275 ,open_n112690}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_0|u2_Display/lt77_cin  (
    .a({\u2_Display/n2309 ,1'b0}),
    .b({1'b0,open_n112696}),
    .fco(\u2_Display/lt77_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_10|u2_Display/lt77_9  (
    .a({\u2_Display/n2299 ,\u2_Display/n2300 }),
    .b(2'b01),
    .fci(\u2_Display/lt77_c9 ),
    .fco(\u2_Display/lt77_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_12|u2_Display/lt77_11  (
    .a({\u2_Display/n2297 ,\u2_Display/n2298 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c11 ),
    .fco(\u2_Display/lt77_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_14|u2_Display/lt77_13  (
    .a({\u2_Display/n2295 ,\u2_Display/n2296 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c13 ),
    .fco(\u2_Display/lt77_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_16|u2_Display/lt77_15  (
    .a({\u2_Display/n2293 ,\u2_Display/n2294 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c15 ),
    .fco(\u2_Display/lt77_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_18|u2_Display/lt77_17  (
    .a({\u2_Display/n2291 ,\u2_Display/n2292 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c17 ),
    .fco(\u2_Display/lt77_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_20|u2_Display/lt77_19  (
    .a({\u2_Display/n2289 ,\u2_Display/n2290 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c19 ),
    .fco(\u2_Display/lt77_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_22|u2_Display/lt77_21  (
    .a({\u2_Display/n2287 ,\u2_Display/n2288 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c21 ),
    .fco(\u2_Display/lt77_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_24|u2_Display/lt77_23  (
    .a({\u2_Display/n2285 ,\u2_Display/n2286 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c23 ),
    .fco(\u2_Display/lt77_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_26|u2_Display/lt77_25  (
    .a({\u2_Display/n2283 ,\u2_Display/n2284 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c25 ),
    .fco(\u2_Display/lt77_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_28|u2_Display/lt77_27  (
    .a({\u2_Display/n2281 ,\u2_Display/n2282 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c27 ),
    .fco(\u2_Display/lt77_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_2|u2_Display/lt77_1  (
    .a({\u2_Display/n2307 ,\u2_Display/n2308 }),
    .b(2'b10),
    .fci(\u2_Display/lt77_c1 ),
    .fco(\u2_Display/lt77_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_30|u2_Display/lt77_29  (
    .a({\u2_Display/n2279 ,\u2_Display/n2280 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c29 ),
    .fco(\u2_Display/lt77_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_4|u2_Display/lt77_3  (
    .a({\u2_Display/n2305 ,\u2_Display/n2306 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c3 ),
    .fco(\u2_Display/lt77_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_6|u2_Display/lt77_5  (
    .a({\u2_Display/n2303 ,\u2_Display/n2304 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c5 ),
    .fco(\u2_Display/lt77_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_8|u2_Display/lt77_7  (
    .a({\u2_Display/n2301 ,\u2_Display/n2302 }),
    .b(2'b11),
    .fci(\u2_Display/lt77_c7 ),
    .fco(\u2_Display/lt77_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_cout|u2_Display/lt77_31  (
    .a({1'b0,\u2_Display/n2278 }),
    .b(2'b10),
    .fci(\u2_Display/lt77_c31 ),
    .f({\u2_Display/n2310 ,open_n113100}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_0|u2_Display/lt7_2_cin  (
    .a({\u2_Display/n102 [0],1'b0}),
    .b({lcd_ypos[0],open_n113106}),
    .fco(\u2_Display/lt7_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_10|u2_Display/lt7_2_9  (
    .a({\u2_Display/n102 [31],\u2_Display/n102 [9]}),
    .b(lcd_ypos[10:9]),
    .fci(\u2_Display/lt7_2_c9 ),
    .fco(\u2_Display/lt7_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_12|u2_Display/lt7_2_11  (
    .a({\u2_Display/n102 [31],\u2_Display/n102 [31]}),
    .b({1'b0,lcd_ypos[11]}),
    .fci(\u2_Display/lt7_2_c11 ),
    .fco(\u2_Display/lt7_2_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_2|u2_Display/lt7_2_1  (
    .a(\u2_Display/n102 [2:1]),
    .b(lcd_ypos[2:1]),
    .fci(\u2_Display/lt7_2_c1 ),
    .fco(\u2_Display/lt7_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_4|u2_Display/lt7_2_3  (
    .a(\u2_Display/n102 [4:3]),
    .b(lcd_ypos[4:3]),
    .fci(\u2_Display/lt7_2_c3 ),
    .fco(\u2_Display/lt7_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_6|u2_Display/lt7_2_5  (
    .a(\u2_Display/n102 [6:5]),
    .b(lcd_ypos[6:5]),
    .fci(\u2_Display/lt7_2_c5 ),
    .fco(\u2_Display/lt7_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_8|u2_Display/lt7_2_7  (
    .a(\u2_Display/n102 [8:7]),
    .b(lcd_ypos[8:7]),
    .fci(\u2_Display/lt7_2_c7 ),
    .fco(\u2_Display/lt7_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_cout_al_u5062  (
    .a({open_n113276,1'b0}),
    .b({open_n113277,1'b1}),
    .fci(\u2_Display/lt7_2_c13 ),
    .f({open_n113296,\u2_Display/n103 }));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_0|u2_Display/lt88_cin  (
    .a({\u2_Display/counta [0],1'b0}),
    .b({1'b0,open_n113302}),
    .fco(\u2_Display/lt88_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_10|u2_Display/lt88_9  (
    .a(\u2_Display/counta [10:9]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c9 ),
    .fco(\u2_Display/lt88_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_12|u2_Display/lt88_11  (
    .a(\u2_Display/counta [12:11]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c11 ),
    .fco(\u2_Display/lt88_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_14|u2_Display/lt88_13  (
    .a(\u2_Display/counta [14:13]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c13 ),
    .fco(\u2_Display/lt88_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_16|u2_Display/lt88_15  (
    .a(\u2_Display/counta [16:15]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c15 ),
    .fco(\u2_Display/lt88_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_18|u2_Display/lt88_17  (
    .a(\u2_Display/counta [18:17]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c17 ),
    .fco(\u2_Display/lt88_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_20|u2_Display/lt88_19  (
    .a(\u2_Display/counta [20:19]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c19 ),
    .fco(\u2_Display/lt88_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_22|u2_Display/lt88_21  (
    .a(\u2_Display/counta [22:21]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c21 ),
    .fco(\u2_Display/lt88_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_24|u2_Display/lt88_23  (
    .a(\u2_Display/counta [24:23]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c23 ),
    .fco(\u2_Display/lt88_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_26|u2_Display/lt88_25  (
    .a(\u2_Display/counta [26:25]),
    .b(2'b11),
    .fci(\u2_Display/lt88_c25 ),
    .fco(\u2_Display/lt88_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_28|u2_Display/lt88_27  (
    .a(\u2_Display/counta [28:27]),
    .b(2'b10),
    .fci(\u2_Display/lt88_c27 ),
    .fco(\u2_Display/lt88_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_2|u2_Display/lt88_1  (
    .a(\u2_Display/counta [2:1]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c1 ),
    .fco(\u2_Display/lt88_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_30|u2_Display/lt88_29  (
    .a(\u2_Display/counta [30:29]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c29 ),
    .fco(\u2_Display/lt88_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_4|u2_Display/lt88_3  (
    .a(\u2_Display/counta [4:3]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c3 ),
    .fco(\u2_Display/lt88_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_6|u2_Display/lt88_5  (
    .a(\u2_Display/counta [6:5]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c5 ),
    .fco(\u2_Display/lt88_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_8|u2_Display/lt88_7  (
    .a(\u2_Display/counta [8:7]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c7 ),
    .fco(\u2_Display/lt88_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_cout|u2_Display/lt88_31  (
    .a({1'b0,\u2_Display/counta [31]}),
    .b(2'b11),
    .fci(\u2_Display/lt88_c31 ),
    .f({\u2_Display/n2663 ,open_n113706}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_0|u2_Display/lt89_cin  (
    .a({\u2_Display/n2697 ,1'b0}),
    .b({1'b0,open_n113712}),
    .fco(\u2_Display/lt89_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_10|u2_Display/lt89_9  (
    .a({\u2_Display/n2687 ,\u2_Display/n2688 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c9 ),
    .fco(\u2_Display/lt89_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_12|u2_Display/lt89_11  (
    .a({\u2_Display/n2685 ,\u2_Display/n2686 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c11 ),
    .fco(\u2_Display/lt89_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_14|u2_Display/lt89_13  (
    .a({\u2_Display/n2683 ,\u2_Display/n2684 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c13 ),
    .fco(\u2_Display/lt89_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_16|u2_Display/lt89_15  (
    .a({\u2_Display/n2681 ,\u2_Display/n2682 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c15 ),
    .fco(\u2_Display/lt89_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_18|u2_Display/lt89_17  (
    .a({\u2_Display/n2679 ,\u2_Display/n2680 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c17 ),
    .fco(\u2_Display/lt89_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_20|u2_Display/lt89_19  (
    .a({\u2_Display/n2677 ,\u2_Display/n2678 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c19 ),
    .fco(\u2_Display/lt89_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_22|u2_Display/lt89_21  (
    .a({\u2_Display/n2675 ,\u2_Display/n2676 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c21 ),
    .fco(\u2_Display/lt89_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_24|u2_Display/lt89_23  (
    .a({\u2_Display/n2673 ,\u2_Display/n2674 }),
    .b(2'b10),
    .fci(\u2_Display/lt89_c23 ),
    .fco(\u2_Display/lt89_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_26|u2_Display/lt89_25  (
    .a({\u2_Display/n2671 ,\u2_Display/n2672 }),
    .b(2'b01),
    .fci(\u2_Display/lt89_c25 ),
    .fco(\u2_Display/lt89_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_28|u2_Display/lt89_27  (
    .a({\u2_Display/n2669 ,\u2_Display/n2670 }),
    .b(2'b01),
    .fci(\u2_Display/lt89_c27 ),
    .fco(\u2_Display/lt89_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_2|u2_Display/lt89_1  (
    .a({\u2_Display/n2695 ,\u2_Display/n2696 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c1 ),
    .fco(\u2_Display/lt89_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_30|u2_Display/lt89_29  (
    .a({\u2_Display/n2667 ,\u2_Display/n2668 }),
    .b(2'b10),
    .fci(\u2_Display/lt89_c29 ),
    .fco(\u2_Display/lt89_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_4|u2_Display/lt89_3  (
    .a({\u2_Display/n2693 ,\u2_Display/n2694 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c3 ),
    .fco(\u2_Display/lt89_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_6|u2_Display/lt89_5  (
    .a({\u2_Display/n2691 ,\u2_Display/n2692 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c5 ),
    .fco(\u2_Display/lt89_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_8|u2_Display/lt89_7  (
    .a({\u2_Display/n2689 ,\u2_Display/n2690 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c7 ),
    .fco(\u2_Display/lt89_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_cout|u2_Display/lt89_31  (
    .a({1'b0,\u2_Display/n2666 }),
    .b(2'b10),
    .fci(\u2_Display/lt89_c31 ),
    .f({\u2_Display/n2698 ,open_n114116}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_0|u2_Display/lt8_2_cin  (
    .a({lcd_xpos[0],1'b0}),
    .b({\u2_Display/j [0],open_n114122}),
    .fco(\u2_Display/lt8_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_10|u2_Display/lt8_2_9  (
    .a(lcd_xpos[10:9]),
    .b({\u2_Display/add6_2_co ,\u2_Display/n135 [2]}),
    .fci(\u2_Display/lt8_2_c9 ),
    .fco(\u2_Display/lt8_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_2|u2_Display/lt8_2_1  (
    .a(lcd_xpos[2:1]),
    .b(\u2_Display/j [2:1]),
    .fci(\u2_Display/lt8_2_c1 ),
    .fco(\u2_Display/lt8_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_4|u2_Display/lt8_2_3  (
    .a(lcd_xpos[4:3]),
    .b(\u2_Display/j [4:3]),
    .fci(\u2_Display/lt8_2_c3 ),
    .fco(\u2_Display/lt8_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_6|u2_Display/lt8_2_5  (
    .a(lcd_xpos[6:5]),
    .b(\u2_Display/j [6:5]),
    .fci(\u2_Display/lt8_2_c5 ),
    .fco(\u2_Display/lt8_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_8|u2_Display/lt8_2_7  (
    .a(lcd_xpos[8:7]),
    .b(\u2_Display/n135 [1:0]),
    .fci(\u2_Display/lt8_2_c7 ),
    .fco(\u2_Display/lt8_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_cout|u2_Display/lt8_2_11  (
    .a({1'b0,lcd_xpos[11]}),
    .b(2'b10),
    .fci(\u2_Display/lt8_2_c11 ),
    .f({\u2_Display/n136 ,open_n114286}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_0|u2_Display/lt90_cin  (
    .a({\u2_Display/n2732 ,1'b0}),
    .b({1'b0,open_n114292}),
    .fco(\u2_Display/lt90_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_10|u2_Display/lt90_9  (
    .a({\u2_Display/n2722 ,\u2_Display/n2723 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c9 ),
    .fco(\u2_Display/lt90_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_12|u2_Display/lt90_11  (
    .a({\u2_Display/n2720 ,\u2_Display/n2721 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c11 ),
    .fco(\u2_Display/lt90_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_14|u2_Display/lt90_13  (
    .a({\u2_Display/n2718 ,\u2_Display/n2719 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c13 ),
    .fco(\u2_Display/lt90_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_16|u2_Display/lt90_15  (
    .a({\u2_Display/n2716 ,\u2_Display/n2717 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c15 ),
    .fco(\u2_Display/lt90_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_18|u2_Display/lt90_17  (
    .a({\u2_Display/n2714 ,\u2_Display/n2715 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c17 ),
    .fco(\u2_Display/lt90_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_20|u2_Display/lt90_19  (
    .a({\u2_Display/n2712 ,\u2_Display/n2713 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c19 ),
    .fco(\u2_Display/lt90_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_22|u2_Display/lt90_21  (
    .a({\u2_Display/n2710 ,\u2_Display/n2711 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c21 ),
    .fco(\u2_Display/lt90_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_24|u2_Display/lt90_23  (
    .a({\u2_Display/n2708 ,\u2_Display/n2709 }),
    .b(2'b11),
    .fci(\u2_Display/lt90_c23 ),
    .fco(\u2_Display/lt90_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_26|u2_Display/lt90_25  (
    .a({\u2_Display/n2706 ,\u2_Display/n2707 }),
    .b(2'b10),
    .fci(\u2_Display/lt90_c25 ),
    .fco(\u2_Display/lt90_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_28|u2_Display/lt90_27  (
    .a({\u2_Display/n2704 ,\u2_Display/n2705 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c27 ),
    .fco(\u2_Display/lt90_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_2|u2_Display/lt90_1  (
    .a({\u2_Display/n2730 ,\u2_Display/n2731 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c1 ),
    .fco(\u2_Display/lt90_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_30|u2_Display/lt90_29  (
    .a({\u2_Display/n2702 ,\u2_Display/n2703 }),
    .b(2'b01),
    .fci(\u2_Display/lt90_c29 ),
    .fco(\u2_Display/lt90_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_4|u2_Display/lt90_3  (
    .a({\u2_Display/n2728 ,\u2_Display/n2729 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c3 ),
    .fco(\u2_Display/lt90_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_6|u2_Display/lt90_5  (
    .a({\u2_Display/n2726 ,\u2_Display/n2727 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c5 ),
    .fco(\u2_Display/lt90_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_8|u2_Display/lt90_7  (
    .a({\u2_Display/n2724 ,\u2_Display/n2725 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c7 ),
    .fco(\u2_Display/lt90_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_cout|u2_Display/lt90_31  (
    .a({1'b0,\u2_Display/n2701 }),
    .b(2'b10),
    .fci(\u2_Display/lt90_c31 ),
    .f({\u2_Display/n2733 ,open_n114696}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_0|u2_Display/lt91_cin  (
    .a({\u2_Display/n2767 ,1'b0}),
    .b({1'b0,open_n114702}),
    .fco(\u2_Display/lt91_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_10|u2_Display/lt91_9  (
    .a({\u2_Display/n2757 ,\u2_Display/n2758 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c9 ),
    .fco(\u2_Display/lt91_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_12|u2_Display/lt91_11  (
    .a({\u2_Display/n2755 ,\u2_Display/n2756 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c11 ),
    .fco(\u2_Display/lt91_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_14|u2_Display/lt91_13  (
    .a({\u2_Display/n2753 ,\u2_Display/n2754 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c13 ),
    .fco(\u2_Display/lt91_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_16|u2_Display/lt91_15  (
    .a({\u2_Display/n2751 ,\u2_Display/n2752 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c15 ),
    .fco(\u2_Display/lt91_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_18|u2_Display/lt91_17  (
    .a({\u2_Display/n2749 ,\u2_Display/n2750 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c17 ),
    .fco(\u2_Display/lt91_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_20|u2_Display/lt91_19  (
    .a({\u2_Display/n2747 ,\u2_Display/n2748 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c19 ),
    .fco(\u2_Display/lt91_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_22|u2_Display/lt91_21  (
    .a({\u2_Display/n2745 ,\u2_Display/n2746 }),
    .b(2'b10),
    .fci(\u2_Display/lt91_c21 ),
    .fco(\u2_Display/lt91_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_24|u2_Display/lt91_23  (
    .a({\u2_Display/n2743 ,\u2_Display/n2744 }),
    .b(2'b01),
    .fci(\u2_Display/lt91_c23 ),
    .fco(\u2_Display/lt91_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_26|u2_Display/lt91_25  (
    .a({\u2_Display/n2741 ,\u2_Display/n2742 }),
    .b(2'b01),
    .fci(\u2_Display/lt91_c25 ),
    .fco(\u2_Display/lt91_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_28|u2_Display/lt91_27  (
    .a({\u2_Display/n2739 ,\u2_Display/n2740 }),
    .b(2'b10),
    .fci(\u2_Display/lt91_c27 ),
    .fco(\u2_Display/lt91_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_2|u2_Display/lt91_1  (
    .a({\u2_Display/n2765 ,\u2_Display/n2766 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c1 ),
    .fco(\u2_Display/lt91_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_30|u2_Display/lt91_29  (
    .a({\u2_Display/n2737 ,\u2_Display/n2738 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c29 ),
    .fco(\u2_Display/lt91_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_4|u2_Display/lt91_3  (
    .a({\u2_Display/n2763 ,\u2_Display/n2764 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c3 ),
    .fco(\u2_Display/lt91_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_6|u2_Display/lt91_5  (
    .a({\u2_Display/n2761 ,\u2_Display/n2762 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c5 ),
    .fco(\u2_Display/lt91_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_8|u2_Display/lt91_7  (
    .a({\u2_Display/n2759 ,\u2_Display/n2760 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c7 ),
    .fco(\u2_Display/lt91_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_cout|u2_Display/lt91_31  (
    .a({1'b0,\u2_Display/n2736 }),
    .b(2'b10),
    .fci(\u2_Display/lt91_c31 ),
    .f({\u2_Display/n2768 ,open_n115106}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_0|u2_Display/lt92_cin  (
    .a({\u2_Display/n2802 ,1'b0}),
    .b({1'b0,open_n115112}),
    .fco(\u2_Display/lt92_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_10|u2_Display/lt92_9  (
    .a({\u2_Display/n2792 ,\u2_Display/n2793 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c9 ),
    .fco(\u2_Display/lt92_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_12|u2_Display/lt92_11  (
    .a({\u2_Display/n2790 ,\u2_Display/n2791 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c11 ),
    .fco(\u2_Display/lt92_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_14|u2_Display/lt92_13  (
    .a({\u2_Display/n2788 ,\u2_Display/n2789 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c13 ),
    .fco(\u2_Display/lt92_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_16|u2_Display/lt92_15  (
    .a({\u2_Display/n2786 ,\u2_Display/n2787 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c15 ),
    .fco(\u2_Display/lt92_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_18|u2_Display/lt92_17  (
    .a({\u2_Display/n2784 ,\u2_Display/n2785 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c17 ),
    .fco(\u2_Display/lt92_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_20|u2_Display/lt92_19  (
    .a({\u2_Display/n2782 ,\u2_Display/n2783 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c19 ),
    .fco(\u2_Display/lt92_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_22|u2_Display/lt92_21  (
    .a({\u2_Display/n2780 ,\u2_Display/n2781 }),
    .b(2'b11),
    .fci(\u2_Display/lt92_c21 ),
    .fco(\u2_Display/lt92_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_24|u2_Display/lt92_23  (
    .a({\u2_Display/n2778 ,\u2_Display/n2779 }),
    .b(2'b10),
    .fci(\u2_Display/lt92_c23 ),
    .fco(\u2_Display/lt92_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_26|u2_Display/lt92_25  (
    .a({\u2_Display/n2776 ,\u2_Display/n2777 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c25 ),
    .fco(\u2_Display/lt92_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_28|u2_Display/lt92_27  (
    .a({\u2_Display/n2774 ,\u2_Display/n2775 }),
    .b(2'b01),
    .fci(\u2_Display/lt92_c27 ),
    .fco(\u2_Display/lt92_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_2|u2_Display/lt92_1  (
    .a({\u2_Display/n2800 ,\u2_Display/n2801 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c1 ),
    .fco(\u2_Display/lt92_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_30|u2_Display/lt92_29  (
    .a({\u2_Display/n2772 ,\u2_Display/n2773 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c29 ),
    .fco(\u2_Display/lt92_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_4|u2_Display/lt92_3  (
    .a({\u2_Display/n2798 ,\u2_Display/n2799 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c3 ),
    .fco(\u2_Display/lt92_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_6|u2_Display/lt92_5  (
    .a({\u2_Display/n2796 ,\u2_Display/n2797 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c5 ),
    .fco(\u2_Display/lt92_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_8|u2_Display/lt92_7  (
    .a({\u2_Display/n2794 ,\u2_Display/n2795 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c7 ),
    .fco(\u2_Display/lt92_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_cout|u2_Display/lt92_31  (
    .a({1'b0,\u2_Display/n2771 }),
    .b(2'b10),
    .fci(\u2_Display/lt92_c31 ),
    .f({\u2_Display/n2803 ,open_n115516}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_0|u2_Display/lt93_cin  (
    .a({\u2_Display/n2837 ,1'b0}),
    .b({1'b0,open_n115522}),
    .fco(\u2_Display/lt93_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_10|u2_Display/lt93_9  (
    .a({\u2_Display/n2827 ,\u2_Display/n2828 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c9 ),
    .fco(\u2_Display/lt93_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_12|u2_Display/lt93_11  (
    .a({\u2_Display/n2825 ,\u2_Display/n2826 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c11 ),
    .fco(\u2_Display/lt93_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_14|u2_Display/lt93_13  (
    .a({\u2_Display/n2823 ,\u2_Display/n2824 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c13 ),
    .fco(\u2_Display/lt93_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_16|u2_Display/lt93_15  (
    .a({\u2_Display/n2821 ,\u2_Display/n2822 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c15 ),
    .fco(\u2_Display/lt93_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_18|u2_Display/lt93_17  (
    .a({\u2_Display/n2819 ,\u2_Display/n2820 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c17 ),
    .fco(\u2_Display/lt93_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_20|u2_Display/lt93_19  (
    .a({\u2_Display/n2817 ,\u2_Display/n2818 }),
    .b(2'b10),
    .fci(\u2_Display/lt93_c19 ),
    .fco(\u2_Display/lt93_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_22|u2_Display/lt93_21  (
    .a({\u2_Display/n2815 ,\u2_Display/n2816 }),
    .b(2'b01),
    .fci(\u2_Display/lt93_c21 ),
    .fco(\u2_Display/lt93_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_24|u2_Display/lt93_23  (
    .a({\u2_Display/n2813 ,\u2_Display/n2814 }),
    .b(2'b01),
    .fci(\u2_Display/lt93_c23 ),
    .fco(\u2_Display/lt93_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_26|u2_Display/lt93_25  (
    .a({\u2_Display/n2811 ,\u2_Display/n2812 }),
    .b(2'b10),
    .fci(\u2_Display/lt93_c25 ),
    .fco(\u2_Display/lt93_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_28|u2_Display/lt93_27  (
    .a({\u2_Display/n2809 ,\u2_Display/n2810 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c27 ),
    .fco(\u2_Display/lt93_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_2|u2_Display/lt93_1  (
    .a({\u2_Display/n2835 ,\u2_Display/n2836 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c1 ),
    .fco(\u2_Display/lt93_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_30|u2_Display/lt93_29  (
    .a({\u2_Display/n2807 ,\u2_Display/n2808 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c29 ),
    .fco(\u2_Display/lt93_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_4|u2_Display/lt93_3  (
    .a({\u2_Display/n2833 ,\u2_Display/n2834 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c3 ),
    .fco(\u2_Display/lt93_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_6|u2_Display/lt93_5  (
    .a({\u2_Display/n2831 ,\u2_Display/n2832 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c5 ),
    .fco(\u2_Display/lt93_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_8|u2_Display/lt93_7  (
    .a({\u2_Display/n2829 ,\u2_Display/n2830 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c7 ),
    .fco(\u2_Display/lt93_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_cout|u2_Display/lt93_31  (
    .a({1'b0,\u2_Display/n2806 }),
    .b(2'b10),
    .fci(\u2_Display/lt93_c31 ),
    .f({\u2_Display/n2838 ,open_n115926}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_0|u2_Display/lt94_cin  (
    .a({\u2_Display/n2872 ,1'b0}),
    .b({1'b0,open_n115932}),
    .fco(\u2_Display/lt94_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_10|u2_Display/lt94_9  (
    .a({\u2_Display/n2862 ,\u2_Display/n2863 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c9 ),
    .fco(\u2_Display/lt94_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_12|u2_Display/lt94_11  (
    .a({\u2_Display/n2860 ,\u2_Display/n2861 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c11 ),
    .fco(\u2_Display/lt94_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_14|u2_Display/lt94_13  (
    .a({\u2_Display/n2858 ,\u2_Display/n2859 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c13 ),
    .fco(\u2_Display/lt94_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_16|u2_Display/lt94_15  (
    .a({\u2_Display/n2856 ,\u2_Display/n2857 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c15 ),
    .fco(\u2_Display/lt94_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_18|u2_Display/lt94_17  (
    .a({\u2_Display/n2854 ,\u2_Display/n2855 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c17 ),
    .fco(\u2_Display/lt94_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_20|u2_Display/lt94_19  (
    .a({\u2_Display/n2852 ,\u2_Display/n2853 }),
    .b(2'b11),
    .fci(\u2_Display/lt94_c19 ),
    .fco(\u2_Display/lt94_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_22|u2_Display/lt94_21  (
    .a({\u2_Display/n2850 ,\u2_Display/n2851 }),
    .b(2'b10),
    .fci(\u2_Display/lt94_c21 ),
    .fco(\u2_Display/lt94_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_24|u2_Display/lt94_23  (
    .a({\u2_Display/n2848 ,\u2_Display/n2849 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c23 ),
    .fco(\u2_Display/lt94_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_26|u2_Display/lt94_25  (
    .a({\u2_Display/n2846 ,\u2_Display/n2847 }),
    .b(2'b01),
    .fci(\u2_Display/lt94_c25 ),
    .fco(\u2_Display/lt94_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_28|u2_Display/lt94_27  (
    .a({\u2_Display/n2844 ,\u2_Display/n2845 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c27 ),
    .fco(\u2_Display/lt94_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_2|u2_Display/lt94_1  (
    .a({\u2_Display/n2870 ,\u2_Display/n2871 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c1 ),
    .fco(\u2_Display/lt94_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_30|u2_Display/lt94_29  (
    .a({\u2_Display/n2842 ,\u2_Display/n2843 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c29 ),
    .fco(\u2_Display/lt94_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_4|u2_Display/lt94_3  (
    .a({\u2_Display/n2868 ,\u2_Display/n2869 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c3 ),
    .fco(\u2_Display/lt94_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_6|u2_Display/lt94_5  (
    .a({\u2_Display/n2866 ,\u2_Display/n2867 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c5 ),
    .fco(\u2_Display/lt94_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_8|u2_Display/lt94_7  (
    .a({\u2_Display/n2864 ,\u2_Display/n2865 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c7 ),
    .fco(\u2_Display/lt94_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_cout|u2_Display/lt94_31  (
    .a({1'b0,\u2_Display/n2841 }),
    .b(2'b10),
    .fci(\u2_Display/lt94_c31 ),
    .f({\u2_Display/n2873 ,open_n116336}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_0|u2_Display/lt95_cin  (
    .a({\u2_Display/n2907 ,1'b0}),
    .b({1'b0,open_n116342}),
    .fco(\u2_Display/lt95_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_10|u2_Display/lt95_9  (
    .a({\u2_Display/n2897 ,\u2_Display/n2898 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c9 ),
    .fco(\u2_Display/lt95_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_12|u2_Display/lt95_11  (
    .a({\u2_Display/n2895 ,\u2_Display/n2896 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c11 ),
    .fco(\u2_Display/lt95_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_14|u2_Display/lt95_13  (
    .a({\u2_Display/n2893 ,\u2_Display/n2894 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c13 ),
    .fco(\u2_Display/lt95_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_16|u2_Display/lt95_15  (
    .a({\u2_Display/n2891 ,\u2_Display/n2892 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c15 ),
    .fco(\u2_Display/lt95_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_18|u2_Display/lt95_17  (
    .a({\u2_Display/n2889 ,\u2_Display/n2890 }),
    .b(2'b10),
    .fci(\u2_Display/lt95_c17 ),
    .fco(\u2_Display/lt95_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_20|u2_Display/lt95_19  (
    .a({\u2_Display/n2887 ,\u2_Display/n2888 }),
    .b(2'b01),
    .fci(\u2_Display/lt95_c19 ),
    .fco(\u2_Display/lt95_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_22|u2_Display/lt95_21  (
    .a({\u2_Display/n2885 ,\u2_Display/n2886 }),
    .b(2'b01),
    .fci(\u2_Display/lt95_c21 ),
    .fco(\u2_Display/lt95_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_24|u2_Display/lt95_23  (
    .a({\u2_Display/n2883 ,\u2_Display/n2884 }),
    .b(2'b10),
    .fci(\u2_Display/lt95_c23 ),
    .fco(\u2_Display/lt95_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_26|u2_Display/lt95_25  (
    .a({\u2_Display/n2881 ,\u2_Display/n2882 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c25 ),
    .fco(\u2_Display/lt95_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_28|u2_Display/lt95_27  (
    .a({\u2_Display/n2879 ,\u2_Display/n2880 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c27 ),
    .fco(\u2_Display/lt95_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_2|u2_Display/lt95_1  (
    .a({\u2_Display/n2905 ,\u2_Display/n2906 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c1 ),
    .fco(\u2_Display/lt95_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_30|u2_Display/lt95_29  (
    .a({\u2_Display/n2877 ,\u2_Display/n2878 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c29 ),
    .fco(\u2_Display/lt95_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_4|u2_Display/lt95_3  (
    .a({\u2_Display/n2903 ,\u2_Display/n2904 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c3 ),
    .fco(\u2_Display/lt95_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_6|u2_Display/lt95_5  (
    .a({\u2_Display/n2901 ,\u2_Display/n2902 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c5 ),
    .fco(\u2_Display/lt95_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_8|u2_Display/lt95_7  (
    .a({\u2_Display/n2899 ,\u2_Display/n2900 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c7 ),
    .fco(\u2_Display/lt95_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_cout|u2_Display/lt95_31  (
    .a({1'b0,\u2_Display/n2876 }),
    .b(2'b10),
    .fci(\u2_Display/lt95_c31 ),
    .f({\u2_Display/n2908 ,open_n116746}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_0|u2_Display/lt96_cin  (
    .a({\u2_Display/n2942 ,1'b0}),
    .b({1'b0,open_n116752}),
    .fco(\u2_Display/lt96_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_10|u2_Display/lt96_9  (
    .a({\u2_Display/n2932 ,\u2_Display/n2933 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c9 ),
    .fco(\u2_Display/lt96_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_12|u2_Display/lt96_11  (
    .a({\u2_Display/n2930 ,\u2_Display/n2931 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c11 ),
    .fco(\u2_Display/lt96_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_14|u2_Display/lt96_13  (
    .a({\u2_Display/n2928 ,\u2_Display/n2929 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c13 ),
    .fco(\u2_Display/lt96_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_16|u2_Display/lt96_15  (
    .a({\u2_Display/n2926 ,\u2_Display/n2927 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c15 ),
    .fco(\u2_Display/lt96_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_18|u2_Display/lt96_17  (
    .a({\u2_Display/n2924 ,\u2_Display/n2925 }),
    .b(2'b11),
    .fci(\u2_Display/lt96_c17 ),
    .fco(\u2_Display/lt96_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_20|u2_Display/lt96_19  (
    .a({\u2_Display/n2922 ,\u2_Display/n2923 }),
    .b(2'b10),
    .fci(\u2_Display/lt96_c19 ),
    .fco(\u2_Display/lt96_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_22|u2_Display/lt96_21  (
    .a({\u2_Display/n2920 ,\u2_Display/n2921 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c21 ),
    .fco(\u2_Display/lt96_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_24|u2_Display/lt96_23  (
    .a({\u2_Display/n2918 ,\u2_Display/n2919 }),
    .b(2'b01),
    .fci(\u2_Display/lt96_c23 ),
    .fco(\u2_Display/lt96_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_26|u2_Display/lt96_25  (
    .a({\u2_Display/n2916 ,\u2_Display/n2917 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c25 ),
    .fco(\u2_Display/lt96_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_28|u2_Display/lt96_27  (
    .a({\u2_Display/n2914 ,\u2_Display/n2915 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c27 ),
    .fco(\u2_Display/lt96_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_2|u2_Display/lt96_1  (
    .a({\u2_Display/n2940 ,\u2_Display/n2941 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c1 ),
    .fco(\u2_Display/lt96_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_30|u2_Display/lt96_29  (
    .a({\u2_Display/n2912 ,\u2_Display/n2913 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c29 ),
    .fco(\u2_Display/lt96_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_4|u2_Display/lt96_3  (
    .a({\u2_Display/n2938 ,\u2_Display/n2939 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c3 ),
    .fco(\u2_Display/lt96_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_6|u2_Display/lt96_5  (
    .a({\u2_Display/n2936 ,\u2_Display/n2937 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c5 ),
    .fco(\u2_Display/lt96_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_8|u2_Display/lt96_7  (
    .a({\u2_Display/n2934 ,\u2_Display/n2935 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c7 ),
    .fco(\u2_Display/lt96_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_cout|u2_Display/lt96_31  (
    .a({1'b0,\u2_Display/n2911 }),
    .b(2'b10),
    .fci(\u2_Display/lt96_c31 ),
    .f({\u2_Display/n2943 ,open_n117156}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_0|u2_Display/lt97_cin  (
    .a({\u2_Display/n2977 ,1'b0}),
    .b({1'b0,open_n117162}),
    .fco(\u2_Display/lt97_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_10|u2_Display/lt97_9  (
    .a({\u2_Display/n2967 ,\u2_Display/n2968 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c9 ),
    .fco(\u2_Display/lt97_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_12|u2_Display/lt97_11  (
    .a({\u2_Display/n2965 ,\u2_Display/n2966 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c11 ),
    .fco(\u2_Display/lt97_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_14|u2_Display/lt97_13  (
    .a({\u2_Display/n2963 ,\u2_Display/n2964 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c13 ),
    .fco(\u2_Display/lt97_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_16|u2_Display/lt97_15  (
    .a({\u2_Display/n2961 ,\u2_Display/n2962 }),
    .b(2'b10),
    .fci(\u2_Display/lt97_c15 ),
    .fco(\u2_Display/lt97_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_18|u2_Display/lt97_17  (
    .a({\u2_Display/n2959 ,\u2_Display/n2960 }),
    .b(2'b01),
    .fci(\u2_Display/lt97_c17 ),
    .fco(\u2_Display/lt97_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_20|u2_Display/lt97_19  (
    .a({\u2_Display/n2957 ,\u2_Display/n2958 }),
    .b(2'b01),
    .fci(\u2_Display/lt97_c19 ),
    .fco(\u2_Display/lt97_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_22|u2_Display/lt97_21  (
    .a({\u2_Display/n2955 ,\u2_Display/n2956 }),
    .b(2'b10),
    .fci(\u2_Display/lt97_c21 ),
    .fco(\u2_Display/lt97_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_24|u2_Display/lt97_23  (
    .a({\u2_Display/n2953 ,\u2_Display/n2954 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c23 ),
    .fco(\u2_Display/lt97_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_26|u2_Display/lt97_25  (
    .a({\u2_Display/n2951 ,\u2_Display/n2952 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c25 ),
    .fco(\u2_Display/lt97_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_28|u2_Display/lt97_27  (
    .a({\u2_Display/n2949 ,\u2_Display/n2950 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c27 ),
    .fco(\u2_Display/lt97_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_2|u2_Display/lt97_1  (
    .a({\u2_Display/n2975 ,\u2_Display/n2976 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c1 ),
    .fco(\u2_Display/lt97_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_30|u2_Display/lt97_29  (
    .a({\u2_Display/n2947 ,\u2_Display/n2948 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c29 ),
    .fco(\u2_Display/lt97_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_4|u2_Display/lt97_3  (
    .a({\u2_Display/n2973 ,\u2_Display/n2974 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c3 ),
    .fco(\u2_Display/lt97_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_6|u2_Display/lt97_5  (
    .a({\u2_Display/n2971 ,\u2_Display/n2972 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c5 ),
    .fco(\u2_Display/lt97_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_8|u2_Display/lt97_7  (
    .a({\u2_Display/n2969 ,\u2_Display/n2970 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c7 ),
    .fco(\u2_Display/lt97_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_cout|u2_Display/lt97_31  (
    .a({1'b0,\u2_Display/n2946 }),
    .b(2'b10),
    .fci(\u2_Display/lt97_c31 ),
    .f({\u2_Display/n2978 ,open_n117566}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_0|u2_Display/lt98_cin  (
    .a({\u2_Display/n3012 ,1'b0}),
    .b({1'b0,open_n117572}),
    .fco(\u2_Display/lt98_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_10|u2_Display/lt98_9  (
    .a({\u2_Display/n3002 ,\u2_Display/n3003 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c9 ),
    .fco(\u2_Display/lt98_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_12|u2_Display/lt98_11  (
    .a({\u2_Display/n3000 ,\u2_Display/n3001 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c11 ),
    .fco(\u2_Display/lt98_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_14|u2_Display/lt98_13  (
    .a({\u2_Display/n2998 ,\u2_Display/n2999 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c13 ),
    .fco(\u2_Display/lt98_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_16|u2_Display/lt98_15  (
    .a({\u2_Display/n2996 ,\u2_Display/n2997 }),
    .b(2'b11),
    .fci(\u2_Display/lt98_c15 ),
    .fco(\u2_Display/lt98_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_18|u2_Display/lt98_17  (
    .a({\u2_Display/n2994 ,\u2_Display/n2995 }),
    .b(2'b10),
    .fci(\u2_Display/lt98_c17 ),
    .fco(\u2_Display/lt98_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_20|u2_Display/lt98_19  (
    .a({\u2_Display/n2992 ,\u2_Display/n2993 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c19 ),
    .fco(\u2_Display/lt98_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_22|u2_Display/lt98_21  (
    .a({\u2_Display/n2990 ,\u2_Display/n2991 }),
    .b(2'b01),
    .fci(\u2_Display/lt98_c21 ),
    .fco(\u2_Display/lt98_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_24|u2_Display/lt98_23  (
    .a({\u2_Display/n2988 ,\u2_Display/n2989 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c23 ),
    .fco(\u2_Display/lt98_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_26|u2_Display/lt98_25  (
    .a({\u2_Display/n2986 ,\u2_Display/n2987 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c25 ),
    .fco(\u2_Display/lt98_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_28|u2_Display/lt98_27  (
    .a({\u2_Display/n2984 ,\u2_Display/n2985 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c27 ),
    .fco(\u2_Display/lt98_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_2|u2_Display/lt98_1  (
    .a({\u2_Display/n3010 ,\u2_Display/n3011 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c1 ),
    .fco(\u2_Display/lt98_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_30|u2_Display/lt98_29  (
    .a({\u2_Display/n2982 ,\u2_Display/n2983 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c29 ),
    .fco(\u2_Display/lt98_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_4|u2_Display/lt98_3  (
    .a({\u2_Display/n3008 ,\u2_Display/n3009 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c3 ),
    .fco(\u2_Display/lt98_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_6|u2_Display/lt98_5  (
    .a({\u2_Display/n3006 ,\u2_Display/n3007 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c5 ),
    .fco(\u2_Display/lt98_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_8|u2_Display/lt98_7  (
    .a({\u2_Display/n3004 ,\u2_Display/n3005 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c7 ),
    .fco(\u2_Display/lt98_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_cout|u2_Display/lt98_31  (
    .a({1'b0,\u2_Display/n2981 }),
    .b(2'b10),
    .fci(\u2_Display/lt98_c31 ),
    .f({\u2_Display/n3013 ,open_n117976}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_0|u2_Display/lt99_cin  (
    .a({\u2_Display/n3047 ,1'b0}),
    .b({1'b0,open_n117982}),
    .fco(\u2_Display/lt99_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_10|u2_Display/lt99_9  (
    .a({\u2_Display/n3037 ,\u2_Display/n3038 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c9 ),
    .fco(\u2_Display/lt99_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_12|u2_Display/lt99_11  (
    .a({\u2_Display/n3035 ,\u2_Display/n3036 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c11 ),
    .fco(\u2_Display/lt99_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_14|u2_Display/lt99_13  (
    .a({\u2_Display/n3033 ,\u2_Display/n3034 }),
    .b(2'b10),
    .fci(\u2_Display/lt99_c13 ),
    .fco(\u2_Display/lt99_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_16|u2_Display/lt99_15  (
    .a({\u2_Display/n3031 ,\u2_Display/n3032 }),
    .b(2'b01),
    .fci(\u2_Display/lt99_c15 ),
    .fco(\u2_Display/lt99_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_18|u2_Display/lt99_17  (
    .a({\u2_Display/n3029 ,\u2_Display/n3030 }),
    .b(2'b01),
    .fci(\u2_Display/lt99_c17 ),
    .fco(\u2_Display/lt99_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_20|u2_Display/lt99_19  (
    .a({\u2_Display/n3027 ,\u2_Display/n3028 }),
    .b(2'b10),
    .fci(\u2_Display/lt99_c19 ),
    .fco(\u2_Display/lt99_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_22|u2_Display/lt99_21  (
    .a({\u2_Display/n3025 ,\u2_Display/n3026 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c21 ),
    .fco(\u2_Display/lt99_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_24|u2_Display/lt99_23  (
    .a({\u2_Display/n3023 ,\u2_Display/n3024 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c23 ),
    .fco(\u2_Display/lt99_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_26|u2_Display/lt99_25  (
    .a({\u2_Display/n3021 ,\u2_Display/n3022 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c25 ),
    .fco(\u2_Display/lt99_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_28|u2_Display/lt99_27  (
    .a({\u2_Display/n3019 ,\u2_Display/n3020 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c27 ),
    .fco(\u2_Display/lt99_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_2|u2_Display/lt99_1  (
    .a({\u2_Display/n3045 ,\u2_Display/n3046 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c1 ),
    .fco(\u2_Display/lt99_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_30|u2_Display/lt99_29  (
    .a({\u2_Display/n3017 ,\u2_Display/n3018 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c29 ),
    .fco(\u2_Display/lt99_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_4|u2_Display/lt99_3  (
    .a({\u2_Display/n3043 ,\u2_Display/n3044 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c3 ),
    .fco(\u2_Display/lt99_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_6|u2_Display/lt99_5  (
    .a({\u2_Display/n3041 ,\u2_Display/n3042 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c5 ),
    .fco(\u2_Display/lt99_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_8|u2_Display/lt99_7  (
    .a({\u2_Display/n3039 ,\u2_Display/n3040 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c7 ),
    .fco(\u2_Display/lt99_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_cout|u2_Display/lt99_31  (
    .a({1'b0,\u2_Display/n3016 }),
    .b(2'b10),
    .fci(\u2_Display/lt99_c31 ),
    .f({\u2_Display/n3048 ,open_n118386}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_0|u2_Display/lt9_2_cin  (
    .a({\u2_Display/n137 [0],1'b0}),
    .b({lcd_xpos[0],open_n118392}),
    .fco(\u2_Display/lt9_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_10|u2_Display/lt9_2_9  (
    .a({\u2_Display/n137 [31],\u2_Display/n137 [9]}),
    .b(lcd_xpos[10:9]),
    .fci(\u2_Display/lt9_2_c9 ),
    .fco(\u2_Display/lt9_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_12|u2_Display/lt9_2_11  (
    .a({\u2_Display/n137 [31],\u2_Display/n137 [31]}),
    .b({1'b0,lcd_xpos[11]}),
    .fci(\u2_Display/lt9_2_c11 ),
    .fco(\u2_Display/lt9_2_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_2|u2_Display/lt9_2_1  (
    .a(\u2_Display/n137 [2:1]),
    .b(lcd_xpos[2:1]),
    .fci(\u2_Display/lt9_2_c1 ),
    .fco(\u2_Display/lt9_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_4|u2_Display/lt9_2_3  (
    .a(\u2_Display/n137 [4:3]),
    .b(lcd_xpos[4:3]),
    .fci(\u2_Display/lt9_2_c3 ),
    .fco(\u2_Display/lt9_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_6|u2_Display/lt9_2_5  (
    .a(\u2_Display/n137 [6:5]),
    .b(lcd_xpos[6:5]),
    .fci(\u2_Display/lt9_2_c5 ),
    .fco(\u2_Display/lt9_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_8|u2_Display/lt9_2_7  (
    .a(\u2_Display/n137 [8:7]),
    .b(lcd_xpos[8:7]),
    .fci(\u2_Display/lt9_2_c7 ),
    .fco(\u2_Display/lt9_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_cout_al_u5063  (
    .a({open_n118562,1'b0}),
    .b({open_n118563,1'b1}),
    .fci(\u2_Display/lt9_2_c13 ),
    .f({open_n118582,\u2_Display/n138 }));
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b0|u2_Display/reg0_b2  (
    .clk(clk_vga),
    .mi({\u2_Display/n37 [0],\u2_Display/n37 [2]}),
    .sr(\u2_Display/n35 ),
    .q({\u2_Display/n [0],\u2_Display/n [2]}));  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b1  (
    .clk(clk_vga),
    .mi({open_n118628,\u2_Display/n37 [1]}),
    .sr(\u2_Display/n35 ),
    .q({open_n118645,\u2_Display/n [1]}));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b10|u2_Display/reg0_b11  (
    .clk(clk_vga),
    .mi({\u2_Display/n37 [10],\u2_Display/n37 [11]}),
    .sr(\u2_Display/n35 ),
    .q({\u2_Display/n [10],\u2_Display/n [11]}));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b12|u2_Display/reg0_b15  (
    .clk(clk_vga),
    .mi({\u2_Display/n37 [12],\u2_Display/n37 [15]}),
    .sr(\u2_Display/n35 ),
    .q({\u2_Display/n [12],\u2_Display/n [15]}));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b13|u2_Display/reg0_b14  (
    .clk(clk_vga),
    .mi({\u2_Display/n37 [13],\u2_Display/n37 [14]}),
    .sr(\u2_Display/n35 ),
    .q({\u2_Display/n [13],\u2_Display/n [14]}));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b16|u2_Display/reg0_b21  (
    .clk(clk_vga),
    .mi({\u2_Display/n37 [16],\u2_Display/n37 [21]}),
    .sr(\u2_Display/n35 ),
    .q({\u2_Display/n [16],\u2_Display/n [21]}));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b17|u2_Display/reg0_b18  (
    .clk(clk_vga),
    .mi({\u2_Display/n37 [17],\u2_Display/n37 [18]}),
    .sr(\u2_Display/n35 ),
    .q({\u2_Display/n [17],\u2_Display/n [18]}));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b19|u2_Display/reg0_b24  (
    .clk(clk_vga),
    .mi({\u2_Display/n37 [19],\u2_Display/n37 [24]}),
    .sr(\u2_Display/n35 ),
    .q({\u2_Display/n [19],\u2_Display/n [24]}));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b20|u2_Display/reg0_b22  (
    .clk(clk_vga),
    .mi({\u2_Display/n37 [20],\u2_Display/n37 [22]}),
    .sr(\u2_Display/n35 ),
    .q({\u2_Display/n [20],\u2_Display/n [22]}));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b23|u2_Display/reg0_b25  (
    .clk(clk_vga),
    .mi({\u2_Display/n37 [23],\u2_Display/n37 [25]}),
    .sr(\u2_Display/n35 ),
    .q({\u2_Display/n [23],\u2_Display/n [25]}));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(C*D*B*A)"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(C*D*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b26|u2_Display/reg0_b3  (
    .a({_al_u1349_o,\u2_Display/n [2]}),
    .b({_al_u1350_o,\u2_Display/n [20]}),
    .c({_al_u1352_o,\u2_Display/n [21]}),
    .clk(clk_vga),
    .d({_al_u1351_o,\u2_Display/n [22]}),
    .mi({\u2_Display/n37 [26],\u2_Display/n37 [3]}),
    .sr(\u2_Display/n35 ),
    .f({_al_u1353_o,_al_u1351_o}),
    .q({\u2_Display/n [26],\u2_Display/n [3]}));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*C*D*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(B*C*D*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b27|u2_Display/reg0_b28  (
    .a({\u2_Display/n [16],_al_u1353_o}),
    .b({\u2_Display/n [17],_al_u1346_o}),
    .c({\u2_Display/n [18],_al_u1345_o}),
    .clk(clk_vga),
    .d({\u2_Display/n [19],_al_u1348_o}),
    .mi({\u2_Display/n37 [27],\u2_Display/n37 [28]}),
    .sr(\u2_Display/n35 ),
    .f({_al_u1352_o,\u2_Display/n35 }),
    .q({\u2_Display/n [27],\u2_Display/n [28]}));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(~D*~A*~C*~B)"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(~D*~A*~C*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b29|u2_Display/reg0_b30  (
    .a({\u2_Display/n [29],\u2_Display/n [23]}),
    .b({\u2_Display/n [27],\u2_Display/n [24]}),
    .c({\u2_Display/n [28],\u2_Display/n [25]}),
    .clk(clk_vga),
    .d({\u2_Display/n [3],\u2_Display/n [26]}),
    .mi({\u2_Display/n37 [29],\u2_Display/n37 [30]}),
    .sr(\u2_Display/n35 ),
    .f({_al_u1345_o,_al_u1346_o}),
    .q({\u2_Display/n [29],\u2_Display/n [30]}));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*~A)"),
    //.LUTF1("(~D*C*~B*~A)"),
    //.LUTG0("(~D*~C*B*~A)"),
    //.LUTG1("(~D*C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000100),
    .INIT_LUTF1(16'b0000000000010000),
    .INIT_LUTG0(16'b0000000000000100),
    .INIT_LUTG1(16'b0000000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b6|u2_Display/reg0_b9  (
    .a({\u2_Display/n [0],\u2_Display/n [30]}),
    .b({\u2_Display/n [1],\u2_Display/n [4]}),
    .c({\u2_Display/n [10],\u2_Display/n [5]}),
    .clk(clk_vga),
    .d({\u2_Display/n [11],\u2_Display/n [6]}),
    .mi({\u2_Display/n37 [6],\u2_Display/n37 [9]}),
    .sr(\u2_Display/n35 ),
    .f({_al_u1350_o,_al_u1347_o}),
    .q({\u2_Display/n [6],\u2_Display/n [9]}));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  // source/rtl/Display.v(61)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~C*B*~A)"),
    //.LUTF1("(C*A*~D*B)"),
    //.LUTG0("(~D*~C*B*~A)"),
    //.LUTG1("(C*A*~D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000100),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000000000100),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b8|u2_Display/reg0_b7  (
    .a({\u2_Display/n [8],\u2_Display/n [12]}),
    .b({_al_u1347_o,\u2_Display/n [13]}),
    .c({\u2_Display/n [9],\u2_Display/n [14]}),
    .clk(clk_vga),
    .d({\u2_Display/n [7],\u2_Display/n [15]}),
    .mi(\u2_Display/n37 [8:7]),
    .sr(\u2_Display/n35 ),
    .f({_al_u1348_o,_al_u1349_o}),
    .q(\u2_Display/n [8:7]));  // source/rtl/Display.v(61)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b0|u2_Display/reg2_b2  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [23],\u2_Display/counta [27]}),
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({\u2_Display/n1542 [23],\u2_Display/n1542 [27]}),
    .mi({\u2_Display/n41 [0],\u2_Display/n41 [2]}),
    .f({\u2_Display/n1551 ,\u2_Display/n1547 }),
    .q({\u2_Display/counta [0],\u2_Display/counta [2]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b10|u2_Display/reg2_b13  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .mi({\u2_Display/n41 [10],\u2_Display/n41 [13]}),
    .q({\u2_Display/counta [10],\u2_Display/counta [13]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b11|u2_Display/reg2_b17  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .mi({\u2_Display/n41 [11],\u2_Display/n41 [17]}),
    .q({\u2_Display/counta [11],\u2_Display/counta [17]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b12|u2_Display/reg2_b14  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .mi({\u2_Display/n41 [12],\u2_Display/n41 [14]}),
    .q({\u2_Display/counta [12],\u2_Display/counta [14]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b15|u2_Display/reg2_b21  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .mi({\u2_Display/n41 [15],\u2_Display/n41 [21]}),
    .q({\u2_Display/counta [15],\u2_Display/counta [21]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b16|u2_Display/reg2_b18  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .mi({\u2_Display/n41 [16],\u2_Display/n41 [18]}),
    .q({\u2_Display/counta [16],\u2_Display/counta [18]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b19|u2_Display/reg2_b25  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .mi({\u2_Display/n41 [19],\u2_Display/n41 [25]}),
    .q({\u2_Display/counta [19],\u2_Display/counta [25]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b1|u2_Display/reg2_b4  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [28],\u2_Display/counta [29]}),
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({\u2_Display/n1542 [28],\u2_Display/n1542 [29]}),
    .mi({\u2_Display/n41 [1],\u2_Display/n41 [4]}),
    .f({\u2_Display/n1546 ,\u2_Display/n1545 }),
    .q({\u2_Display/counta [1],\u2_Display/counta [4]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b20|u2_Display/reg2_b22  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .mi({\u2_Display/n41 [20],\u2_Display/n41 [22]}),
    .q({\u2_Display/counta [20],\u2_Display/counta [22]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b23|u2_Display/reg2_b28  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .mi({\u2_Display/n41 [23],\u2_Display/n41 [28]}),
    .q({\u2_Display/counta [23],\u2_Display/counta [28]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b24|u2_Display/reg2_b26  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .mi({\u2_Display/n41 [24],\u2_Display/n41 [26]}),
    .q({\u2_Display/counta [24],\u2_Display/counta [26]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b27|u2_Display/reg2_b29  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .mi({\u2_Display/n41 [27],\u2_Display/n41 [29]}),
    .q({\u2_Display/counta [27],\u2_Display/counta [29]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTF1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG0("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    //.LUTG1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111001111000000),
    .INIT_LUTG0(16'b1111001111000000),
    .INIT_LUTG1(16'b1111001111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b3|u2_Display/reg2_b9  (
    .b({\u2_Display/n1540 ,\u2_Display/n1540 }),
    .c({\u2_Display/counta [30],\u2_Display/counta [31]}),
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({\u2_Display/n1542 [30],\u2_Display/n1542 [31]}),
    .mi({\u2_Display/n41 [3],\u2_Display/n41 [9]}),
    .f({\u2_Display/n1544 ,\u2_Display/n1543 }),
    .q({\u2_Display/counta [3],\u2_Display/counta [9]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b7|u2_Display/reg2_b8  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s_gclk_net ),
    .mi({\u2_Display/n41 [7],\u2_Display/n41 [8]}),
    .q({\u2_Display/counta [7],\u2_Display/counta [8]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110011111100),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000110011111100),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b0|u2_Display/reg3_b8  (
    .b({_al_u3956_o,_al_u3991_o}),
    .c({\u2_Display/mux19_b0_sel_is_0_o ,\u2_Display/mux19_b0_sel_is_0_o }),
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({_al_u3958_o,_al_u3993_o}),
    .q({\u2_Display/i [0],\u2_Display/i [8]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~C*~A))"),
    //.LUTF1("~(B*~(C*~D))"),
    //.LUTG0("(B*~(D*~C*~A))"),
    //.LUTG1("~(B*~(C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100100011001100),
    .INIT_LUTF1(16'b0011001111110011),
    .INIT_LUTG0(16'b1100100011001100),
    .INIT_LUTG1(16'b0011001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b1|u2_Display/reg3_b5  (
    .a({open_n119352,_al_u3980_o}),
    .b({_al_u3963_o,_al_u3978_o}),
    .c({\u2_Display/mux19_b0_sel_is_0_o ,_al_u3981_o}),
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({_al_u3962_o,\u2_Display/mux19_b0_sel_is_0_o }),
    .q({\u2_Display/i [1],\u2_Display/i [5]}));  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C*~D))"),
    //.LUTG0("~(B*~(C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001111110011),
    .INIT_LUTG0(16'b0011001111110011),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b3  (
    .b({open_n119377,_al_u3972_o}),
    .c({open_n119378,\u2_Display/mux19_b0_sel_is_0_o }),
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({open_n119379,_al_u3971_o}),
    .q({open_n119402,\u2_Display/i [3]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*(~B*~(A)*~(0)+~B*A*~(0)+~(~B)*A*0+~B*A*0)))"),
    //.LUTF1("~(C*~(D*(~B*~(A)*~(0)+~B*A*~(0)+~(~B)*A*0+~B*A*0)))"),
    //.LUTG0("~(C*~(D*(~B*~(A)*~(1)+~B*A*~(1)+~(~B)*A*1+~B*A*1)))"),
    //.LUTG1("~(C*~(D*(~B*~(A)*~(1)+~B*A*~(1)+~(~B)*A*1+~B*A*1)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011111100001111),
    .INIT_LUTF1(16'b0011111100001111),
    .INIT_LUTG0(16'b1010111100001111),
    .INIT_LUTG1(16'b1010111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b4|u2_Display/reg3_b6  (
    .a({_al_u3974_o,_al_u3983_o}),
    .b({_al_u3975_o,_al_u3984_o}),
    .c({_al_u3976_o,_al_u3985_o}),
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({\u2_Display/mux19_b0_sel_is_0_o ,\u2_Display/mux19_b0_sel_is_0_o }),
    .e({on_off_pad[2],on_off_pad[2]}),
    .q({\u2_Display/i [4],\u2_Display/i [6]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTF1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG0("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    //.LUTG1("~(~B*~(D)*~(C)+~B*D*~(C)+~(~B)*D*C+~B*D*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110011111100),
    .INIT_LUTF1(16'b0000110011111100),
    .INIT_LUTG0(16'b0000110011111100),
    .INIT_LUTG1(16'b0000110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b7|u2_Display/reg3_b9  (
    .b({_al_u3987_o,_al_u3995_o}),
    .c({\u2_Display/mux19_b0_sel_is_0_o ,\u2_Display/mux19_b0_sel_is_0_o }),
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({_al_u3989_o,_al_u3997_o}),
    .q({\u2_Display/i [7],\u2_Display/i [9]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0011000011111100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0011000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b1|u2_Display/reg4_b2  (
    .b({\u2_Display/mux19_b0_sel_is_0_o ,\u2_Display/mux19_b0_sel_is_0_o }),
    .c({\u2_Display/counta [1],\u2_Display/counta [2]}),
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({_al_u3922_o,_al_u3926_o}),
    .q({\u2_Display/j [1],\u2_Display/j [2]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0011000011111100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0011000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b3|u2_Display/reg4_b6  (
    .b({\u2_Display/mux19_b0_sel_is_0_o ,\u2_Display/mux19_b0_sel_is_0_o }),
    .c({\u2_Display/counta [3],\u2_Display/counta [6]}),
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({_al_u3930_o,_al_u3942_o}),
    .q({\u2_Display/j [3],\u2_Display/j [6]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTF1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG0("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000011111100),
    .INIT_LUTF1(16'b0011000011111100),
    .INIT_LUTG0(16'b0011000011111100),
    .INIT_LUTG1(16'b0011000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b4|u2_Display/reg4_b5  (
    .b({\u2_Display/mux19_b0_sel_is_0_o ,\u2_Display/mux19_b0_sel_is_0_o }),
    .c({\u2_Display/counta [4],\u2_Display/counta [5]}),
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({_al_u3934_o,_al_u3938_o}),
    .q({\u2_Display/j [4],\u2_Display/j [5]}));  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTF1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    //.LUTG0("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    //.LUTG1("~(~C*~(D)*~(B)+~C*D*~(B)+~(~C)*D*B+~C*D*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0011000011111100),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b0011000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b7|u2_Display/reg4_b8  (
    .b({\u2_Display/mux19_b0_sel_is_0_o ,\u2_Display/mux19_b0_sel_is_0_o }),
    .c({\u2_Display/counta [7],\u2_Display/counta [8]}),
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s_gclk_net ),
    .d({_al_u3946_o,_al_u3950_o}),
    .q({\u2_Display/j [7],\u2_Display/j [8]}));  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub0_2/ucin_al_u5029"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub0_2/u3_al_u5030  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/i [5],\u2_Display/i [3]}),
    .e({\u2_Display/i [6],\u2_Display/i [4]}),
    .fci(\u2_Display/sub0_2/c3 ),
    .f({\u2_Display/n96 [5],\u2_Display/n96 [3]}),
    .fco(\u2_Display/sub0_2/c7 ),
    .fx({\u2_Display/n96 [6],\u2_Display/n96 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub0_2/ucin_al_u5029"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub0_2/u7_al_u5031  (
    .a(2'b11),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/i [9],\u2_Display/i [7]}),
    .e({\u2_Display/i [10],\u2_Display/i [8]}),
    .fci(\u2_Display/sub0_2/c7 ),
    .f({\u2_Display/n96 [9],\u2_Display/n96 [7]}),
    .fco(\u2_Display/sub0_2/c11 ),
    .fx({\u2_Display/n96 [10],\u2_Display/n96 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub0_2/ucin_al_u5029"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub0_2/ucin_al_u5029  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/i [1],1'b1}),
    .e({\u2_Display/i [2],\u2_Display/i [0]}),
    .f({\u2_Display/n96 [1],open_n119596}),
    .fco(\u2_Display/sub0_2/c3 ),
    .fx({\u2_Display/n96 [2],\u2_Display/n96 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub0_2/ucin_al_u5029"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub0_2/ucout_al_u5032  (
    .c(2'b11),
    .fci(\u2_Display/sub0_2/c11 ),
    .f({open_n119623,\u2_Display/n96 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub1_2/ucin_al_u5037"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub1_2/u3_al_u5038  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/j [5],\u2_Display/j [3]}),
    .e({\u2_Display/j [6],\u2_Display/j [4]}),
    .fci(\u2_Display/sub1_2/c3 ),
    .f({\u2_Display/n102 [5],\u2_Display/n102 [3]}),
    .fco(\u2_Display/sub1_2/c7 ),
    .fx({\u2_Display/n102 [6],\u2_Display/n102 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub1_2/ucin_al_u5037"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub1_2/u7_al_u5039  (
    .a(2'b10),
    .b({open_n119647,1'b0}),
    .c(2'b11),
    .d({\u2_Display/j [9],\u2_Display/j [7]}),
    .e({open_n119650,\u2_Display/j [8]}),
    .fci(\u2_Display/sub1_2/c7 ),
    .f({\u2_Display/n102 [9],\u2_Display/n102 [7]}),
    .fx({\u2_Display/n102 [31],\u2_Display/n102 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub1_2/ucin_al_u5037"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub1_2/ucin_al_u5037  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/j [1],1'b1}),
    .e({\u2_Display/j [2],\u2_Display/j [0]}),
    .f({\u2_Display/n102 [1],open_n119685}),
    .fco(\u2_Display/sub1_2/c3 ),
    .fx({\u2_Display/n102 [2],\u2_Display/n102 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub2_2/ucin_al_u5040"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub2_2/u3_al_u5041  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/j [5],\u2_Display/j [3]}),
    .e({\u2_Display/j [6],\u2_Display/j [4]}),
    .fci(\u2_Display/sub2_2/c3 ),
    .f({\u2_Display/n137 [5],\u2_Display/n137 [3]}),
    .fco(\u2_Display/sub2_2/c7 ),
    .fx({\u2_Display/n137 [6],\u2_Display/n137 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub2_2/ucin_al_u5040"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub2_2/u7_al_u5042  (
    .a(2'b11),
    .b({open_n119706,1'b0}),
    .c(2'b11),
    .d({\u2_Display/j [9],\u2_Display/j [7]}),
    .e({open_n119709,\u2_Display/j [8]}),
    .fci(\u2_Display/sub2_2/c7 ),
    .f({\u2_Display/n137 [9],\u2_Display/n137 [7]}),
    .fx({\u2_Display/n137 [31],\u2_Display/n137 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub2_2/ucin_al_u5040"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub2_2/ucin_al_u5040  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/j [1],1'b1}),
    .e({\u2_Display/j [2],\u2_Display/j [0]}),
    .f({\u2_Display/n137 [1],open_n119744}),
    .fco(\u2_Display/sub2_2/c3 ),
    .fx({\u2_Display/n137 [2],\u2_Display/n137 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub3_2/ucin_al_u5033"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub3_2/u3_al_u5034  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/i [5],\u2_Display/i [3]}),
    .e({\u2_Display/i [6],\u2_Display/i [4]}),
    .fci(\u2_Display/sub3_2/c3 ),
    .f({\u2_Display/n143 [5],\u2_Display/n143 [3]}),
    .fco(\u2_Display/sub3_2/c7 ),
    .fx({\u2_Display/n143 [6],\u2_Display/n143 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub3_2/ucin_al_u5033"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub3_2/u7_al_u5035  (
    .a(2'b10),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/i [9],\u2_Display/i [7]}),
    .e({\u2_Display/i [10],\u2_Display/i [8]}),
    .fci(\u2_Display/sub3_2/c7 ),
    .f({\u2_Display/n143 [9],\u2_Display/n143 [7]}),
    .fco(\u2_Display/sub3_2/c11 ),
    .fx({\u2_Display/n143 [10],\u2_Display/n143 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub3_2/ucin_al_u5033"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub3_2/ucin_al_u5033  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/i [1],1'b1}),
    .e({\u2_Display/i [2],\u2_Display/i [0]}),
    .f({\u2_Display/n143 [1],open_n119800}),
    .fco(\u2_Display/sub3_2/c3 ),
    .fx({\u2_Display/n143 [2],\u2_Display/n143 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub3_2/ucin_al_u5033"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub3_2/ucout_al_u5036  (
    .c(2'b11),
    .fci(\u2_Display/sub3_2/c11 ),
    .f({open_n119827,\u2_Display/n143 [31]}));

endmodule 

