// Verilog netlist created by TD v5.0.19080
// Sun May 31 12:04:53 2020

`timescale 1ns / 1ps
module VGA_Demo  // source/rtl/VGA_Demo.v(2)
  (
  clk_24m,
  on_off,
  rst_n,
  vga_b,
  vga_clk,
  vga_de,
  vga_g,
  vga_hs,
  vga_r,
  vga_vs
  );

  input clk_24m;  // source/rtl/VGA_Demo.v(4)
  input [7:0] on_off;  // source/rtl/VGA_Demo.v(6)
  input rst_n;  // source/rtl/VGA_Demo.v(5)
  output [7:0] vga_b;  // source/rtl/VGA_Demo.v(17)
  output vga_clk;  // source/rtl/VGA_Demo.v(9)
  output vga_de;  // source/rtl/VGA_Demo.v(13)
  output [7:0] vga_g;  // source/rtl/VGA_Demo.v(16)
  output vga_hs;  // source/rtl/VGA_Demo.v(10)
  output [7:0] vga_r;  // source/rtl/VGA_Demo.v(15)
  output vga_vs;  // source/rtl/VGA_Demo.v(11)

  wire [23:0] lcd_data;  // source/rtl/VGA_Demo.v(23)
  wire [11:0] lcd_xpos;  // source/rtl/VGA_Demo.v(21)
  wire [11:0] lcd_ypos;  // source/rtl/VGA_Demo.v(22)
  wire [7:0] on_off_pad;  // source/rtl/VGA_Demo.v(6)
  wire [11:0] \u1_Driver/hcnt ;  // source/rtl/Driver.v(44)
  wire [11:0] \u1_Driver/n2 ;
  wire [12:0] \u1_Driver/n20 ;
  wire [12:0] \u1_Driver/n21 ;
  wire [11:0] \u1_Driver/n3 ;
  wire [11:0] \u1_Driver/n7 ;
  wire [11:0] \u1_Driver/n8 ;
  wire [11:0] \u1_Driver/vcnt ;  // source/rtl/Driver.v(45)
  wire [31:0] \u2_Display/counta ;  // source/rtl/Display.v(39)
  wire [31:0] \u2_Display/i ;  // source/rtl/Display.v(41)
  wire [31:0] \u2_Display/j ;  // source/rtl/Display.v(42)
  wire [30:0] \u2_Display/n ;  // source/rtl/Display.v(48)
  wire [31:0] \u2_Display/n1014 ;
  wire [31:0] \u2_Display/n102 ;
  wire [31:0] \u2_Display/n1049 ;
  wire [31:0] \u2_Display/n1084 ;
  wire [31:0] \u2_Display/n1119 ;
  wire [31:0] \u2_Display/n1154 ;
  wire [31:0] \u2_Display/n1189 ;
  wire [24:0] \u2_Display/n135 ;
  wire [31:0] \u2_Display/n137 ;
  wire [22:0] \u2_Display/n140 ;
  wire [31:0] \u2_Display/n143 ;
  wire [31:0] \u2_Display/n1542 ;
  wire [31:0] \u2_Display/n1577 ;
  wire [31:0] \u2_Display/n1612 ;
  wire [31:0] \u2_Display/n1647 ;
  wire [31:0] \u2_Display/n1682 ;
  wire [31:0] \u2_Display/n1717 ;
  wire [31:0] \u2_Display/n1752 ;
  wire [31:0] \u2_Display/n1787 ;
  wire [31:0] \u2_Display/n1822 ;
  wire [31:0] \u2_Display/n1857 ;
  wire [31:0] \u2_Display/n1892 ;
  wire [31:0] \u2_Display/n1927 ;
  wire [31:0] \u2_Display/n1962 ;
  wire [31:0] \u2_Display/n1997 ;
  wire [31:0] \u2_Display/n2032 ;
  wire [31:0] \u2_Display/n2067 ;
  wire [31:0] \u2_Display/n2102 ;
  wire [31:0] \u2_Display/n2137 ;
  wire [31:0] \u2_Display/n2172 ;
  wire [31:0] \u2_Display/n2207 ;
  wire [31:0] \u2_Display/n2242 ;
  wire [31:0] \u2_Display/n2277 ;
  wire [31:0] \u2_Display/n2312 ;
  wire [23:0] \u2_Display/n236 ;
  wire [31:0] \u2_Display/n238 ;
  wire [31:0] \u2_Display/n239 ;
  wire [23:0] \u2_Display/n240 ;
  wire [31:0] \u2_Display/n2665 ;
  wire [31:0] \u2_Display/n2700 ;
  wire [31:0] \u2_Display/n2735 ;
  wire [31:0] \u2_Display/n2770 ;
  wire [31:0] \u2_Display/n2805 ;
  wire [31:0] \u2_Display/n2840 ;
  wire [31:0] \u2_Display/n2875 ;
  wire [31:0] \u2_Display/n2910 ;
  wire [31:0] \u2_Display/n2945 ;
  wire [31:0] \u2_Display/n2980 ;
  wire [31:0] \u2_Display/n3015 ;
  wire [31:0] \u2_Display/n3050 ;
  wire [31:0] \u2_Display/n3085 ;
  wire [31:0] \u2_Display/n3120 ;
  wire [31:0] \u2_Display/n3155 ;
  wire [31:0] \u2_Display/n3190 ;
  wire [31:0] \u2_Display/n3225 ;
  wire [31:0] \u2_Display/n3260 ;
  wire [31:0] \u2_Display/n3295 ;
  wire [31:0] \u2_Display/n3330 ;
  wire [31:0] \u2_Display/n3365 ;
  wire [31:0] \u2_Display/n3400 ;
  wire [31:0] \u2_Display/n3435 ;
  wire [30:0] \u2_Display/n37 ;
  wire [31:0] \u2_Display/n3788 ;
  wire [31:0] \u2_Display/n3823 ;
  wire [31:0] \u2_Display/n3858 ;
  wire [31:0] \u2_Display/n3893 ;
  wire [31:0] \u2_Display/n3928 ;
  wire [31:0] \u2_Display/n3963 ;
  wire [31:0] \u2_Display/n3998 ;
  wire [31:0] \u2_Display/n4033 ;
  wire [31:0] \u2_Display/n4068 ;
  wire [31:0] \u2_Display/n41 ;
  wire [31:0] \u2_Display/n4103 ;
  wire [31:0] \u2_Display/n4138 ;
  wire [31:0] \u2_Display/n4173 ;
  wire [31:0] \u2_Display/n419 ;
  wire [31:0] \u2_Display/n4208 ;
  wire [31:0] \u2_Display/n4243 ;
  wire [31:0] \u2_Display/n4278 ;
  wire [23:0] \u2_Display/n43 ;
  wire [31:0] \u2_Display/n4313 ;
  wire [31:0] \u2_Display/n4348 ;
  wire [31:0] \u2_Display/n4383 ;
  wire [31:0] \u2_Display/n4418 ;
  wire [31:0] \u2_Display/n4453 ;
  wire [31:0] \u2_Display/n4488 ;
  wire [31:0] \u2_Display/n4523 ;
  wire [31:0] \u2_Display/n454 ;
  wire [31:0] \u2_Display/n4558 ;
  wire [31:0] \u2_Display/n489 ;
  wire [31:0] \u2_Display/n4911 ;
  wire [31:0] \u2_Display/n4946 ;
  wire [31:0] \u2_Display/n4981 ;
  wire [31:0] \u2_Display/n5016 ;
  wire [31:0] \u2_Display/n5051 ;
  wire [31:0] \u2_Display/n5086 ;
  wire [31:0] \u2_Display/n5121 ;
  wire [31:0] \u2_Display/n5156 ;
  wire [31:0] \u2_Display/n5191 ;
  wire [31:0] \u2_Display/n5226 ;
  wire [31:0] \u2_Display/n524 ;
  wire [31:0] \u2_Display/n5261 ;
  wire [31:0] \u2_Display/n5296 ;
  wire [31:0] \u2_Display/n5331 ;
  wire [31:0] \u2_Display/n5366 ;
  wire [31:0] \u2_Display/n5401 ;
  wire [31:0] \u2_Display/n5436 ;
  wire [31:0] \u2_Display/n5471 ;
  wire [31:0] \u2_Display/n5506 ;
  wire [31:0] \u2_Display/n5541 ;
  wire [31:0] \u2_Display/n5576 ;
  wire [31:0] \u2_Display/n559 ;
  wire [31:0] \u2_Display/n5611 ;
  wire [31:0] \u2_Display/n5646 ;
  wire [31:0] \u2_Display/n5681 ;
  wire [31:0] \u2_Display/n594 ;
  wire [31:0] \u2_Display/n629 ;
  wire [31:0] \u2_Display/n664 ;
  wire [31:0] \u2_Display/n699 ;
  wire [31:0] \u2_Display/n734 ;
  wire [31:0] \u2_Display/n769 ;
  wire [31:0] \u2_Display/n804 ;
  wire [31:0] \u2_Display/n839 ;
  wire [31:0] \u2_Display/n874 ;
  wire [31:0] \u2_Display/n909 ;
  wire [24:0] \u2_Display/n94 ;
  wire [31:0] \u2_Display/n944 ;
  wire [31:0] \u2_Display/n96 ;
  wire [31:0] \u2_Display/n979 ;
  wire [22:0] \u2_Display/n99 ;
  wire [7:0] vga_b_pad;  // source/rtl/VGA_Demo.v(17)
  wire _al_u1168_o;
  wire _al_u1170_o;
  wire _al_u1171_o;
  wire _al_u1345_o;
  wire _al_u1346_o;
  wire _al_u1347_o;
  wire _al_u1348_o;
  wire _al_u1349_o;
  wire _al_u1350_o;
  wire _al_u1351_o;
  wire _al_u1352_o;
  wire _al_u1353_o;
  wire _al_u3916_o;
  wire _al_u3917_o;
  wire _al_u3918_o;
  wire _al_u3920_o;
  wire _al_u3921_o;
  wire _al_u3922_o;
  wire _al_u3924_o;
  wire _al_u3925_o;
  wire _al_u3926_o;
  wire _al_u3928_o;
  wire _al_u3929_o;
  wire _al_u3930_o;
  wire _al_u3932_o;
  wire _al_u3933_o;
  wire _al_u3934_o;
  wire _al_u3936_o;
  wire _al_u3937_o;
  wire _al_u3938_o;
  wire _al_u3940_o;
  wire _al_u3941_o;
  wire _al_u3942_o;
  wire _al_u3944_o;
  wire _al_u3945_o;
  wire _al_u3946_o;
  wire _al_u3948_o;
  wire _al_u3949_o;
  wire _al_u3950_o;
  wire _al_u3952_o;
  wire _al_u3953_o;
  wire _al_u3954_o;
  wire _al_u3956_o;
  wire _al_u3957_o;
  wire _al_u3958_o;
  wire _al_u3960_o;
  wire _al_u3961_o;
  wire _al_u3962_o;
  wire _al_u3963_o;
  wire _al_u3965_o;
  wire _al_u3966_o;
  wire _al_u3967_o;
  wire _al_u3969_o;
  wire _al_u3970_o;
  wire _al_u3971_o;
  wire _al_u3972_o;
  wire _al_u3974_o;
  wire _al_u3975_o;
  wire _al_u3976_o;
  wire _al_u3978_o;
  wire _al_u3979_o;
  wire _al_u3980_o;
  wire _al_u3981_o;
  wire _al_u3983_o;
  wire _al_u3984_o;
  wire _al_u3985_o;
  wire _al_u3987_o;
  wire _al_u3988_o;
  wire _al_u3989_o;
  wire _al_u3991_o;
  wire _al_u3992_o;
  wire _al_u3993_o;
  wire _al_u3995_o;
  wire _al_u3996_o;
  wire _al_u3997_o;
  wire _al_u997_o;
  wire _al_u998_o;
  wire clk_24m_pad;  // source/rtl/VGA_Demo.v(4)
  wire clk_vga;  // source/rtl/VGA_Demo.v(20)
  wire rst_n_pad;  // source/rtl/VGA_Demo.v(5)
  wire \u0_PLL/n0 ;
  wire \u0_PLL/uut/clk0_buf ;  // al_ip/PLL.v(32)
  wire \u1_Driver/add0/c11 ;
  wire \u1_Driver/add0/c3 ;
  wire \u1_Driver/add0/c7 ;
  wire \u1_Driver/add1/c11 ;
  wire \u1_Driver/add1/c3 ;
  wire \u1_Driver/add1/c7 ;
  wire \u1_Driver/lcd_request ;  // source/rtl/Driver.v(46)
  wire \u1_Driver/lt0_c1 ;
  wire \u1_Driver/lt0_c11 ;
  wire \u1_Driver/lt0_c3 ;
  wire \u1_Driver/lt0_c5 ;
  wire \u1_Driver/lt0_c7 ;
  wire \u1_Driver/lt0_c9 ;
  wire \u1_Driver/lt1_c1 ;
  wire \u1_Driver/lt1_c11 ;
  wire \u1_Driver/lt1_c3 ;
  wire \u1_Driver/lt1_c5 ;
  wire \u1_Driver/lt1_c7 ;
  wire \u1_Driver/lt1_c9 ;
  wire \u1_Driver/lt2_c1 ;
  wire \u1_Driver/lt2_c11 ;
  wire \u1_Driver/lt2_c3 ;
  wire \u1_Driver/lt2_c5 ;
  wire \u1_Driver/lt2_c7 ;
  wire \u1_Driver/lt2_c9 ;
  wire \u1_Driver/lt3_c1 ;
  wire \u1_Driver/lt3_c11 ;
  wire \u1_Driver/lt3_c3 ;
  wire \u1_Driver/lt3_c5 ;
  wire \u1_Driver/lt3_c7 ;
  wire \u1_Driver/lt3_c9 ;
  wire \u1_Driver/lt4_c1 ;
  wire \u1_Driver/lt4_c11 ;
  wire \u1_Driver/lt4_c3 ;
  wire \u1_Driver/lt4_c5 ;
  wire \u1_Driver/lt4_c7 ;
  wire \u1_Driver/lt4_c9 ;
  wire \u1_Driver/lt5_c1 ;
  wire \u1_Driver/lt5_c11 ;
  wire \u1_Driver/lt5_c3 ;
  wire \u1_Driver/lt5_c5 ;
  wire \u1_Driver/lt5_c7 ;
  wire \u1_Driver/lt5_c9 ;
  wire \u1_Driver/lt6_c1 ;
  wire \u1_Driver/lt6_c11 ;
  wire \u1_Driver/lt6_c3 ;
  wire \u1_Driver/lt6_c5 ;
  wire \u1_Driver/lt6_c7 ;
  wire \u1_Driver/lt6_c9 ;
  wire \u1_Driver/lt7_c1 ;
  wire \u1_Driver/lt7_c11 ;
  wire \u1_Driver/lt7_c3 ;
  wire \u1_Driver/lt7_c5 ;
  wire \u1_Driver/lt7_c7 ;
  wire \u1_Driver/lt7_c9 ;
  wire \u1_Driver/lt8_c1 ;
  wire \u1_Driver/lt8_c11 ;
  wire \u1_Driver/lt8_c3 ;
  wire \u1_Driver/lt8_c5 ;
  wire \u1_Driver/lt8_c7 ;
  wire \u1_Driver/lt8_c9 ;
  wire \u1_Driver/n1 ;
  wire \u1_Driver/n10 ;
  wire \u1_Driver/n11 ;
  wire \u1_Driver/n12 ;
  wire \u1_Driver/n14 ;
  wire \u1_Driver/n15 ;
  wire \u1_Driver/n17 ;
  wire \u1_Driver/n18 ;
  wire \u1_Driver/n4 ;
  wire \u1_Driver/n5 ;
  wire \u1_Driver/n6_lutinv ;
  wire \u1_Driver/sub0/c11 ;
  wire \u1_Driver/sub0/c3 ;
  wire \u1_Driver/sub0/c7 ;
  wire \u1_Driver/sub1/c11 ;
  wire \u1_Driver/sub1/c3 ;
  wire \u1_Driver/sub1/c7 ;
  wire \u2_Display/add0/c11 ;
  wire \u2_Display/add0/c15 ;
  wire \u2_Display/add0/c19 ;
  wire \u2_Display/add0/c23 ;
  wire \u2_Display/add0/c27 ;
  wire \u2_Display/add0/c3 ;
  wire \u2_Display/add0/c7 ;
  wire \u2_Display/add1/c11 ;
  wire \u2_Display/add1/c15 ;
  wire \u2_Display/add1/c19 ;
  wire \u2_Display/add1/c23 ;
  wire \u2_Display/add1/c27 ;
  wire \u2_Display/add1/c3 ;
  wire \u2_Display/add1/c31 ;
  wire \u2_Display/add1/c7 ;
  wire \u2_Display/add100/c11 ;
  wire \u2_Display/add100/c15 ;
  wire \u2_Display/add100/c19 ;
  wire \u2_Display/add100/c23 ;
  wire \u2_Display/add100/c27 ;
  wire \u2_Display/add100/c3 ;
  wire \u2_Display/add100/c31 ;
  wire \u2_Display/add100/c7 ;
  wire \u2_Display/add101/c11 ;
  wire \u2_Display/add101/c15 ;
  wire \u2_Display/add101/c19 ;
  wire \u2_Display/add101/c23 ;
  wire \u2_Display/add101/c27 ;
  wire \u2_Display/add101/c3 ;
  wire \u2_Display/add101/c31 ;
  wire \u2_Display/add101/c7 ;
  wire \u2_Display/add102/c11 ;
  wire \u2_Display/add102/c15 ;
  wire \u2_Display/add102/c19 ;
  wire \u2_Display/add102/c23 ;
  wire \u2_Display/add102/c27 ;
  wire \u2_Display/add102/c3 ;
  wire \u2_Display/add102/c31 ;
  wire \u2_Display/add102/c7 ;
  wire \u2_Display/add103/c11 ;
  wire \u2_Display/add103/c15 ;
  wire \u2_Display/add103/c19 ;
  wire \u2_Display/add103/c23 ;
  wire \u2_Display/add103/c27 ;
  wire \u2_Display/add103/c3 ;
  wire \u2_Display/add103/c31 ;
  wire \u2_Display/add103/c7 ;
  wire \u2_Display/add104/c11 ;
  wire \u2_Display/add104/c15 ;
  wire \u2_Display/add104/c19 ;
  wire \u2_Display/add104/c23 ;
  wire \u2_Display/add104/c27 ;
  wire \u2_Display/add104/c3 ;
  wire \u2_Display/add104/c31 ;
  wire \u2_Display/add104/c7 ;
  wire \u2_Display/add105/c11 ;
  wire \u2_Display/add105/c15 ;
  wire \u2_Display/add105/c19 ;
  wire \u2_Display/add105/c23 ;
  wire \u2_Display/add105/c27 ;
  wire \u2_Display/add105/c3 ;
  wire \u2_Display/add105/c31 ;
  wire \u2_Display/add105/c7 ;
  wire \u2_Display/add106/c3 ;
  wire \u2_Display/add106/c7 ;
  wire \u2_Display/add117/c11 ;
  wire \u2_Display/add117/c15 ;
  wire \u2_Display/add117/c19 ;
  wire \u2_Display/add117/c23 ;
  wire \u2_Display/add117/c27 ;
  wire \u2_Display/add117/c3 ;
  wire \u2_Display/add117/c31 ;
  wire \u2_Display/add117/c7 ;
  wire \u2_Display/add118/c11 ;
  wire \u2_Display/add118/c15 ;
  wire \u2_Display/add118/c19 ;
  wire \u2_Display/add118/c23 ;
  wire \u2_Display/add118/c27 ;
  wire \u2_Display/add118/c3 ;
  wire \u2_Display/add118/c31 ;
  wire \u2_Display/add118/c7 ;
  wire \u2_Display/add119/c11 ;
  wire \u2_Display/add119/c15 ;
  wire \u2_Display/add119/c19 ;
  wire \u2_Display/add119/c23 ;
  wire \u2_Display/add119/c27 ;
  wire \u2_Display/add119/c3 ;
  wire \u2_Display/add119/c31 ;
  wire \u2_Display/add119/c7 ;
  wire \u2_Display/add120/c11 ;
  wire \u2_Display/add120/c15 ;
  wire \u2_Display/add120/c19 ;
  wire \u2_Display/add120/c23 ;
  wire \u2_Display/add120/c27 ;
  wire \u2_Display/add120/c3 ;
  wire \u2_Display/add120/c31 ;
  wire \u2_Display/add120/c7 ;
  wire \u2_Display/add121/c11 ;
  wire \u2_Display/add121/c15 ;
  wire \u2_Display/add121/c19 ;
  wire \u2_Display/add121/c23 ;
  wire \u2_Display/add121/c27 ;
  wire \u2_Display/add121/c3 ;
  wire \u2_Display/add121/c31 ;
  wire \u2_Display/add121/c7 ;
  wire \u2_Display/add122/c11 ;
  wire \u2_Display/add122/c15 ;
  wire \u2_Display/add122/c19 ;
  wire \u2_Display/add122/c23 ;
  wire \u2_Display/add122/c27 ;
  wire \u2_Display/add122/c3 ;
  wire \u2_Display/add122/c31 ;
  wire \u2_Display/add122/c7 ;
  wire \u2_Display/add123/c11 ;
  wire \u2_Display/add123/c15 ;
  wire \u2_Display/add123/c19 ;
  wire \u2_Display/add123/c23 ;
  wire \u2_Display/add123/c27 ;
  wire \u2_Display/add123/c3 ;
  wire \u2_Display/add123/c31 ;
  wire \u2_Display/add123/c7 ;
  wire \u2_Display/add124/c11 ;
  wire \u2_Display/add124/c15 ;
  wire \u2_Display/add124/c19 ;
  wire \u2_Display/add124/c23 ;
  wire \u2_Display/add124/c27 ;
  wire \u2_Display/add124/c3 ;
  wire \u2_Display/add124/c31 ;
  wire \u2_Display/add124/c7 ;
  wire \u2_Display/add125/c11 ;
  wire \u2_Display/add125/c15 ;
  wire \u2_Display/add125/c19 ;
  wire \u2_Display/add125/c23 ;
  wire \u2_Display/add125/c27 ;
  wire \u2_Display/add125/c3 ;
  wire \u2_Display/add125/c31 ;
  wire \u2_Display/add125/c7 ;
  wire \u2_Display/add126/c11 ;
  wire \u2_Display/add126/c15 ;
  wire \u2_Display/add126/c19 ;
  wire \u2_Display/add126/c23 ;
  wire \u2_Display/add126/c27 ;
  wire \u2_Display/add126/c3 ;
  wire \u2_Display/add126/c31 ;
  wire \u2_Display/add126/c7 ;
  wire \u2_Display/add127/c11 ;
  wire \u2_Display/add127/c15 ;
  wire \u2_Display/add127/c19 ;
  wire \u2_Display/add127/c23 ;
  wire \u2_Display/add127/c27 ;
  wire \u2_Display/add127/c3 ;
  wire \u2_Display/add127/c31 ;
  wire \u2_Display/add127/c7 ;
  wire \u2_Display/add128/c11 ;
  wire \u2_Display/add128/c15 ;
  wire \u2_Display/add128/c19 ;
  wire \u2_Display/add128/c23 ;
  wire \u2_Display/add128/c27 ;
  wire \u2_Display/add128/c3 ;
  wire \u2_Display/add128/c31 ;
  wire \u2_Display/add128/c7 ;
  wire \u2_Display/add129/c11 ;
  wire \u2_Display/add129/c15 ;
  wire \u2_Display/add129/c19 ;
  wire \u2_Display/add129/c23 ;
  wire \u2_Display/add129/c27 ;
  wire \u2_Display/add129/c3 ;
  wire \u2_Display/add129/c31 ;
  wire \u2_Display/add129/c7 ;
  wire \u2_Display/add130/c11 ;
  wire \u2_Display/add130/c15 ;
  wire \u2_Display/add130/c19 ;
  wire \u2_Display/add130/c23 ;
  wire \u2_Display/add130/c27 ;
  wire \u2_Display/add130/c3 ;
  wire \u2_Display/add130/c31 ;
  wire \u2_Display/add130/c7 ;
  wire \u2_Display/add131/c11 ;
  wire \u2_Display/add131/c15 ;
  wire \u2_Display/add131/c19 ;
  wire \u2_Display/add131/c23 ;
  wire \u2_Display/add131/c27 ;
  wire \u2_Display/add131/c3 ;
  wire \u2_Display/add131/c31 ;
  wire \u2_Display/add131/c7 ;
  wire \u2_Display/add132/c11 ;
  wire \u2_Display/add132/c15 ;
  wire \u2_Display/add132/c19 ;
  wire \u2_Display/add132/c23 ;
  wire \u2_Display/add132/c27 ;
  wire \u2_Display/add132/c3 ;
  wire \u2_Display/add132/c31 ;
  wire \u2_Display/add132/c7 ;
  wire \u2_Display/add133/c11 ;
  wire \u2_Display/add133/c15 ;
  wire \u2_Display/add133/c19 ;
  wire \u2_Display/add133/c23 ;
  wire \u2_Display/add133/c27 ;
  wire \u2_Display/add133/c3 ;
  wire \u2_Display/add133/c31 ;
  wire \u2_Display/add133/c7 ;
  wire \u2_Display/add134/c11 ;
  wire \u2_Display/add134/c15 ;
  wire \u2_Display/add134/c19 ;
  wire \u2_Display/add134/c23 ;
  wire \u2_Display/add134/c27 ;
  wire \u2_Display/add134/c3 ;
  wire \u2_Display/add134/c31 ;
  wire \u2_Display/add134/c7 ;
  wire \u2_Display/add135/c11 ;
  wire \u2_Display/add135/c15 ;
  wire \u2_Display/add135/c19 ;
  wire \u2_Display/add135/c23 ;
  wire \u2_Display/add135/c27 ;
  wire \u2_Display/add135/c3 ;
  wire \u2_Display/add135/c31 ;
  wire \u2_Display/add135/c7 ;
  wire \u2_Display/add136/c11 ;
  wire \u2_Display/add136/c15 ;
  wire \u2_Display/add136/c19 ;
  wire \u2_Display/add136/c23 ;
  wire \u2_Display/add136/c27 ;
  wire \u2_Display/add136/c3 ;
  wire \u2_Display/add136/c31 ;
  wire \u2_Display/add136/c7 ;
  wire \u2_Display/add137/c11 ;
  wire \u2_Display/add137/c15 ;
  wire \u2_Display/add137/c19 ;
  wire \u2_Display/add137/c23 ;
  wire \u2_Display/add137/c27 ;
  wire \u2_Display/add137/c3 ;
  wire \u2_Display/add137/c31 ;
  wire \u2_Display/add137/c7 ;
  wire \u2_Display/add138/c11 ;
  wire \u2_Display/add138/c15 ;
  wire \u2_Display/add138/c19 ;
  wire \u2_Display/add138/c23 ;
  wire \u2_Display/add138/c27 ;
  wire \u2_Display/add138/c3 ;
  wire \u2_Display/add138/c31 ;
  wire \u2_Display/add138/c7 ;
  wire \u2_Display/add139/c3 ;
  wire \u2_Display/add139/c7 ;
  wire \u2_Display/add14/c11 ;
  wire \u2_Display/add14/c15 ;
  wire \u2_Display/add14/c19 ;
  wire \u2_Display/add14/c23 ;
  wire \u2_Display/add14/c27 ;
  wire \u2_Display/add14/c3 ;
  wire \u2_Display/add14/c31 ;
  wire \u2_Display/add14/c7 ;
  wire \u2_Display/add151/c11 ;
  wire \u2_Display/add151/c15 ;
  wire \u2_Display/add151/c19 ;
  wire \u2_Display/add151/c23 ;
  wire \u2_Display/add151/c27 ;
  wire \u2_Display/add151/c3 ;
  wire \u2_Display/add151/c31 ;
  wire \u2_Display/add151/c7 ;
  wire \u2_Display/add152/c11 ;
  wire \u2_Display/add152/c15 ;
  wire \u2_Display/add152/c19 ;
  wire \u2_Display/add152/c23 ;
  wire \u2_Display/add152/c27 ;
  wire \u2_Display/add152/c3 ;
  wire \u2_Display/add152/c31 ;
  wire \u2_Display/add152/c7 ;
  wire \u2_Display/add153/c11 ;
  wire \u2_Display/add153/c15 ;
  wire \u2_Display/add153/c19 ;
  wire \u2_Display/add153/c23 ;
  wire \u2_Display/add153/c27 ;
  wire \u2_Display/add153/c3 ;
  wire \u2_Display/add153/c31 ;
  wire \u2_Display/add153/c7 ;
  wire \u2_Display/add154/c11 ;
  wire \u2_Display/add154/c15 ;
  wire \u2_Display/add154/c19 ;
  wire \u2_Display/add154/c23 ;
  wire \u2_Display/add154/c27 ;
  wire \u2_Display/add154/c3 ;
  wire \u2_Display/add154/c31 ;
  wire \u2_Display/add154/c7 ;
  wire \u2_Display/add155/c11 ;
  wire \u2_Display/add155/c15 ;
  wire \u2_Display/add155/c19 ;
  wire \u2_Display/add155/c23 ;
  wire \u2_Display/add155/c27 ;
  wire \u2_Display/add155/c3 ;
  wire \u2_Display/add155/c31 ;
  wire \u2_Display/add155/c7 ;
  wire \u2_Display/add156/c11 ;
  wire \u2_Display/add156/c15 ;
  wire \u2_Display/add156/c19 ;
  wire \u2_Display/add156/c23 ;
  wire \u2_Display/add156/c27 ;
  wire \u2_Display/add156/c3 ;
  wire \u2_Display/add156/c31 ;
  wire \u2_Display/add156/c7 ;
  wire \u2_Display/add157/c11 ;
  wire \u2_Display/add157/c15 ;
  wire \u2_Display/add157/c19 ;
  wire \u2_Display/add157/c23 ;
  wire \u2_Display/add157/c27 ;
  wire \u2_Display/add157/c3 ;
  wire \u2_Display/add157/c31 ;
  wire \u2_Display/add157/c7 ;
  wire \u2_Display/add158/c11 ;
  wire \u2_Display/add158/c15 ;
  wire \u2_Display/add158/c19 ;
  wire \u2_Display/add158/c23 ;
  wire \u2_Display/add158/c27 ;
  wire \u2_Display/add158/c3 ;
  wire \u2_Display/add158/c31 ;
  wire \u2_Display/add158/c7 ;
  wire \u2_Display/add159/c11 ;
  wire \u2_Display/add159/c15 ;
  wire \u2_Display/add159/c19 ;
  wire \u2_Display/add159/c23 ;
  wire \u2_Display/add159/c27 ;
  wire \u2_Display/add159/c3 ;
  wire \u2_Display/add159/c31 ;
  wire \u2_Display/add159/c7 ;
  wire \u2_Display/add160/c11 ;
  wire \u2_Display/add160/c15 ;
  wire \u2_Display/add160/c19 ;
  wire \u2_Display/add160/c23 ;
  wire \u2_Display/add160/c27 ;
  wire \u2_Display/add160/c3 ;
  wire \u2_Display/add160/c31 ;
  wire \u2_Display/add160/c7 ;
  wire \u2_Display/add161/c11 ;
  wire \u2_Display/add161/c15 ;
  wire \u2_Display/add161/c19 ;
  wire \u2_Display/add161/c23 ;
  wire \u2_Display/add161/c27 ;
  wire \u2_Display/add161/c3 ;
  wire \u2_Display/add161/c31 ;
  wire \u2_Display/add161/c7 ;
  wire \u2_Display/add162/c11 ;
  wire \u2_Display/add162/c15 ;
  wire \u2_Display/add162/c19 ;
  wire \u2_Display/add162/c23 ;
  wire \u2_Display/add162/c27 ;
  wire \u2_Display/add162/c3 ;
  wire \u2_Display/add162/c31 ;
  wire \u2_Display/add162/c7 ;
  wire \u2_Display/add163/c11 ;
  wire \u2_Display/add163/c15 ;
  wire \u2_Display/add163/c19 ;
  wire \u2_Display/add163/c23 ;
  wire \u2_Display/add163/c27 ;
  wire \u2_Display/add163/c3 ;
  wire \u2_Display/add163/c31 ;
  wire \u2_Display/add163/c7 ;
  wire \u2_Display/add164/c11 ;
  wire \u2_Display/add164/c15 ;
  wire \u2_Display/add164/c19 ;
  wire \u2_Display/add164/c23 ;
  wire \u2_Display/add164/c27 ;
  wire \u2_Display/add164/c3 ;
  wire \u2_Display/add164/c31 ;
  wire \u2_Display/add164/c7 ;
  wire \u2_Display/add165/c11 ;
  wire \u2_Display/add165/c15 ;
  wire \u2_Display/add165/c19 ;
  wire \u2_Display/add165/c23 ;
  wire \u2_Display/add165/c27 ;
  wire \u2_Display/add165/c3 ;
  wire \u2_Display/add165/c31 ;
  wire \u2_Display/add165/c7 ;
  wire \u2_Display/add166/c11 ;
  wire \u2_Display/add166/c15 ;
  wire \u2_Display/add166/c19 ;
  wire \u2_Display/add166/c23 ;
  wire \u2_Display/add166/c27 ;
  wire \u2_Display/add166/c3 ;
  wire \u2_Display/add166/c31 ;
  wire \u2_Display/add166/c7 ;
  wire \u2_Display/add167/c11 ;
  wire \u2_Display/add167/c15 ;
  wire \u2_Display/add167/c19 ;
  wire \u2_Display/add167/c23 ;
  wire \u2_Display/add167/c27 ;
  wire \u2_Display/add167/c3 ;
  wire \u2_Display/add167/c31 ;
  wire \u2_Display/add167/c7 ;
  wire \u2_Display/add168/c11 ;
  wire \u2_Display/add168/c15 ;
  wire \u2_Display/add168/c19 ;
  wire \u2_Display/add168/c23 ;
  wire \u2_Display/add168/c27 ;
  wire \u2_Display/add168/c3 ;
  wire \u2_Display/add168/c31 ;
  wire \u2_Display/add168/c7 ;
  wire \u2_Display/add169/c11 ;
  wire \u2_Display/add169/c15 ;
  wire \u2_Display/add169/c19 ;
  wire \u2_Display/add169/c23 ;
  wire \u2_Display/add169/c27 ;
  wire \u2_Display/add169/c3 ;
  wire \u2_Display/add169/c31 ;
  wire \u2_Display/add169/c7 ;
  wire \u2_Display/add170/c11 ;
  wire \u2_Display/add170/c15 ;
  wire \u2_Display/add170/c19 ;
  wire \u2_Display/add170/c23 ;
  wire \u2_Display/add170/c27 ;
  wire \u2_Display/add170/c3 ;
  wire \u2_Display/add170/c31 ;
  wire \u2_Display/add170/c7 ;
  wire \u2_Display/add171/c11 ;
  wire \u2_Display/add171/c15 ;
  wire \u2_Display/add171/c19 ;
  wire \u2_Display/add171/c23 ;
  wire \u2_Display/add171/c27 ;
  wire \u2_Display/add171/c3 ;
  wire \u2_Display/add171/c31 ;
  wire \u2_Display/add171/c7 ;
  wire \u2_Display/add172/c3 ;
  wire \u2_Display/add172/c7 ;
  wire \u2_Display/add18/c11 ;
  wire \u2_Display/add18/c15 ;
  wire \u2_Display/add18/c19 ;
  wire \u2_Display/add18/c23 ;
  wire \u2_Display/add18/c27 ;
  wire \u2_Display/add18/c3 ;
  wire \u2_Display/add18/c31 ;
  wire \u2_Display/add18/c7 ;
  wire \u2_Display/add19/c11 ;
  wire \u2_Display/add19/c15 ;
  wire \u2_Display/add19/c19 ;
  wire \u2_Display/add19/c23 ;
  wire \u2_Display/add19/c27 ;
  wire \u2_Display/add19/c3 ;
  wire \u2_Display/add19/c31 ;
  wire \u2_Display/add19/c7 ;
  wire \u2_Display/add20/c11 ;
  wire \u2_Display/add20/c15 ;
  wire \u2_Display/add20/c19 ;
  wire \u2_Display/add20/c23 ;
  wire \u2_Display/add20/c27 ;
  wire \u2_Display/add20/c3 ;
  wire \u2_Display/add20/c31 ;
  wire \u2_Display/add20/c7 ;
  wire \u2_Display/add21/c11 ;
  wire \u2_Display/add21/c15 ;
  wire \u2_Display/add21/c19 ;
  wire \u2_Display/add21/c23 ;
  wire \u2_Display/add21/c27 ;
  wire \u2_Display/add21/c3 ;
  wire \u2_Display/add21/c31 ;
  wire \u2_Display/add21/c7 ;
  wire \u2_Display/add22/c11 ;
  wire \u2_Display/add22/c15 ;
  wire \u2_Display/add22/c19 ;
  wire \u2_Display/add22/c23 ;
  wire \u2_Display/add22/c27 ;
  wire \u2_Display/add22/c3 ;
  wire \u2_Display/add22/c31 ;
  wire \u2_Display/add22/c7 ;
  wire \u2_Display/add23/c11 ;
  wire \u2_Display/add23/c15 ;
  wire \u2_Display/add23/c19 ;
  wire \u2_Display/add23/c23 ;
  wire \u2_Display/add23/c27 ;
  wire \u2_Display/add23/c3 ;
  wire \u2_Display/add23/c31 ;
  wire \u2_Display/add23/c7 ;
  wire \u2_Display/add24/c11 ;
  wire \u2_Display/add24/c15 ;
  wire \u2_Display/add24/c19 ;
  wire \u2_Display/add24/c23 ;
  wire \u2_Display/add24/c27 ;
  wire \u2_Display/add24/c3 ;
  wire \u2_Display/add24/c31 ;
  wire \u2_Display/add24/c7 ;
  wire \u2_Display/add25/c11 ;
  wire \u2_Display/add25/c15 ;
  wire \u2_Display/add25/c19 ;
  wire \u2_Display/add25/c23 ;
  wire \u2_Display/add25/c27 ;
  wire \u2_Display/add25/c3 ;
  wire \u2_Display/add25/c31 ;
  wire \u2_Display/add25/c7 ;
  wire \u2_Display/add26/c11 ;
  wire \u2_Display/add26/c15 ;
  wire \u2_Display/add26/c19 ;
  wire \u2_Display/add26/c23 ;
  wire \u2_Display/add26/c27 ;
  wire \u2_Display/add26/c3 ;
  wire \u2_Display/add26/c31 ;
  wire \u2_Display/add26/c7 ;
  wire \u2_Display/add27/c11 ;
  wire \u2_Display/add27/c15 ;
  wire \u2_Display/add27/c19 ;
  wire \u2_Display/add27/c23 ;
  wire \u2_Display/add27/c27 ;
  wire \u2_Display/add27/c3 ;
  wire \u2_Display/add27/c31 ;
  wire \u2_Display/add27/c7 ;
  wire \u2_Display/add28/c11 ;
  wire \u2_Display/add28/c15 ;
  wire \u2_Display/add28/c19 ;
  wire \u2_Display/add28/c23 ;
  wire \u2_Display/add28/c27 ;
  wire \u2_Display/add28/c3 ;
  wire \u2_Display/add28/c31 ;
  wire \u2_Display/add28/c7 ;
  wire \u2_Display/add29/c11 ;
  wire \u2_Display/add29/c15 ;
  wire \u2_Display/add29/c19 ;
  wire \u2_Display/add29/c23 ;
  wire \u2_Display/add29/c27 ;
  wire \u2_Display/add29/c3 ;
  wire \u2_Display/add29/c31 ;
  wire \u2_Display/add29/c7 ;
  wire \u2_Display/add2_2/c1 ;
  wire \u2_Display/add2_2/c3 ;
  wire \u2_Display/add2_2_co ;
  wire \u2_Display/add30/c11 ;
  wire \u2_Display/add30/c15 ;
  wire \u2_Display/add30/c19 ;
  wire \u2_Display/add30/c23 ;
  wire \u2_Display/add30/c27 ;
  wire \u2_Display/add30/c3 ;
  wire \u2_Display/add30/c31 ;
  wire \u2_Display/add30/c7 ;
  wire \u2_Display/add31/c11 ;
  wire \u2_Display/add31/c15 ;
  wire \u2_Display/add31/c19 ;
  wire \u2_Display/add31/c23 ;
  wire \u2_Display/add31/c27 ;
  wire \u2_Display/add31/c3 ;
  wire \u2_Display/add31/c31 ;
  wire \u2_Display/add31/c7 ;
  wire \u2_Display/add32/c11 ;
  wire \u2_Display/add32/c15 ;
  wire \u2_Display/add32/c19 ;
  wire \u2_Display/add32/c23 ;
  wire \u2_Display/add32/c27 ;
  wire \u2_Display/add32/c3 ;
  wire \u2_Display/add32/c31 ;
  wire \u2_Display/add32/c7 ;
  wire \u2_Display/add33/c11 ;
  wire \u2_Display/add33/c15 ;
  wire \u2_Display/add33/c19 ;
  wire \u2_Display/add33/c23 ;
  wire \u2_Display/add33/c27 ;
  wire \u2_Display/add33/c3 ;
  wire \u2_Display/add33/c31 ;
  wire \u2_Display/add33/c7 ;
  wire \u2_Display/add34/c11 ;
  wire \u2_Display/add34/c15 ;
  wire \u2_Display/add34/c19 ;
  wire \u2_Display/add34/c23 ;
  wire \u2_Display/add34/c27 ;
  wire \u2_Display/add34/c3 ;
  wire \u2_Display/add34/c31 ;
  wire \u2_Display/add34/c7 ;
  wire \u2_Display/add35/c11 ;
  wire \u2_Display/add35/c15 ;
  wire \u2_Display/add35/c19 ;
  wire \u2_Display/add35/c23 ;
  wire \u2_Display/add35/c27 ;
  wire \u2_Display/add35/c3 ;
  wire \u2_Display/add35/c31 ;
  wire \u2_Display/add35/c7 ;
  wire \u2_Display/add36/c11 ;
  wire \u2_Display/add36/c15 ;
  wire \u2_Display/add36/c19 ;
  wire \u2_Display/add36/c23 ;
  wire \u2_Display/add36/c27 ;
  wire \u2_Display/add36/c3 ;
  wire \u2_Display/add36/c31 ;
  wire \u2_Display/add36/c7 ;
  wire \u2_Display/add37/c11 ;
  wire \u2_Display/add37/c15 ;
  wire \u2_Display/add37/c19 ;
  wire \u2_Display/add37/c23 ;
  wire \u2_Display/add37/c27 ;
  wire \u2_Display/add37/c3 ;
  wire \u2_Display/add37/c31 ;
  wire \u2_Display/add37/c7 ;
  wire \u2_Display/add38/c11 ;
  wire \u2_Display/add38/c15 ;
  wire \u2_Display/add38/c19 ;
  wire \u2_Display/add38/c23 ;
  wire \u2_Display/add38/c27 ;
  wire \u2_Display/add38/c3 ;
  wire \u2_Display/add38/c31 ;
  wire \u2_Display/add38/c7 ;
  wire \u2_Display/add39/c11 ;
  wire \u2_Display/add39/c15 ;
  wire \u2_Display/add39/c19 ;
  wire \u2_Display/add39/c23 ;
  wire \u2_Display/add39/c27 ;
  wire \u2_Display/add39/c3 ;
  wire \u2_Display/add39/c31 ;
  wire \u2_Display/add39/c7 ;
  wire \u2_Display/add40/c3 ;
  wire \u2_Display/add40/c7 ;
  wire \u2_Display/add4_2/c1 ;
  wire \u2_Display/add4_2/c3 ;
  wire \u2_Display/add4_2_co ;
  wire \u2_Display/add51/c11 ;
  wire \u2_Display/add51/c15 ;
  wire \u2_Display/add51/c19 ;
  wire \u2_Display/add51/c23 ;
  wire \u2_Display/add51/c27 ;
  wire \u2_Display/add51/c3 ;
  wire \u2_Display/add51/c31 ;
  wire \u2_Display/add51/c7 ;
  wire \u2_Display/add52/c11 ;
  wire \u2_Display/add52/c15 ;
  wire \u2_Display/add52/c19 ;
  wire \u2_Display/add52/c23 ;
  wire \u2_Display/add52/c27 ;
  wire \u2_Display/add52/c3 ;
  wire \u2_Display/add52/c31 ;
  wire \u2_Display/add52/c7 ;
  wire \u2_Display/add53/c11 ;
  wire \u2_Display/add53/c15 ;
  wire \u2_Display/add53/c19 ;
  wire \u2_Display/add53/c23 ;
  wire \u2_Display/add53/c27 ;
  wire \u2_Display/add53/c3 ;
  wire \u2_Display/add53/c31 ;
  wire \u2_Display/add53/c7 ;
  wire \u2_Display/add54/c11 ;
  wire \u2_Display/add54/c15 ;
  wire \u2_Display/add54/c19 ;
  wire \u2_Display/add54/c23 ;
  wire \u2_Display/add54/c27 ;
  wire \u2_Display/add54/c3 ;
  wire \u2_Display/add54/c31 ;
  wire \u2_Display/add54/c7 ;
  wire \u2_Display/add55/c11 ;
  wire \u2_Display/add55/c15 ;
  wire \u2_Display/add55/c19 ;
  wire \u2_Display/add55/c23 ;
  wire \u2_Display/add55/c27 ;
  wire \u2_Display/add55/c3 ;
  wire \u2_Display/add55/c31 ;
  wire \u2_Display/add55/c7 ;
  wire \u2_Display/add56/c11 ;
  wire \u2_Display/add56/c15 ;
  wire \u2_Display/add56/c19 ;
  wire \u2_Display/add56/c23 ;
  wire \u2_Display/add56/c27 ;
  wire \u2_Display/add56/c3 ;
  wire \u2_Display/add56/c31 ;
  wire \u2_Display/add56/c7 ;
  wire \u2_Display/add57/c11 ;
  wire \u2_Display/add57/c15 ;
  wire \u2_Display/add57/c19 ;
  wire \u2_Display/add57/c23 ;
  wire \u2_Display/add57/c27 ;
  wire \u2_Display/add57/c3 ;
  wire \u2_Display/add57/c31 ;
  wire \u2_Display/add57/c7 ;
  wire \u2_Display/add58/c11 ;
  wire \u2_Display/add58/c15 ;
  wire \u2_Display/add58/c19 ;
  wire \u2_Display/add58/c23 ;
  wire \u2_Display/add58/c27 ;
  wire \u2_Display/add58/c3 ;
  wire \u2_Display/add58/c31 ;
  wire \u2_Display/add58/c7 ;
  wire \u2_Display/add59/c11 ;
  wire \u2_Display/add59/c15 ;
  wire \u2_Display/add59/c19 ;
  wire \u2_Display/add59/c23 ;
  wire \u2_Display/add59/c27 ;
  wire \u2_Display/add59/c3 ;
  wire \u2_Display/add59/c31 ;
  wire \u2_Display/add59/c7 ;
  wire \u2_Display/add60/c11 ;
  wire \u2_Display/add60/c15 ;
  wire \u2_Display/add60/c19 ;
  wire \u2_Display/add60/c23 ;
  wire \u2_Display/add60/c27 ;
  wire \u2_Display/add60/c3 ;
  wire \u2_Display/add60/c31 ;
  wire \u2_Display/add60/c7 ;
  wire \u2_Display/add61/c11 ;
  wire \u2_Display/add61/c15 ;
  wire \u2_Display/add61/c19 ;
  wire \u2_Display/add61/c23 ;
  wire \u2_Display/add61/c27 ;
  wire \u2_Display/add61/c3 ;
  wire \u2_Display/add61/c31 ;
  wire \u2_Display/add61/c7 ;
  wire \u2_Display/add62/c11 ;
  wire \u2_Display/add62/c15 ;
  wire \u2_Display/add62/c19 ;
  wire \u2_Display/add62/c23 ;
  wire \u2_Display/add62/c27 ;
  wire \u2_Display/add62/c3 ;
  wire \u2_Display/add62/c31 ;
  wire \u2_Display/add62/c7 ;
  wire \u2_Display/add63/c11 ;
  wire \u2_Display/add63/c15 ;
  wire \u2_Display/add63/c19 ;
  wire \u2_Display/add63/c23 ;
  wire \u2_Display/add63/c27 ;
  wire \u2_Display/add63/c3 ;
  wire \u2_Display/add63/c31 ;
  wire \u2_Display/add63/c7 ;
  wire \u2_Display/add64/c11 ;
  wire \u2_Display/add64/c15 ;
  wire \u2_Display/add64/c19 ;
  wire \u2_Display/add64/c23 ;
  wire \u2_Display/add64/c27 ;
  wire \u2_Display/add64/c3 ;
  wire \u2_Display/add64/c31 ;
  wire \u2_Display/add64/c7 ;
  wire \u2_Display/add65/c11 ;
  wire \u2_Display/add65/c15 ;
  wire \u2_Display/add65/c19 ;
  wire \u2_Display/add65/c23 ;
  wire \u2_Display/add65/c27 ;
  wire \u2_Display/add65/c3 ;
  wire \u2_Display/add65/c31 ;
  wire \u2_Display/add65/c7 ;
  wire \u2_Display/add66/c11 ;
  wire \u2_Display/add66/c15 ;
  wire \u2_Display/add66/c19 ;
  wire \u2_Display/add66/c23 ;
  wire \u2_Display/add66/c27 ;
  wire \u2_Display/add66/c3 ;
  wire \u2_Display/add66/c31 ;
  wire \u2_Display/add66/c7 ;
  wire \u2_Display/add67/c11 ;
  wire \u2_Display/add67/c15 ;
  wire \u2_Display/add67/c19 ;
  wire \u2_Display/add67/c23 ;
  wire \u2_Display/add67/c27 ;
  wire \u2_Display/add67/c3 ;
  wire \u2_Display/add67/c31 ;
  wire \u2_Display/add67/c7 ;
  wire \u2_Display/add68/c11 ;
  wire \u2_Display/add68/c15 ;
  wire \u2_Display/add68/c19 ;
  wire \u2_Display/add68/c23 ;
  wire \u2_Display/add68/c27 ;
  wire \u2_Display/add68/c3 ;
  wire \u2_Display/add68/c31 ;
  wire \u2_Display/add68/c7 ;
  wire \u2_Display/add69/c11 ;
  wire \u2_Display/add69/c15 ;
  wire \u2_Display/add69/c19 ;
  wire \u2_Display/add69/c23 ;
  wire \u2_Display/add69/c27 ;
  wire \u2_Display/add69/c3 ;
  wire \u2_Display/add69/c31 ;
  wire \u2_Display/add69/c7 ;
  wire \u2_Display/add6_2/c1 ;
  wire \u2_Display/add6_2/c3 ;
  wire \u2_Display/add6_2_co ;
  wire \u2_Display/add70/c11 ;
  wire \u2_Display/add70/c15 ;
  wire \u2_Display/add70/c19 ;
  wire \u2_Display/add70/c23 ;
  wire \u2_Display/add70/c27 ;
  wire \u2_Display/add70/c3 ;
  wire \u2_Display/add70/c31 ;
  wire \u2_Display/add70/c7 ;
  wire \u2_Display/add71/c11 ;
  wire \u2_Display/add71/c15 ;
  wire \u2_Display/add71/c19 ;
  wire \u2_Display/add71/c23 ;
  wire \u2_Display/add71/c27 ;
  wire \u2_Display/add71/c3 ;
  wire \u2_Display/add71/c31 ;
  wire \u2_Display/add71/c7 ;
  wire \u2_Display/add72/c11 ;
  wire \u2_Display/add72/c15 ;
  wire \u2_Display/add72/c19 ;
  wire \u2_Display/add72/c23 ;
  wire \u2_Display/add72/c27 ;
  wire \u2_Display/add72/c3 ;
  wire \u2_Display/add72/c31 ;
  wire \u2_Display/add72/c7 ;
  wire \u2_Display/add73/c3 ;
  wire \u2_Display/add73/c7 ;
  wire \u2_Display/add7_2_co ;
  wire \u2_Display/add84/c11 ;
  wire \u2_Display/add84/c15 ;
  wire \u2_Display/add84/c19 ;
  wire \u2_Display/add84/c23 ;
  wire \u2_Display/add84/c27 ;
  wire \u2_Display/add84/c3 ;
  wire \u2_Display/add84/c31 ;
  wire \u2_Display/add84/c7 ;
  wire \u2_Display/add85/c11 ;
  wire \u2_Display/add85/c15 ;
  wire \u2_Display/add85/c19 ;
  wire \u2_Display/add85/c23 ;
  wire \u2_Display/add85/c27 ;
  wire \u2_Display/add85/c3 ;
  wire \u2_Display/add85/c31 ;
  wire \u2_Display/add85/c7 ;
  wire \u2_Display/add86/c11 ;
  wire \u2_Display/add86/c15 ;
  wire \u2_Display/add86/c19 ;
  wire \u2_Display/add86/c23 ;
  wire \u2_Display/add86/c27 ;
  wire \u2_Display/add86/c3 ;
  wire \u2_Display/add86/c31 ;
  wire \u2_Display/add86/c7 ;
  wire \u2_Display/add87/c11 ;
  wire \u2_Display/add87/c15 ;
  wire \u2_Display/add87/c19 ;
  wire \u2_Display/add87/c23 ;
  wire \u2_Display/add87/c27 ;
  wire \u2_Display/add87/c3 ;
  wire \u2_Display/add87/c31 ;
  wire \u2_Display/add87/c7 ;
  wire \u2_Display/add88/c11 ;
  wire \u2_Display/add88/c15 ;
  wire \u2_Display/add88/c19 ;
  wire \u2_Display/add88/c23 ;
  wire \u2_Display/add88/c27 ;
  wire \u2_Display/add88/c3 ;
  wire \u2_Display/add88/c31 ;
  wire \u2_Display/add88/c7 ;
  wire \u2_Display/add89/c11 ;
  wire \u2_Display/add89/c15 ;
  wire \u2_Display/add89/c19 ;
  wire \u2_Display/add89/c23 ;
  wire \u2_Display/add89/c27 ;
  wire \u2_Display/add89/c3 ;
  wire \u2_Display/add89/c31 ;
  wire \u2_Display/add89/c7 ;
  wire \u2_Display/add90/c11 ;
  wire \u2_Display/add90/c15 ;
  wire \u2_Display/add90/c19 ;
  wire \u2_Display/add90/c23 ;
  wire \u2_Display/add90/c27 ;
  wire \u2_Display/add90/c3 ;
  wire \u2_Display/add90/c31 ;
  wire \u2_Display/add90/c7 ;
  wire \u2_Display/add91/c11 ;
  wire \u2_Display/add91/c15 ;
  wire \u2_Display/add91/c19 ;
  wire \u2_Display/add91/c23 ;
  wire \u2_Display/add91/c27 ;
  wire \u2_Display/add91/c3 ;
  wire \u2_Display/add91/c31 ;
  wire \u2_Display/add91/c7 ;
  wire \u2_Display/add92/c11 ;
  wire \u2_Display/add92/c15 ;
  wire \u2_Display/add92/c19 ;
  wire \u2_Display/add92/c23 ;
  wire \u2_Display/add92/c27 ;
  wire \u2_Display/add92/c3 ;
  wire \u2_Display/add92/c31 ;
  wire \u2_Display/add92/c7 ;
  wire \u2_Display/add93/c11 ;
  wire \u2_Display/add93/c15 ;
  wire \u2_Display/add93/c19 ;
  wire \u2_Display/add93/c23 ;
  wire \u2_Display/add93/c27 ;
  wire \u2_Display/add93/c3 ;
  wire \u2_Display/add93/c31 ;
  wire \u2_Display/add93/c7 ;
  wire \u2_Display/add94/c11 ;
  wire \u2_Display/add94/c15 ;
  wire \u2_Display/add94/c19 ;
  wire \u2_Display/add94/c23 ;
  wire \u2_Display/add94/c27 ;
  wire \u2_Display/add94/c3 ;
  wire \u2_Display/add94/c31 ;
  wire \u2_Display/add94/c7 ;
  wire \u2_Display/add95/c11 ;
  wire \u2_Display/add95/c15 ;
  wire \u2_Display/add95/c19 ;
  wire \u2_Display/add95/c23 ;
  wire \u2_Display/add95/c27 ;
  wire \u2_Display/add95/c3 ;
  wire \u2_Display/add95/c31 ;
  wire \u2_Display/add95/c7 ;
  wire \u2_Display/add96/c11 ;
  wire \u2_Display/add96/c15 ;
  wire \u2_Display/add96/c19 ;
  wire \u2_Display/add96/c23 ;
  wire \u2_Display/add96/c27 ;
  wire \u2_Display/add96/c3 ;
  wire \u2_Display/add96/c31 ;
  wire \u2_Display/add96/c7 ;
  wire \u2_Display/add97/c11 ;
  wire \u2_Display/add97/c15 ;
  wire \u2_Display/add97/c19 ;
  wire \u2_Display/add97/c23 ;
  wire \u2_Display/add97/c27 ;
  wire \u2_Display/add97/c3 ;
  wire \u2_Display/add97/c31 ;
  wire \u2_Display/add97/c7 ;
  wire \u2_Display/add98/c11 ;
  wire \u2_Display/add98/c15 ;
  wire \u2_Display/add98/c19 ;
  wire \u2_Display/add98/c23 ;
  wire \u2_Display/add98/c27 ;
  wire \u2_Display/add98/c3 ;
  wire \u2_Display/add98/c31 ;
  wire \u2_Display/add98/c7 ;
  wire \u2_Display/add99/c11 ;
  wire \u2_Display/add99/c15 ;
  wire \u2_Display/add99/c19 ;
  wire \u2_Display/add99/c23 ;
  wire \u2_Display/add99/c27 ;
  wire \u2_Display/add99/c3 ;
  wire \u2_Display/add99/c31 ;
  wire \u2_Display/add99/c7 ;
  wire \u2_Display/clk1s ;  // source/rtl/Display.v(46)
  wire \u2_Display/lt0_2_c1 ;
  wire \u2_Display/lt0_2_c11 ;
  wire \u2_Display/lt0_2_c3 ;
  wire \u2_Display/lt0_2_c5 ;
  wire \u2_Display/lt0_2_c7 ;
  wire \u2_Display/lt0_2_c9 ;
  wire \u2_Display/lt100_c1 ;
  wire \u2_Display/lt100_c11 ;
  wire \u2_Display/lt100_c13 ;
  wire \u2_Display/lt100_c15 ;
  wire \u2_Display/lt100_c17 ;
  wire \u2_Display/lt100_c19 ;
  wire \u2_Display/lt100_c21 ;
  wire \u2_Display/lt100_c23 ;
  wire \u2_Display/lt100_c25 ;
  wire \u2_Display/lt100_c27 ;
  wire \u2_Display/lt100_c29 ;
  wire \u2_Display/lt100_c3 ;
  wire \u2_Display/lt100_c31 ;
  wire \u2_Display/lt100_c5 ;
  wire \u2_Display/lt100_c7 ;
  wire \u2_Display/lt100_c9 ;
  wire \u2_Display/lt101_c1 ;
  wire \u2_Display/lt101_c11 ;
  wire \u2_Display/lt101_c13 ;
  wire \u2_Display/lt101_c15 ;
  wire \u2_Display/lt101_c17 ;
  wire \u2_Display/lt101_c19 ;
  wire \u2_Display/lt101_c21 ;
  wire \u2_Display/lt101_c23 ;
  wire \u2_Display/lt101_c25 ;
  wire \u2_Display/lt101_c27 ;
  wire \u2_Display/lt101_c29 ;
  wire \u2_Display/lt101_c3 ;
  wire \u2_Display/lt101_c31 ;
  wire \u2_Display/lt101_c5 ;
  wire \u2_Display/lt101_c7 ;
  wire \u2_Display/lt101_c9 ;
  wire \u2_Display/lt102_c1 ;
  wire \u2_Display/lt102_c11 ;
  wire \u2_Display/lt102_c13 ;
  wire \u2_Display/lt102_c15 ;
  wire \u2_Display/lt102_c17 ;
  wire \u2_Display/lt102_c19 ;
  wire \u2_Display/lt102_c21 ;
  wire \u2_Display/lt102_c23 ;
  wire \u2_Display/lt102_c25 ;
  wire \u2_Display/lt102_c27 ;
  wire \u2_Display/lt102_c29 ;
  wire \u2_Display/lt102_c3 ;
  wire \u2_Display/lt102_c31 ;
  wire \u2_Display/lt102_c5 ;
  wire \u2_Display/lt102_c7 ;
  wire \u2_Display/lt102_c9 ;
  wire \u2_Display/lt103_c1 ;
  wire \u2_Display/lt103_c11 ;
  wire \u2_Display/lt103_c13 ;
  wire \u2_Display/lt103_c15 ;
  wire \u2_Display/lt103_c17 ;
  wire \u2_Display/lt103_c19 ;
  wire \u2_Display/lt103_c21 ;
  wire \u2_Display/lt103_c23 ;
  wire \u2_Display/lt103_c25 ;
  wire \u2_Display/lt103_c27 ;
  wire \u2_Display/lt103_c29 ;
  wire \u2_Display/lt103_c3 ;
  wire \u2_Display/lt103_c31 ;
  wire \u2_Display/lt103_c5 ;
  wire \u2_Display/lt103_c7 ;
  wire \u2_Display/lt103_c9 ;
  wire \u2_Display/lt104_c1 ;
  wire \u2_Display/lt104_c11 ;
  wire \u2_Display/lt104_c13 ;
  wire \u2_Display/lt104_c15 ;
  wire \u2_Display/lt104_c17 ;
  wire \u2_Display/lt104_c19 ;
  wire \u2_Display/lt104_c21 ;
  wire \u2_Display/lt104_c23 ;
  wire \u2_Display/lt104_c25 ;
  wire \u2_Display/lt104_c27 ;
  wire \u2_Display/lt104_c29 ;
  wire \u2_Display/lt104_c3 ;
  wire \u2_Display/lt104_c31 ;
  wire \u2_Display/lt104_c5 ;
  wire \u2_Display/lt104_c7 ;
  wire \u2_Display/lt104_c9 ;
  wire \u2_Display/lt105_c1 ;
  wire \u2_Display/lt105_c11 ;
  wire \u2_Display/lt105_c13 ;
  wire \u2_Display/lt105_c15 ;
  wire \u2_Display/lt105_c17 ;
  wire \u2_Display/lt105_c19 ;
  wire \u2_Display/lt105_c21 ;
  wire \u2_Display/lt105_c23 ;
  wire \u2_Display/lt105_c25 ;
  wire \u2_Display/lt105_c27 ;
  wire \u2_Display/lt105_c29 ;
  wire \u2_Display/lt105_c3 ;
  wire \u2_Display/lt105_c31 ;
  wire \u2_Display/lt105_c5 ;
  wire \u2_Display/lt105_c7 ;
  wire \u2_Display/lt105_c9 ;
  wire \u2_Display/lt106_c1 ;
  wire \u2_Display/lt106_c11 ;
  wire \u2_Display/lt106_c13 ;
  wire \u2_Display/lt106_c15 ;
  wire \u2_Display/lt106_c17 ;
  wire \u2_Display/lt106_c19 ;
  wire \u2_Display/lt106_c21 ;
  wire \u2_Display/lt106_c23 ;
  wire \u2_Display/lt106_c25 ;
  wire \u2_Display/lt106_c27 ;
  wire \u2_Display/lt106_c29 ;
  wire \u2_Display/lt106_c3 ;
  wire \u2_Display/lt106_c31 ;
  wire \u2_Display/lt106_c5 ;
  wire \u2_Display/lt106_c7 ;
  wire \u2_Display/lt106_c9 ;
  wire \u2_Display/lt107_c1 ;
  wire \u2_Display/lt107_c11 ;
  wire \u2_Display/lt107_c13 ;
  wire \u2_Display/lt107_c15 ;
  wire \u2_Display/lt107_c17 ;
  wire \u2_Display/lt107_c19 ;
  wire \u2_Display/lt107_c21 ;
  wire \u2_Display/lt107_c23 ;
  wire \u2_Display/lt107_c25 ;
  wire \u2_Display/lt107_c27 ;
  wire \u2_Display/lt107_c29 ;
  wire \u2_Display/lt107_c3 ;
  wire \u2_Display/lt107_c31 ;
  wire \u2_Display/lt107_c5 ;
  wire \u2_Display/lt107_c7 ;
  wire \u2_Display/lt107_c9 ;
  wire \u2_Display/lt108_c1 ;
  wire \u2_Display/lt108_c11 ;
  wire \u2_Display/lt108_c13 ;
  wire \u2_Display/lt108_c15 ;
  wire \u2_Display/lt108_c17 ;
  wire \u2_Display/lt108_c19 ;
  wire \u2_Display/lt108_c21 ;
  wire \u2_Display/lt108_c23 ;
  wire \u2_Display/lt108_c25 ;
  wire \u2_Display/lt108_c27 ;
  wire \u2_Display/lt108_c29 ;
  wire \u2_Display/lt108_c3 ;
  wire \u2_Display/lt108_c31 ;
  wire \u2_Display/lt108_c5 ;
  wire \u2_Display/lt108_c7 ;
  wire \u2_Display/lt108_c9 ;
  wire \u2_Display/lt109_c1 ;
  wire \u2_Display/lt109_c11 ;
  wire \u2_Display/lt109_c13 ;
  wire \u2_Display/lt109_c15 ;
  wire \u2_Display/lt109_c17 ;
  wire \u2_Display/lt109_c19 ;
  wire \u2_Display/lt109_c21 ;
  wire \u2_Display/lt109_c23 ;
  wire \u2_Display/lt109_c25 ;
  wire \u2_Display/lt109_c27 ;
  wire \u2_Display/lt109_c29 ;
  wire \u2_Display/lt109_c3 ;
  wire \u2_Display/lt109_c31 ;
  wire \u2_Display/lt109_c5 ;
  wire \u2_Display/lt109_c7 ;
  wire \u2_Display/lt109_c9 ;
  wire \u2_Display/lt10_2_c1 ;
  wire \u2_Display/lt10_2_c11 ;
  wire \u2_Display/lt10_2_c3 ;
  wire \u2_Display/lt10_2_c5 ;
  wire \u2_Display/lt10_2_c7 ;
  wire \u2_Display/lt10_2_c9 ;
  wire \u2_Display/lt110_c1 ;
  wire \u2_Display/lt110_c11 ;
  wire \u2_Display/lt110_c13 ;
  wire \u2_Display/lt110_c15 ;
  wire \u2_Display/lt110_c17 ;
  wire \u2_Display/lt110_c19 ;
  wire \u2_Display/lt110_c21 ;
  wire \u2_Display/lt110_c23 ;
  wire \u2_Display/lt110_c25 ;
  wire \u2_Display/lt110_c27 ;
  wire \u2_Display/lt110_c29 ;
  wire \u2_Display/lt110_c3 ;
  wire \u2_Display/lt110_c31 ;
  wire \u2_Display/lt110_c5 ;
  wire \u2_Display/lt110_c7 ;
  wire \u2_Display/lt110_c9 ;
  wire \u2_Display/lt11_2_c1 ;
  wire \u2_Display/lt11_2_c11 ;
  wire \u2_Display/lt11_2_c13 ;
  wire \u2_Display/lt11_2_c3 ;
  wire \u2_Display/lt11_2_c5 ;
  wire \u2_Display/lt11_2_c7 ;
  wire \u2_Display/lt11_2_c9 ;
  wire \u2_Display/lt121_c1 ;
  wire \u2_Display/lt121_c11 ;
  wire \u2_Display/lt121_c13 ;
  wire \u2_Display/lt121_c15 ;
  wire \u2_Display/lt121_c17 ;
  wire \u2_Display/lt121_c19 ;
  wire \u2_Display/lt121_c21 ;
  wire \u2_Display/lt121_c23 ;
  wire \u2_Display/lt121_c25 ;
  wire \u2_Display/lt121_c27 ;
  wire \u2_Display/lt121_c29 ;
  wire \u2_Display/lt121_c3 ;
  wire \u2_Display/lt121_c31 ;
  wire \u2_Display/lt121_c5 ;
  wire \u2_Display/lt121_c7 ;
  wire \u2_Display/lt121_c9 ;
  wire \u2_Display/lt122_c1 ;
  wire \u2_Display/lt122_c11 ;
  wire \u2_Display/lt122_c13 ;
  wire \u2_Display/lt122_c15 ;
  wire \u2_Display/lt122_c17 ;
  wire \u2_Display/lt122_c19 ;
  wire \u2_Display/lt122_c21 ;
  wire \u2_Display/lt122_c23 ;
  wire \u2_Display/lt122_c25 ;
  wire \u2_Display/lt122_c27 ;
  wire \u2_Display/lt122_c29 ;
  wire \u2_Display/lt122_c3 ;
  wire \u2_Display/lt122_c31 ;
  wire \u2_Display/lt122_c5 ;
  wire \u2_Display/lt122_c7 ;
  wire \u2_Display/lt122_c9 ;
  wire \u2_Display/lt123_c1 ;
  wire \u2_Display/lt123_c11 ;
  wire \u2_Display/lt123_c13 ;
  wire \u2_Display/lt123_c15 ;
  wire \u2_Display/lt123_c17 ;
  wire \u2_Display/lt123_c19 ;
  wire \u2_Display/lt123_c21 ;
  wire \u2_Display/lt123_c23 ;
  wire \u2_Display/lt123_c25 ;
  wire \u2_Display/lt123_c27 ;
  wire \u2_Display/lt123_c29 ;
  wire \u2_Display/lt123_c3 ;
  wire \u2_Display/lt123_c31 ;
  wire \u2_Display/lt123_c5 ;
  wire \u2_Display/lt123_c7 ;
  wire \u2_Display/lt123_c9 ;
  wire \u2_Display/lt124_c1 ;
  wire \u2_Display/lt124_c11 ;
  wire \u2_Display/lt124_c13 ;
  wire \u2_Display/lt124_c15 ;
  wire \u2_Display/lt124_c17 ;
  wire \u2_Display/lt124_c19 ;
  wire \u2_Display/lt124_c21 ;
  wire \u2_Display/lt124_c23 ;
  wire \u2_Display/lt124_c25 ;
  wire \u2_Display/lt124_c27 ;
  wire \u2_Display/lt124_c29 ;
  wire \u2_Display/lt124_c3 ;
  wire \u2_Display/lt124_c31 ;
  wire \u2_Display/lt124_c5 ;
  wire \u2_Display/lt124_c7 ;
  wire \u2_Display/lt124_c9 ;
  wire \u2_Display/lt125_c1 ;
  wire \u2_Display/lt125_c11 ;
  wire \u2_Display/lt125_c13 ;
  wire \u2_Display/lt125_c15 ;
  wire \u2_Display/lt125_c17 ;
  wire \u2_Display/lt125_c19 ;
  wire \u2_Display/lt125_c21 ;
  wire \u2_Display/lt125_c23 ;
  wire \u2_Display/lt125_c25 ;
  wire \u2_Display/lt125_c27 ;
  wire \u2_Display/lt125_c29 ;
  wire \u2_Display/lt125_c3 ;
  wire \u2_Display/lt125_c31 ;
  wire \u2_Display/lt125_c5 ;
  wire \u2_Display/lt125_c7 ;
  wire \u2_Display/lt125_c9 ;
  wire \u2_Display/lt126_c1 ;
  wire \u2_Display/lt126_c11 ;
  wire \u2_Display/lt126_c13 ;
  wire \u2_Display/lt126_c15 ;
  wire \u2_Display/lt126_c17 ;
  wire \u2_Display/lt126_c19 ;
  wire \u2_Display/lt126_c21 ;
  wire \u2_Display/lt126_c23 ;
  wire \u2_Display/lt126_c25 ;
  wire \u2_Display/lt126_c27 ;
  wire \u2_Display/lt126_c29 ;
  wire \u2_Display/lt126_c3 ;
  wire \u2_Display/lt126_c31 ;
  wire \u2_Display/lt126_c5 ;
  wire \u2_Display/lt126_c7 ;
  wire \u2_Display/lt126_c9 ;
  wire \u2_Display/lt127_c1 ;
  wire \u2_Display/lt127_c11 ;
  wire \u2_Display/lt127_c13 ;
  wire \u2_Display/lt127_c15 ;
  wire \u2_Display/lt127_c17 ;
  wire \u2_Display/lt127_c19 ;
  wire \u2_Display/lt127_c21 ;
  wire \u2_Display/lt127_c23 ;
  wire \u2_Display/lt127_c25 ;
  wire \u2_Display/lt127_c27 ;
  wire \u2_Display/lt127_c29 ;
  wire \u2_Display/lt127_c3 ;
  wire \u2_Display/lt127_c31 ;
  wire \u2_Display/lt127_c5 ;
  wire \u2_Display/lt127_c7 ;
  wire \u2_Display/lt127_c9 ;
  wire \u2_Display/lt128_c1 ;
  wire \u2_Display/lt128_c11 ;
  wire \u2_Display/lt128_c13 ;
  wire \u2_Display/lt128_c15 ;
  wire \u2_Display/lt128_c17 ;
  wire \u2_Display/lt128_c19 ;
  wire \u2_Display/lt128_c21 ;
  wire \u2_Display/lt128_c23 ;
  wire \u2_Display/lt128_c25 ;
  wire \u2_Display/lt128_c27 ;
  wire \u2_Display/lt128_c29 ;
  wire \u2_Display/lt128_c3 ;
  wire \u2_Display/lt128_c31 ;
  wire \u2_Display/lt128_c5 ;
  wire \u2_Display/lt128_c7 ;
  wire \u2_Display/lt128_c9 ;
  wire \u2_Display/lt129_c1 ;
  wire \u2_Display/lt129_c11 ;
  wire \u2_Display/lt129_c13 ;
  wire \u2_Display/lt129_c15 ;
  wire \u2_Display/lt129_c17 ;
  wire \u2_Display/lt129_c19 ;
  wire \u2_Display/lt129_c21 ;
  wire \u2_Display/lt129_c23 ;
  wire \u2_Display/lt129_c25 ;
  wire \u2_Display/lt129_c27 ;
  wire \u2_Display/lt129_c29 ;
  wire \u2_Display/lt129_c3 ;
  wire \u2_Display/lt129_c31 ;
  wire \u2_Display/lt129_c5 ;
  wire \u2_Display/lt129_c7 ;
  wire \u2_Display/lt129_c9 ;
  wire \u2_Display/lt130_c1 ;
  wire \u2_Display/lt130_c11 ;
  wire \u2_Display/lt130_c13 ;
  wire \u2_Display/lt130_c15 ;
  wire \u2_Display/lt130_c17 ;
  wire \u2_Display/lt130_c19 ;
  wire \u2_Display/lt130_c21 ;
  wire \u2_Display/lt130_c23 ;
  wire \u2_Display/lt130_c25 ;
  wire \u2_Display/lt130_c27 ;
  wire \u2_Display/lt130_c29 ;
  wire \u2_Display/lt130_c3 ;
  wire \u2_Display/lt130_c31 ;
  wire \u2_Display/lt130_c5 ;
  wire \u2_Display/lt130_c7 ;
  wire \u2_Display/lt130_c9 ;
  wire \u2_Display/lt131_c1 ;
  wire \u2_Display/lt131_c11 ;
  wire \u2_Display/lt131_c13 ;
  wire \u2_Display/lt131_c15 ;
  wire \u2_Display/lt131_c17 ;
  wire \u2_Display/lt131_c19 ;
  wire \u2_Display/lt131_c21 ;
  wire \u2_Display/lt131_c23 ;
  wire \u2_Display/lt131_c25 ;
  wire \u2_Display/lt131_c27 ;
  wire \u2_Display/lt131_c29 ;
  wire \u2_Display/lt131_c3 ;
  wire \u2_Display/lt131_c31 ;
  wire \u2_Display/lt131_c5 ;
  wire \u2_Display/lt131_c7 ;
  wire \u2_Display/lt131_c9 ;
  wire \u2_Display/lt132_c1 ;
  wire \u2_Display/lt132_c11 ;
  wire \u2_Display/lt132_c13 ;
  wire \u2_Display/lt132_c15 ;
  wire \u2_Display/lt132_c17 ;
  wire \u2_Display/lt132_c19 ;
  wire \u2_Display/lt132_c21 ;
  wire \u2_Display/lt132_c23 ;
  wire \u2_Display/lt132_c25 ;
  wire \u2_Display/lt132_c27 ;
  wire \u2_Display/lt132_c29 ;
  wire \u2_Display/lt132_c3 ;
  wire \u2_Display/lt132_c31 ;
  wire \u2_Display/lt132_c5 ;
  wire \u2_Display/lt132_c7 ;
  wire \u2_Display/lt132_c9 ;
  wire \u2_Display/lt133_c1 ;
  wire \u2_Display/lt133_c11 ;
  wire \u2_Display/lt133_c13 ;
  wire \u2_Display/lt133_c15 ;
  wire \u2_Display/lt133_c17 ;
  wire \u2_Display/lt133_c19 ;
  wire \u2_Display/lt133_c21 ;
  wire \u2_Display/lt133_c23 ;
  wire \u2_Display/lt133_c25 ;
  wire \u2_Display/lt133_c27 ;
  wire \u2_Display/lt133_c29 ;
  wire \u2_Display/lt133_c3 ;
  wire \u2_Display/lt133_c31 ;
  wire \u2_Display/lt133_c5 ;
  wire \u2_Display/lt133_c7 ;
  wire \u2_Display/lt133_c9 ;
  wire \u2_Display/lt134_c1 ;
  wire \u2_Display/lt134_c11 ;
  wire \u2_Display/lt134_c13 ;
  wire \u2_Display/lt134_c15 ;
  wire \u2_Display/lt134_c17 ;
  wire \u2_Display/lt134_c19 ;
  wire \u2_Display/lt134_c21 ;
  wire \u2_Display/lt134_c23 ;
  wire \u2_Display/lt134_c25 ;
  wire \u2_Display/lt134_c27 ;
  wire \u2_Display/lt134_c29 ;
  wire \u2_Display/lt134_c3 ;
  wire \u2_Display/lt134_c31 ;
  wire \u2_Display/lt134_c5 ;
  wire \u2_Display/lt134_c7 ;
  wire \u2_Display/lt134_c9 ;
  wire \u2_Display/lt135_c1 ;
  wire \u2_Display/lt135_c11 ;
  wire \u2_Display/lt135_c13 ;
  wire \u2_Display/lt135_c15 ;
  wire \u2_Display/lt135_c17 ;
  wire \u2_Display/lt135_c19 ;
  wire \u2_Display/lt135_c21 ;
  wire \u2_Display/lt135_c23 ;
  wire \u2_Display/lt135_c25 ;
  wire \u2_Display/lt135_c27 ;
  wire \u2_Display/lt135_c29 ;
  wire \u2_Display/lt135_c3 ;
  wire \u2_Display/lt135_c31 ;
  wire \u2_Display/lt135_c5 ;
  wire \u2_Display/lt135_c7 ;
  wire \u2_Display/lt135_c9 ;
  wire \u2_Display/lt136_c1 ;
  wire \u2_Display/lt136_c11 ;
  wire \u2_Display/lt136_c13 ;
  wire \u2_Display/lt136_c15 ;
  wire \u2_Display/lt136_c17 ;
  wire \u2_Display/lt136_c19 ;
  wire \u2_Display/lt136_c21 ;
  wire \u2_Display/lt136_c23 ;
  wire \u2_Display/lt136_c25 ;
  wire \u2_Display/lt136_c27 ;
  wire \u2_Display/lt136_c29 ;
  wire \u2_Display/lt136_c3 ;
  wire \u2_Display/lt136_c31 ;
  wire \u2_Display/lt136_c5 ;
  wire \u2_Display/lt136_c7 ;
  wire \u2_Display/lt136_c9 ;
  wire \u2_Display/lt137_c1 ;
  wire \u2_Display/lt137_c11 ;
  wire \u2_Display/lt137_c13 ;
  wire \u2_Display/lt137_c15 ;
  wire \u2_Display/lt137_c17 ;
  wire \u2_Display/lt137_c19 ;
  wire \u2_Display/lt137_c21 ;
  wire \u2_Display/lt137_c23 ;
  wire \u2_Display/lt137_c25 ;
  wire \u2_Display/lt137_c27 ;
  wire \u2_Display/lt137_c29 ;
  wire \u2_Display/lt137_c3 ;
  wire \u2_Display/lt137_c31 ;
  wire \u2_Display/lt137_c5 ;
  wire \u2_Display/lt137_c7 ;
  wire \u2_Display/lt137_c9 ;
  wire \u2_Display/lt138_c1 ;
  wire \u2_Display/lt138_c11 ;
  wire \u2_Display/lt138_c13 ;
  wire \u2_Display/lt138_c15 ;
  wire \u2_Display/lt138_c17 ;
  wire \u2_Display/lt138_c19 ;
  wire \u2_Display/lt138_c21 ;
  wire \u2_Display/lt138_c23 ;
  wire \u2_Display/lt138_c25 ;
  wire \u2_Display/lt138_c27 ;
  wire \u2_Display/lt138_c29 ;
  wire \u2_Display/lt138_c3 ;
  wire \u2_Display/lt138_c31 ;
  wire \u2_Display/lt138_c5 ;
  wire \u2_Display/lt138_c7 ;
  wire \u2_Display/lt138_c9 ;
  wire \u2_Display/lt139_c1 ;
  wire \u2_Display/lt139_c11 ;
  wire \u2_Display/lt139_c13 ;
  wire \u2_Display/lt139_c15 ;
  wire \u2_Display/lt139_c17 ;
  wire \u2_Display/lt139_c19 ;
  wire \u2_Display/lt139_c21 ;
  wire \u2_Display/lt139_c23 ;
  wire \u2_Display/lt139_c25 ;
  wire \u2_Display/lt139_c27 ;
  wire \u2_Display/lt139_c29 ;
  wire \u2_Display/lt139_c3 ;
  wire \u2_Display/lt139_c31 ;
  wire \u2_Display/lt139_c5 ;
  wire \u2_Display/lt139_c7 ;
  wire \u2_Display/lt139_c9 ;
  wire \u2_Display/lt140_c1 ;
  wire \u2_Display/lt140_c11 ;
  wire \u2_Display/lt140_c13 ;
  wire \u2_Display/lt140_c15 ;
  wire \u2_Display/lt140_c17 ;
  wire \u2_Display/lt140_c19 ;
  wire \u2_Display/lt140_c21 ;
  wire \u2_Display/lt140_c23 ;
  wire \u2_Display/lt140_c25 ;
  wire \u2_Display/lt140_c27 ;
  wire \u2_Display/lt140_c29 ;
  wire \u2_Display/lt140_c3 ;
  wire \u2_Display/lt140_c31 ;
  wire \u2_Display/lt140_c5 ;
  wire \u2_Display/lt140_c7 ;
  wire \u2_Display/lt140_c9 ;
  wire \u2_Display/lt141_c1 ;
  wire \u2_Display/lt141_c11 ;
  wire \u2_Display/lt141_c13 ;
  wire \u2_Display/lt141_c15 ;
  wire \u2_Display/lt141_c17 ;
  wire \u2_Display/lt141_c19 ;
  wire \u2_Display/lt141_c21 ;
  wire \u2_Display/lt141_c23 ;
  wire \u2_Display/lt141_c25 ;
  wire \u2_Display/lt141_c27 ;
  wire \u2_Display/lt141_c29 ;
  wire \u2_Display/lt141_c3 ;
  wire \u2_Display/lt141_c31 ;
  wire \u2_Display/lt141_c5 ;
  wire \u2_Display/lt141_c7 ;
  wire \u2_Display/lt141_c9 ;
  wire \u2_Display/lt142_c1 ;
  wire \u2_Display/lt142_c11 ;
  wire \u2_Display/lt142_c13 ;
  wire \u2_Display/lt142_c15 ;
  wire \u2_Display/lt142_c17 ;
  wire \u2_Display/lt142_c19 ;
  wire \u2_Display/lt142_c21 ;
  wire \u2_Display/lt142_c23 ;
  wire \u2_Display/lt142_c25 ;
  wire \u2_Display/lt142_c27 ;
  wire \u2_Display/lt142_c29 ;
  wire \u2_Display/lt142_c3 ;
  wire \u2_Display/lt142_c31 ;
  wire \u2_Display/lt142_c5 ;
  wire \u2_Display/lt142_c7 ;
  wire \u2_Display/lt142_c9 ;
  wire \u2_Display/lt143_c1 ;
  wire \u2_Display/lt143_c11 ;
  wire \u2_Display/lt143_c13 ;
  wire \u2_Display/lt143_c15 ;
  wire \u2_Display/lt143_c17 ;
  wire \u2_Display/lt143_c19 ;
  wire \u2_Display/lt143_c21 ;
  wire \u2_Display/lt143_c23 ;
  wire \u2_Display/lt143_c25 ;
  wire \u2_Display/lt143_c27 ;
  wire \u2_Display/lt143_c29 ;
  wire \u2_Display/lt143_c3 ;
  wire \u2_Display/lt143_c31 ;
  wire \u2_Display/lt143_c5 ;
  wire \u2_Display/lt143_c7 ;
  wire \u2_Display/lt143_c9 ;
  wire \u2_Display/lt154_c1 ;
  wire \u2_Display/lt154_c11 ;
  wire \u2_Display/lt154_c13 ;
  wire \u2_Display/lt154_c15 ;
  wire \u2_Display/lt154_c17 ;
  wire \u2_Display/lt154_c19 ;
  wire \u2_Display/lt154_c21 ;
  wire \u2_Display/lt154_c23 ;
  wire \u2_Display/lt154_c25 ;
  wire \u2_Display/lt154_c27 ;
  wire \u2_Display/lt154_c29 ;
  wire \u2_Display/lt154_c3 ;
  wire \u2_Display/lt154_c31 ;
  wire \u2_Display/lt154_c5 ;
  wire \u2_Display/lt154_c7 ;
  wire \u2_Display/lt154_c9 ;
  wire \u2_Display/lt155_c1 ;
  wire \u2_Display/lt155_c11 ;
  wire \u2_Display/lt155_c13 ;
  wire \u2_Display/lt155_c15 ;
  wire \u2_Display/lt155_c17 ;
  wire \u2_Display/lt155_c19 ;
  wire \u2_Display/lt155_c21 ;
  wire \u2_Display/lt155_c23 ;
  wire \u2_Display/lt155_c25 ;
  wire \u2_Display/lt155_c27 ;
  wire \u2_Display/lt155_c29 ;
  wire \u2_Display/lt155_c3 ;
  wire \u2_Display/lt155_c31 ;
  wire \u2_Display/lt155_c5 ;
  wire \u2_Display/lt155_c7 ;
  wire \u2_Display/lt155_c9 ;
  wire \u2_Display/lt156_c1 ;
  wire \u2_Display/lt156_c11 ;
  wire \u2_Display/lt156_c13 ;
  wire \u2_Display/lt156_c15 ;
  wire \u2_Display/lt156_c17 ;
  wire \u2_Display/lt156_c19 ;
  wire \u2_Display/lt156_c21 ;
  wire \u2_Display/lt156_c23 ;
  wire \u2_Display/lt156_c25 ;
  wire \u2_Display/lt156_c27 ;
  wire \u2_Display/lt156_c29 ;
  wire \u2_Display/lt156_c3 ;
  wire \u2_Display/lt156_c31 ;
  wire \u2_Display/lt156_c5 ;
  wire \u2_Display/lt156_c7 ;
  wire \u2_Display/lt156_c9 ;
  wire \u2_Display/lt157_c1 ;
  wire \u2_Display/lt157_c11 ;
  wire \u2_Display/lt157_c13 ;
  wire \u2_Display/lt157_c15 ;
  wire \u2_Display/lt157_c17 ;
  wire \u2_Display/lt157_c19 ;
  wire \u2_Display/lt157_c21 ;
  wire \u2_Display/lt157_c23 ;
  wire \u2_Display/lt157_c25 ;
  wire \u2_Display/lt157_c27 ;
  wire \u2_Display/lt157_c29 ;
  wire \u2_Display/lt157_c3 ;
  wire \u2_Display/lt157_c31 ;
  wire \u2_Display/lt157_c5 ;
  wire \u2_Display/lt157_c7 ;
  wire \u2_Display/lt157_c9 ;
  wire \u2_Display/lt158_c1 ;
  wire \u2_Display/lt158_c11 ;
  wire \u2_Display/lt158_c13 ;
  wire \u2_Display/lt158_c15 ;
  wire \u2_Display/lt158_c17 ;
  wire \u2_Display/lt158_c19 ;
  wire \u2_Display/lt158_c21 ;
  wire \u2_Display/lt158_c23 ;
  wire \u2_Display/lt158_c25 ;
  wire \u2_Display/lt158_c27 ;
  wire \u2_Display/lt158_c29 ;
  wire \u2_Display/lt158_c3 ;
  wire \u2_Display/lt158_c31 ;
  wire \u2_Display/lt158_c5 ;
  wire \u2_Display/lt158_c7 ;
  wire \u2_Display/lt158_c9 ;
  wire \u2_Display/lt159_c1 ;
  wire \u2_Display/lt159_c11 ;
  wire \u2_Display/lt159_c13 ;
  wire \u2_Display/lt159_c15 ;
  wire \u2_Display/lt159_c17 ;
  wire \u2_Display/lt159_c19 ;
  wire \u2_Display/lt159_c21 ;
  wire \u2_Display/lt159_c23 ;
  wire \u2_Display/lt159_c25 ;
  wire \u2_Display/lt159_c27 ;
  wire \u2_Display/lt159_c29 ;
  wire \u2_Display/lt159_c3 ;
  wire \u2_Display/lt159_c31 ;
  wire \u2_Display/lt159_c5 ;
  wire \u2_Display/lt159_c7 ;
  wire \u2_Display/lt159_c9 ;
  wire \u2_Display/lt160_c1 ;
  wire \u2_Display/lt160_c11 ;
  wire \u2_Display/lt160_c13 ;
  wire \u2_Display/lt160_c15 ;
  wire \u2_Display/lt160_c17 ;
  wire \u2_Display/lt160_c19 ;
  wire \u2_Display/lt160_c21 ;
  wire \u2_Display/lt160_c23 ;
  wire \u2_Display/lt160_c25 ;
  wire \u2_Display/lt160_c27 ;
  wire \u2_Display/lt160_c29 ;
  wire \u2_Display/lt160_c3 ;
  wire \u2_Display/lt160_c31 ;
  wire \u2_Display/lt160_c5 ;
  wire \u2_Display/lt160_c7 ;
  wire \u2_Display/lt160_c9 ;
  wire \u2_Display/lt161_c1 ;
  wire \u2_Display/lt161_c11 ;
  wire \u2_Display/lt161_c13 ;
  wire \u2_Display/lt161_c15 ;
  wire \u2_Display/lt161_c17 ;
  wire \u2_Display/lt161_c19 ;
  wire \u2_Display/lt161_c21 ;
  wire \u2_Display/lt161_c23 ;
  wire \u2_Display/lt161_c25 ;
  wire \u2_Display/lt161_c27 ;
  wire \u2_Display/lt161_c29 ;
  wire \u2_Display/lt161_c3 ;
  wire \u2_Display/lt161_c31 ;
  wire \u2_Display/lt161_c5 ;
  wire \u2_Display/lt161_c7 ;
  wire \u2_Display/lt161_c9 ;
  wire \u2_Display/lt162_c1 ;
  wire \u2_Display/lt162_c11 ;
  wire \u2_Display/lt162_c13 ;
  wire \u2_Display/lt162_c15 ;
  wire \u2_Display/lt162_c17 ;
  wire \u2_Display/lt162_c19 ;
  wire \u2_Display/lt162_c21 ;
  wire \u2_Display/lt162_c23 ;
  wire \u2_Display/lt162_c25 ;
  wire \u2_Display/lt162_c27 ;
  wire \u2_Display/lt162_c29 ;
  wire \u2_Display/lt162_c3 ;
  wire \u2_Display/lt162_c31 ;
  wire \u2_Display/lt162_c5 ;
  wire \u2_Display/lt162_c7 ;
  wire \u2_Display/lt162_c9 ;
  wire \u2_Display/lt163_c1 ;
  wire \u2_Display/lt163_c11 ;
  wire \u2_Display/lt163_c13 ;
  wire \u2_Display/lt163_c15 ;
  wire \u2_Display/lt163_c17 ;
  wire \u2_Display/lt163_c19 ;
  wire \u2_Display/lt163_c21 ;
  wire \u2_Display/lt163_c23 ;
  wire \u2_Display/lt163_c25 ;
  wire \u2_Display/lt163_c27 ;
  wire \u2_Display/lt163_c29 ;
  wire \u2_Display/lt163_c3 ;
  wire \u2_Display/lt163_c31 ;
  wire \u2_Display/lt163_c5 ;
  wire \u2_Display/lt163_c7 ;
  wire \u2_Display/lt163_c9 ;
  wire \u2_Display/lt164_c1 ;
  wire \u2_Display/lt164_c11 ;
  wire \u2_Display/lt164_c13 ;
  wire \u2_Display/lt164_c15 ;
  wire \u2_Display/lt164_c17 ;
  wire \u2_Display/lt164_c19 ;
  wire \u2_Display/lt164_c21 ;
  wire \u2_Display/lt164_c23 ;
  wire \u2_Display/lt164_c25 ;
  wire \u2_Display/lt164_c27 ;
  wire \u2_Display/lt164_c29 ;
  wire \u2_Display/lt164_c3 ;
  wire \u2_Display/lt164_c31 ;
  wire \u2_Display/lt164_c5 ;
  wire \u2_Display/lt164_c7 ;
  wire \u2_Display/lt164_c9 ;
  wire \u2_Display/lt165_c1 ;
  wire \u2_Display/lt165_c11 ;
  wire \u2_Display/lt165_c13 ;
  wire \u2_Display/lt165_c15 ;
  wire \u2_Display/lt165_c17 ;
  wire \u2_Display/lt165_c19 ;
  wire \u2_Display/lt165_c21 ;
  wire \u2_Display/lt165_c23 ;
  wire \u2_Display/lt165_c25 ;
  wire \u2_Display/lt165_c27 ;
  wire \u2_Display/lt165_c29 ;
  wire \u2_Display/lt165_c3 ;
  wire \u2_Display/lt165_c31 ;
  wire \u2_Display/lt165_c5 ;
  wire \u2_Display/lt165_c7 ;
  wire \u2_Display/lt165_c9 ;
  wire \u2_Display/lt166_c1 ;
  wire \u2_Display/lt166_c11 ;
  wire \u2_Display/lt166_c13 ;
  wire \u2_Display/lt166_c15 ;
  wire \u2_Display/lt166_c17 ;
  wire \u2_Display/lt166_c19 ;
  wire \u2_Display/lt166_c21 ;
  wire \u2_Display/lt166_c23 ;
  wire \u2_Display/lt166_c25 ;
  wire \u2_Display/lt166_c27 ;
  wire \u2_Display/lt166_c29 ;
  wire \u2_Display/lt166_c3 ;
  wire \u2_Display/lt166_c31 ;
  wire \u2_Display/lt166_c5 ;
  wire \u2_Display/lt166_c7 ;
  wire \u2_Display/lt166_c9 ;
  wire \u2_Display/lt167_c1 ;
  wire \u2_Display/lt167_c11 ;
  wire \u2_Display/lt167_c13 ;
  wire \u2_Display/lt167_c15 ;
  wire \u2_Display/lt167_c17 ;
  wire \u2_Display/lt167_c19 ;
  wire \u2_Display/lt167_c21 ;
  wire \u2_Display/lt167_c23 ;
  wire \u2_Display/lt167_c25 ;
  wire \u2_Display/lt167_c27 ;
  wire \u2_Display/lt167_c29 ;
  wire \u2_Display/lt167_c3 ;
  wire \u2_Display/lt167_c31 ;
  wire \u2_Display/lt167_c5 ;
  wire \u2_Display/lt167_c7 ;
  wire \u2_Display/lt167_c9 ;
  wire \u2_Display/lt168_c1 ;
  wire \u2_Display/lt168_c11 ;
  wire \u2_Display/lt168_c13 ;
  wire \u2_Display/lt168_c15 ;
  wire \u2_Display/lt168_c17 ;
  wire \u2_Display/lt168_c19 ;
  wire \u2_Display/lt168_c21 ;
  wire \u2_Display/lt168_c23 ;
  wire \u2_Display/lt168_c25 ;
  wire \u2_Display/lt168_c27 ;
  wire \u2_Display/lt168_c29 ;
  wire \u2_Display/lt168_c3 ;
  wire \u2_Display/lt168_c31 ;
  wire \u2_Display/lt168_c5 ;
  wire \u2_Display/lt168_c7 ;
  wire \u2_Display/lt168_c9 ;
  wire \u2_Display/lt169_c1 ;
  wire \u2_Display/lt169_c11 ;
  wire \u2_Display/lt169_c13 ;
  wire \u2_Display/lt169_c15 ;
  wire \u2_Display/lt169_c17 ;
  wire \u2_Display/lt169_c19 ;
  wire \u2_Display/lt169_c21 ;
  wire \u2_Display/lt169_c23 ;
  wire \u2_Display/lt169_c25 ;
  wire \u2_Display/lt169_c27 ;
  wire \u2_Display/lt169_c29 ;
  wire \u2_Display/lt169_c3 ;
  wire \u2_Display/lt169_c31 ;
  wire \u2_Display/lt169_c5 ;
  wire \u2_Display/lt169_c7 ;
  wire \u2_Display/lt169_c9 ;
  wire \u2_Display/lt170_c1 ;
  wire \u2_Display/lt170_c11 ;
  wire \u2_Display/lt170_c13 ;
  wire \u2_Display/lt170_c15 ;
  wire \u2_Display/lt170_c17 ;
  wire \u2_Display/lt170_c19 ;
  wire \u2_Display/lt170_c21 ;
  wire \u2_Display/lt170_c23 ;
  wire \u2_Display/lt170_c25 ;
  wire \u2_Display/lt170_c27 ;
  wire \u2_Display/lt170_c29 ;
  wire \u2_Display/lt170_c3 ;
  wire \u2_Display/lt170_c31 ;
  wire \u2_Display/lt170_c5 ;
  wire \u2_Display/lt170_c7 ;
  wire \u2_Display/lt170_c9 ;
  wire \u2_Display/lt171_c1 ;
  wire \u2_Display/lt171_c11 ;
  wire \u2_Display/lt171_c13 ;
  wire \u2_Display/lt171_c15 ;
  wire \u2_Display/lt171_c17 ;
  wire \u2_Display/lt171_c19 ;
  wire \u2_Display/lt171_c21 ;
  wire \u2_Display/lt171_c23 ;
  wire \u2_Display/lt171_c25 ;
  wire \u2_Display/lt171_c27 ;
  wire \u2_Display/lt171_c29 ;
  wire \u2_Display/lt171_c3 ;
  wire \u2_Display/lt171_c31 ;
  wire \u2_Display/lt171_c5 ;
  wire \u2_Display/lt171_c7 ;
  wire \u2_Display/lt171_c9 ;
  wire \u2_Display/lt172_c1 ;
  wire \u2_Display/lt172_c11 ;
  wire \u2_Display/lt172_c13 ;
  wire \u2_Display/lt172_c15 ;
  wire \u2_Display/lt172_c17 ;
  wire \u2_Display/lt172_c19 ;
  wire \u2_Display/lt172_c21 ;
  wire \u2_Display/lt172_c23 ;
  wire \u2_Display/lt172_c25 ;
  wire \u2_Display/lt172_c27 ;
  wire \u2_Display/lt172_c29 ;
  wire \u2_Display/lt172_c3 ;
  wire \u2_Display/lt172_c31 ;
  wire \u2_Display/lt172_c5 ;
  wire \u2_Display/lt172_c7 ;
  wire \u2_Display/lt172_c9 ;
  wire \u2_Display/lt173_c1 ;
  wire \u2_Display/lt173_c11 ;
  wire \u2_Display/lt173_c13 ;
  wire \u2_Display/lt173_c15 ;
  wire \u2_Display/lt173_c17 ;
  wire \u2_Display/lt173_c19 ;
  wire \u2_Display/lt173_c21 ;
  wire \u2_Display/lt173_c23 ;
  wire \u2_Display/lt173_c25 ;
  wire \u2_Display/lt173_c27 ;
  wire \u2_Display/lt173_c29 ;
  wire \u2_Display/lt173_c3 ;
  wire \u2_Display/lt173_c31 ;
  wire \u2_Display/lt173_c5 ;
  wire \u2_Display/lt173_c7 ;
  wire \u2_Display/lt173_c9 ;
  wire \u2_Display/lt174_c1 ;
  wire \u2_Display/lt174_c11 ;
  wire \u2_Display/lt174_c13 ;
  wire \u2_Display/lt174_c15 ;
  wire \u2_Display/lt174_c17 ;
  wire \u2_Display/lt174_c19 ;
  wire \u2_Display/lt174_c21 ;
  wire \u2_Display/lt174_c23 ;
  wire \u2_Display/lt174_c25 ;
  wire \u2_Display/lt174_c27 ;
  wire \u2_Display/lt174_c29 ;
  wire \u2_Display/lt174_c3 ;
  wire \u2_Display/lt174_c31 ;
  wire \u2_Display/lt174_c5 ;
  wire \u2_Display/lt174_c7 ;
  wire \u2_Display/lt174_c9 ;
  wire \u2_Display/lt175_c1 ;
  wire \u2_Display/lt175_c11 ;
  wire \u2_Display/lt175_c13 ;
  wire \u2_Display/lt175_c15 ;
  wire \u2_Display/lt175_c17 ;
  wire \u2_Display/lt175_c19 ;
  wire \u2_Display/lt175_c21 ;
  wire \u2_Display/lt175_c23 ;
  wire \u2_Display/lt175_c25 ;
  wire \u2_Display/lt175_c27 ;
  wire \u2_Display/lt175_c29 ;
  wire \u2_Display/lt175_c3 ;
  wire \u2_Display/lt175_c31 ;
  wire \u2_Display/lt175_c5 ;
  wire \u2_Display/lt175_c7 ;
  wire \u2_Display/lt175_c9 ;
  wire \u2_Display/lt176_c1 ;
  wire \u2_Display/lt176_c11 ;
  wire \u2_Display/lt176_c13 ;
  wire \u2_Display/lt176_c15 ;
  wire \u2_Display/lt176_c17 ;
  wire \u2_Display/lt176_c19 ;
  wire \u2_Display/lt176_c21 ;
  wire \u2_Display/lt176_c23 ;
  wire \u2_Display/lt176_c25 ;
  wire \u2_Display/lt176_c27 ;
  wire \u2_Display/lt176_c29 ;
  wire \u2_Display/lt176_c3 ;
  wire \u2_Display/lt176_c31 ;
  wire \u2_Display/lt176_c5 ;
  wire \u2_Display/lt176_c7 ;
  wire \u2_Display/lt176_c9 ;
  wire \u2_Display/lt1_c1 ;
  wire \u2_Display/lt1_c11 ;
  wire \u2_Display/lt1_c3 ;
  wire \u2_Display/lt1_c5 ;
  wire \u2_Display/lt1_c7 ;
  wire \u2_Display/lt1_c9 ;
  wire \u2_Display/lt22_c1 ;
  wire \u2_Display/lt22_c11 ;
  wire \u2_Display/lt22_c13 ;
  wire \u2_Display/lt22_c15 ;
  wire \u2_Display/lt22_c17 ;
  wire \u2_Display/lt22_c19 ;
  wire \u2_Display/lt22_c21 ;
  wire \u2_Display/lt22_c23 ;
  wire \u2_Display/lt22_c25 ;
  wire \u2_Display/lt22_c27 ;
  wire \u2_Display/lt22_c29 ;
  wire \u2_Display/lt22_c3 ;
  wire \u2_Display/lt22_c31 ;
  wire \u2_Display/lt22_c5 ;
  wire \u2_Display/lt22_c7 ;
  wire \u2_Display/lt22_c9 ;
  wire \u2_Display/lt23_c1 ;
  wire \u2_Display/lt23_c11 ;
  wire \u2_Display/lt23_c13 ;
  wire \u2_Display/lt23_c15 ;
  wire \u2_Display/lt23_c17 ;
  wire \u2_Display/lt23_c19 ;
  wire \u2_Display/lt23_c21 ;
  wire \u2_Display/lt23_c23 ;
  wire \u2_Display/lt23_c25 ;
  wire \u2_Display/lt23_c27 ;
  wire \u2_Display/lt23_c29 ;
  wire \u2_Display/lt23_c3 ;
  wire \u2_Display/lt23_c31 ;
  wire \u2_Display/lt23_c5 ;
  wire \u2_Display/lt23_c7 ;
  wire \u2_Display/lt23_c9 ;
  wire \u2_Display/lt24_c1 ;
  wire \u2_Display/lt24_c11 ;
  wire \u2_Display/lt24_c13 ;
  wire \u2_Display/lt24_c15 ;
  wire \u2_Display/lt24_c17 ;
  wire \u2_Display/lt24_c19 ;
  wire \u2_Display/lt24_c21 ;
  wire \u2_Display/lt24_c23 ;
  wire \u2_Display/lt24_c25 ;
  wire \u2_Display/lt24_c27 ;
  wire \u2_Display/lt24_c29 ;
  wire \u2_Display/lt24_c3 ;
  wire \u2_Display/lt24_c31 ;
  wire \u2_Display/lt24_c5 ;
  wire \u2_Display/lt24_c7 ;
  wire \u2_Display/lt24_c9 ;
  wire \u2_Display/lt25_c1 ;
  wire \u2_Display/lt25_c11 ;
  wire \u2_Display/lt25_c13 ;
  wire \u2_Display/lt25_c15 ;
  wire \u2_Display/lt25_c17 ;
  wire \u2_Display/lt25_c19 ;
  wire \u2_Display/lt25_c21 ;
  wire \u2_Display/lt25_c23 ;
  wire \u2_Display/lt25_c25 ;
  wire \u2_Display/lt25_c27 ;
  wire \u2_Display/lt25_c29 ;
  wire \u2_Display/lt25_c3 ;
  wire \u2_Display/lt25_c31 ;
  wire \u2_Display/lt25_c5 ;
  wire \u2_Display/lt25_c7 ;
  wire \u2_Display/lt25_c9 ;
  wire \u2_Display/lt26_c1 ;
  wire \u2_Display/lt26_c11 ;
  wire \u2_Display/lt26_c13 ;
  wire \u2_Display/lt26_c15 ;
  wire \u2_Display/lt26_c17 ;
  wire \u2_Display/lt26_c19 ;
  wire \u2_Display/lt26_c21 ;
  wire \u2_Display/lt26_c23 ;
  wire \u2_Display/lt26_c25 ;
  wire \u2_Display/lt26_c27 ;
  wire \u2_Display/lt26_c29 ;
  wire \u2_Display/lt26_c3 ;
  wire \u2_Display/lt26_c31 ;
  wire \u2_Display/lt26_c5 ;
  wire \u2_Display/lt26_c7 ;
  wire \u2_Display/lt26_c9 ;
  wire \u2_Display/lt27_c1 ;
  wire \u2_Display/lt27_c11 ;
  wire \u2_Display/lt27_c13 ;
  wire \u2_Display/lt27_c15 ;
  wire \u2_Display/lt27_c17 ;
  wire \u2_Display/lt27_c19 ;
  wire \u2_Display/lt27_c21 ;
  wire \u2_Display/lt27_c23 ;
  wire \u2_Display/lt27_c25 ;
  wire \u2_Display/lt27_c27 ;
  wire \u2_Display/lt27_c29 ;
  wire \u2_Display/lt27_c3 ;
  wire \u2_Display/lt27_c31 ;
  wire \u2_Display/lt27_c5 ;
  wire \u2_Display/lt27_c7 ;
  wire \u2_Display/lt27_c9 ;
  wire \u2_Display/lt28_c1 ;
  wire \u2_Display/lt28_c11 ;
  wire \u2_Display/lt28_c13 ;
  wire \u2_Display/lt28_c15 ;
  wire \u2_Display/lt28_c17 ;
  wire \u2_Display/lt28_c19 ;
  wire \u2_Display/lt28_c21 ;
  wire \u2_Display/lt28_c23 ;
  wire \u2_Display/lt28_c25 ;
  wire \u2_Display/lt28_c27 ;
  wire \u2_Display/lt28_c29 ;
  wire \u2_Display/lt28_c3 ;
  wire \u2_Display/lt28_c31 ;
  wire \u2_Display/lt28_c5 ;
  wire \u2_Display/lt28_c7 ;
  wire \u2_Display/lt28_c9 ;
  wire \u2_Display/lt29_c1 ;
  wire \u2_Display/lt29_c11 ;
  wire \u2_Display/lt29_c13 ;
  wire \u2_Display/lt29_c15 ;
  wire \u2_Display/lt29_c17 ;
  wire \u2_Display/lt29_c19 ;
  wire \u2_Display/lt29_c21 ;
  wire \u2_Display/lt29_c23 ;
  wire \u2_Display/lt29_c25 ;
  wire \u2_Display/lt29_c27 ;
  wire \u2_Display/lt29_c29 ;
  wire \u2_Display/lt29_c3 ;
  wire \u2_Display/lt29_c31 ;
  wire \u2_Display/lt29_c5 ;
  wire \u2_Display/lt29_c7 ;
  wire \u2_Display/lt29_c9 ;
  wire \u2_Display/lt2_2_c1 ;
  wire \u2_Display/lt2_2_c11 ;
  wire \u2_Display/lt2_2_c3 ;
  wire \u2_Display/lt2_2_c5 ;
  wire \u2_Display/lt2_2_c7 ;
  wire \u2_Display/lt2_2_c9 ;
  wire \u2_Display/lt30_c1 ;
  wire \u2_Display/lt30_c11 ;
  wire \u2_Display/lt30_c13 ;
  wire \u2_Display/lt30_c15 ;
  wire \u2_Display/lt30_c17 ;
  wire \u2_Display/lt30_c19 ;
  wire \u2_Display/lt30_c21 ;
  wire \u2_Display/lt30_c23 ;
  wire \u2_Display/lt30_c25 ;
  wire \u2_Display/lt30_c27 ;
  wire \u2_Display/lt30_c29 ;
  wire \u2_Display/lt30_c3 ;
  wire \u2_Display/lt30_c31 ;
  wire \u2_Display/lt30_c5 ;
  wire \u2_Display/lt30_c7 ;
  wire \u2_Display/lt30_c9 ;
  wire \u2_Display/lt31_c1 ;
  wire \u2_Display/lt31_c11 ;
  wire \u2_Display/lt31_c13 ;
  wire \u2_Display/lt31_c15 ;
  wire \u2_Display/lt31_c17 ;
  wire \u2_Display/lt31_c19 ;
  wire \u2_Display/lt31_c21 ;
  wire \u2_Display/lt31_c23 ;
  wire \u2_Display/lt31_c25 ;
  wire \u2_Display/lt31_c27 ;
  wire \u2_Display/lt31_c29 ;
  wire \u2_Display/lt31_c3 ;
  wire \u2_Display/lt31_c31 ;
  wire \u2_Display/lt31_c5 ;
  wire \u2_Display/lt31_c7 ;
  wire \u2_Display/lt31_c9 ;
  wire \u2_Display/lt32_c1 ;
  wire \u2_Display/lt32_c11 ;
  wire \u2_Display/lt32_c13 ;
  wire \u2_Display/lt32_c15 ;
  wire \u2_Display/lt32_c17 ;
  wire \u2_Display/lt32_c19 ;
  wire \u2_Display/lt32_c21 ;
  wire \u2_Display/lt32_c23 ;
  wire \u2_Display/lt32_c25 ;
  wire \u2_Display/lt32_c27 ;
  wire \u2_Display/lt32_c29 ;
  wire \u2_Display/lt32_c3 ;
  wire \u2_Display/lt32_c31 ;
  wire \u2_Display/lt32_c5 ;
  wire \u2_Display/lt32_c7 ;
  wire \u2_Display/lt32_c9 ;
  wire \u2_Display/lt33_c1 ;
  wire \u2_Display/lt33_c11 ;
  wire \u2_Display/lt33_c13 ;
  wire \u2_Display/lt33_c15 ;
  wire \u2_Display/lt33_c17 ;
  wire \u2_Display/lt33_c19 ;
  wire \u2_Display/lt33_c21 ;
  wire \u2_Display/lt33_c23 ;
  wire \u2_Display/lt33_c25 ;
  wire \u2_Display/lt33_c27 ;
  wire \u2_Display/lt33_c29 ;
  wire \u2_Display/lt33_c3 ;
  wire \u2_Display/lt33_c31 ;
  wire \u2_Display/lt33_c5 ;
  wire \u2_Display/lt33_c7 ;
  wire \u2_Display/lt33_c9 ;
  wire \u2_Display/lt34_c1 ;
  wire \u2_Display/lt34_c11 ;
  wire \u2_Display/lt34_c13 ;
  wire \u2_Display/lt34_c15 ;
  wire \u2_Display/lt34_c17 ;
  wire \u2_Display/lt34_c19 ;
  wire \u2_Display/lt34_c21 ;
  wire \u2_Display/lt34_c23 ;
  wire \u2_Display/lt34_c25 ;
  wire \u2_Display/lt34_c27 ;
  wire \u2_Display/lt34_c29 ;
  wire \u2_Display/lt34_c3 ;
  wire \u2_Display/lt34_c31 ;
  wire \u2_Display/lt34_c5 ;
  wire \u2_Display/lt34_c7 ;
  wire \u2_Display/lt34_c9 ;
  wire \u2_Display/lt35_c1 ;
  wire \u2_Display/lt35_c11 ;
  wire \u2_Display/lt35_c13 ;
  wire \u2_Display/lt35_c15 ;
  wire \u2_Display/lt35_c17 ;
  wire \u2_Display/lt35_c19 ;
  wire \u2_Display/lt35_c21 ;
  wire \u2_Display/lt35_c23 ;
  wire \u2_Display/lt35_c25 ;
  wire \u2_Display/lt35_c27 ;
  wire \u2_Display/lt35_c29 ;
  wire \u2_Display/lt35_c3 ;
  wire \u2_Display/lt35_c31 ;
  wire \u2_Display/lt35_c5 ;
  wire \u2_Display/lt35_c7 ;
  wire \u2_Display/lt35_c9 ;
  wire \u2_Display/lt36_c1 ;
  wire \u2_Display/lt36_c11 ;
  wire \u2_Display/lt36_c13 ;
  wire \u2_Display/lt36_c15 ;
  wire \u2_Display/lt36_c17 ;
  wire \u2_Display/lt36_c19 ;
  wire \u2_Display/lt36_c21 ;
  wire \u2_Display/lt36_c23 ;
  wire \u2_Display/lt36_c25 ;
  wire \u2_Display/lt36_c27 ;
  wire \u2_Display/lt36_c29 ;
  wire \u2_Display/lt36_c3 ;
  wire \u2_Display/lt36_c31 ;
  wire \u2_Display/lt36_c5 ;
  wire \u2_Display/lt36_c7 ;
  wire \u2_Display/lt36_c9 ;
  wire \u2_Display/lt37_c1 ;
  wire \u2_Display/lt37_c11 ;
  wire \u2_Display/lt37_c13 ;
  wire \u2_Display/lt37_c15 ;
  wire \u2_Display/lt37_c17 ;
  wire \u2_Display/lt37_c19 ;
  wire \u2_Display/lt37_c21 ;
  wire \u2_Display/lt37_c23 ;
  wire \u2_Display/lt37_c25 ;
  wire \u2_Display/lt37_c27 ;
  wire \u2_Display/lt37_c29 ;
  wire \u2_Display/lt37_c3 ;
  wire \u2_Display/lt37_c31 ;
  wire \u2_Display/lt37_c5 ;
  wire \u2_Display/lt37_c7 ;
  wire \u2_Display/lt37_c9 ;
  wire \u2_Display/lt38_c1 ;
  wire \u2_Display/lt38_c11 ;
  wire \u2_Display/lt38_c13 ;
  wire \u2_Display/lt38_c15 ;
  wire \u2_Display/lt38_c17 ;
  wire \u2_Display/lt38_c19 ;
  wire \u2_Display/lt38_c21 ;
  wire \u2_Display/lt38_c23 ;
  wire \u2_Display/lt38_c25 ;
  wire \u2_Display/lt38_c27 ;
  wire \u2_Display/lt38_c29 ;
  wire \u2_Display/lt38_c3 ;
  wire \u2_Display/lt38_c31 ;
  wire \u2_Display/lt38_c5 ;
  wire \u2_Display/lt38_c7 ;
  wire \u2_Display/lt38_c9 ;
  wire \u2_Display/lt39_c1 ;
  wire \u2_Display/lt39_c11 ;
  wire \u2_Display/lt39_c13 ;
  wire \u2_Display/lt39_c15 ;
  wire \u2_Display/lt39_c17 ;
  wire \u2_Display/lt39_c19 ;
  wire \u2_Display/lt39_c21 ;
  wire \u2_Display/lt39_c23 ;
  wire \u2_Display/lt39_c25 ;
  wire \u2_Display/lt39_c27 ;
  wire \u2_Display/lt39_c29 ;
  wire \u2_Display/lt39_c3 ;
  wire \u2_Display/lt39_c31 ;
  wire \u2_Display/lt39_c5 ;
  wire \u2_Display/lt39_c7 ;
  wire \u2_Display/lt39_c9 ;
  wire \u2_Display/lt3_c1 ;
  wire \u2_Display/lt3_c11 ;
  wire \u2_Display/lt3_c3 ;
  wire \u2_Display/lt3_c5 ;
  wire \u2_Display/lt3_c7 ;
  wire \u2_Display/lt3_c9 ;
  wire \u2_Display/lt40_c1 ;
  wire \u2_Display/lt40_c11 ;
  wire \u2_Display/lt40_c13 ;
  wire \u2_Display/lt40_c15 ;
  wire \u2_Display/lt40_c17 ;
  wire \u2_Display/lt40_c19 ;
  wire \u2_Display/lt40_c21 ;
  wire \u2_Display/lt40_c23 ;
  wire \u2_Display/lt40_c25 ;
  wire \u2_Display/lt40_c27 ;
  wire \u2_Display/lt40_c29 ;
  wire \u2_Display/lt40_c3 ;
  wire \u2_Display/lt40_c31 ;
  wire \u2_Display/lt40_c5 ;
  wire \u2_Display/lt40_c7 ;
  wire \u2_Display/lt40_c9 ;
  wire \u2_Display/lt41_c1 ;
  wire \u2_Display/lt41_c11 ;
  wire \u2_Display/lt41_c13 ;
  wire \u2_Display/lt41_c15 ;
  wire \u2_Display/lt41_c17 ;
  wire \u2_Display/lt41_c19 ;
  wire \u2_Display/lt41_c21 ;
  wire \u2_Display/lt41_c23 ;
  wire \u2_Display/lt41_c25 ;
  wire \u2_Display/lt41_c27 ;
  wire \u2_Display/lt41_c29 ;
  wire \u2_Display/lt41_c3 ;
  wire \u2_Display/lt41_c31 ;
  wire \u2_Display/lt41_c5 ;
  wire \u2_Display/lt41_c7 ;
  wire \u2_Display/lt41_c9 ;
  wire \u2_Display/lt42_c1 ;
  wire \u2_Display/lt42_c11 ;
  wire \u2_Display/lt42_c13 ;
  wire \u2_Display/lt42_c15 ;
  wire \u2_Display/lt42_c17 ;
  wire \u2_Display/lt42_c19 ;
  wire \u2_Display/lt42_c21 ;
  wire \u2_Display/lt42_c23 ;
  wire \u2_Display/lt42_c25 ;
  wire \u2_Display/lt42_c27 ;
  wire \u2_Display/lt42_c29 ;
  wire \u2_Display/lt42_c3 ;
  wire \u2_Display/lt42_c31 ;
  wire \u2_Display/lt42_c5 ;
  wire \u2_Display/lt42_c7 ;
  wire \u2_Display/lt42_c9 ;
  wire \u2_Display/lt43_c1 ;
  wire \u2_Display/lt43_c11 ;
  wire \u2_Display/lt43_c13 ;
  wire \u2_Display/lt43_c15 ;
  wire \u2_Display/lt43_c17 ;
  wire \u2_Display/lt43_c19 ;
  wire \u2_Display/lt43_c21 ;
  wire \u2_Display/lt43_c23 ;
  wire \u2_Display/lt43_c25 ;
  wire \u2_Display/lt43_c27 ;
  wire \u2_Display/lt43_c29 ;
  wire \u2_Display/lt43_c3 ;
  wire \u2_Display/lt43_c31 ;
  wire \u2_Display/lt43_c5 ;
  wire \u2_Display/lt43_c7 ;
  wire \u2_Display/lt43_c9 ;
  wire \u2_Display/lt44_c1 ;
  wire \u2_Display/lt44_c11 ;
  wire \u2_Display/lt44_c13 ;
  wire \u2_Display/lt44_c15 ;
  wire \u2_Display/lt44_c17 ;
  wire \u2_Display/lt44_c19 ;
  wire \u2_Display/lt44_c21 ;
  wire \u2_Display/lt44_c23 ;
  wire \u2_Display/lt44_c25 ;
  wire \u2_Display/lt44_c27 ;
  wire \u2_Display/lt44_c29 ;
  wire \u2_Display/lt44_c3 ;
  wire \u2_Display/lt44_c31 ;
  wire \u2_Display/lt44_c5 ;
  wire \u2_Display/lt44_c7 ;
  wire \u2_Display/lt44_c9 ;
  wire \u2_Display/lt4_2_c1 ;
  wire \u2_Display/lt4_2_c11 ;
  wire \u2_Display/lt4_2_c3 ;
  wire \u2_Display/lt4_2_c5 ;
  wire \u2_Display/lt4_2_c7 ;
  wire \u2_Display/lt4_2_c9 ;
  wire \u2_Display/lt55_c1 ;
  wire \u2_Display/lt55_c11 ;
  wire \u2_Display/lt55_c13 ;
  wire \u2_Display/lt55_c15 ;
  wire \u2_Display/lt55_c17 ;
  wire \u2_Display/lt55_c19 ;
  wire \u2_Display/lt55_c21 ;
  wire \u2_Display/lt55_c23 ;
  wire \u2_Display/lt55_c25 ;
  wire \u2_Display/lt55_c27 ;
  wire \u2_Display/lt55_c29 ;
  wire \u2_Display/lt55_c3 ;
  wire \u2_Display/lt55_c31 ;
  wire \u2_Display/lt55_c5 ;
  wire \u2_Display/lt55_c7 ;
  wire \u2_Display/lt55_c9 ;
  wire \u2_Display/lt56_c1 ;
  wire \u2_Display/lt56_c11 ;
  wire \u2_Display/lt56_c13 ;
  wire \u2_Display/lt56_c15 ;
  wire \u2_Display/lt56_c17 ;
  wire \u2_Display/lt56_c19 ;
  wire \u2_Display/lt56_c21 ;
  wire \u2_Display/lt56_c23 ;
  wire \u2_Display/lt56_c25 ;
  wire \u2_Display/lt56_c27 ;
  wire \u2_Display/lt56_c29 ;
  wire \u2_Display/lt56_c3 ;
  wire \u2_Display/lt56_c31 ;
  wire \u2_Display/lt56_c5 ;
  wire \u2_Display/lt56_c7 ;
  wire \u2_Display/lt56_c9 ;
  wire \u2_Display/lt57_c1 ;
  wire \u2_Display/lt57_c11 ;
  wire \u2_Display/lt57_c13 ;
  wire \u2_Display/lt57_c15 ;
  wire \u2_Display/lt57_c17 ;
  wire \u2_Display/lt57_c19 ;
  wire \u2_Display/lt57_c21 ;
  wire \u2_Display/lt57_c23 ;
  wire \u2_Display/lt57_c25 ;
  wire \u2_Display/lt57_c27 ;
  wire \u2_Display/lt57_c29 ;
  wire \u2_Display/lt57_c3 ;
  wire \u2_Display/lt57_c31 ;
  wire \u2_Display/lt57_c5 ;
  wire \u2_Display/lt57_c7 ;
  wire \u2_Display/lt57_c9 ;
  wire \u2_Display/lt58_c1 ;
  wire \u2_Display/lt58_c11 ;
  wire \u2_Display/lt58_c13 ;
  wire \u2_Display/lt58_c15 ;
  wire \u2_Display/lt58_c17 ;
  wire \u2_Display/lt58_c19 ;
  wire \u2_Display/lt58_c21 ;
  wire \u2_Display/lt58_c23 ;
  wire \u2_Display/lt58_c25 ;
  wire \u2_Display/lt58_c27 ;
  wire \u2_Display/lt58_c29 ;
  wire \u2_Display/lt58_c3 ;
  wire \u2_Display/lt58_c31 ;
  wire \u2_Display/lt58_c5 ;
  wire \u2_Display/lt58_c7 ;
  wire \u2_Display/lt58_c9 ;
  wire \u2_Display/lt59_c1 ;
  wire \u2_Display/lt59_c11 ;
  wire \u2_Display/lt59_c13 ;
  wire \u2_Display/lt59_c15 ;
  wire \u2_Display/lt59_c17 ;
  wire \u2_Display/lt59_c19 ;
  wire \u2_Display/lt59_c21 ;
  wire \u2_Display/lt59_c23 ;
  wire \u2_Display/lt59_c25 ;
  wire \u2_Display/lt59_c27 ;
  wire \u2_Display/lt59_c29 ;
  wire \u2_Display/lt59_c3 ;
  wire \u2_Display/lt59_c31 ;
  wire \u2_Display/lt59_c5 ;
  wire \u2_Display/lt59_c7 ;
  wire \u2_Display/lt59_c9 ;
  wire \u2_Display/lt5_2_c1 ;
  wire \u2_Display/lt5_2_c11 ;
  wire \u2_Display/lt5_2_c13 ;
  wire \u2_Display/lt5_2_c3 ;
  wire \u2_Display/lt5_2_c5 ;
  wire \u2_Display/lt5_2_c7 ;
  wire \u2_Display/lt5_2_c9 ;
  wire \u2_Display/lt60_c1 ;
  wire \u2_Display/lt60_c11 ;
  wire \u2_Display/lt60_c13 ;
  wire \u2_Display/lt60_c15 ;
  wire \u2_Display/lt60_c17 ;
  wire \u2_Display/lt60_c19 ;
  wire \u2_Display/lt60_c21 ;
  wire \u2_Display/lt60_c23 ;
  wire \u2_Display/lt60_c25 ;
  wire \u2_Display/lt60_c27 ;
  wire \u2_Display/lt60_c29 ;
  wire \u2_Display/lt60_c3 ;
  wire \u2_Display/lt60_c31 ;
  wire \u2_Display/lt60_c5 ;
  wire \u2_Display/lt60_c7 ;
  wire \u2_Display/lt60_c9 ;
  wire \u2_Display/lt61_c1 ;
  wire \u2_Display/lt61_c11 ;
  wire \u2_Display/lt61_c13 ;
  wire \u2_Display/lt61_c15 ;
  wire \u2_Display/lt61_c17 ;
  wire \u2_Display/lt61_c19 ;
  wire \u2_Display/lt61_c21 ;
  wire \u2_Display/lt61_c23 ;
  wire \u2_Display/lt61_c25 ;
  wire \u2_Display/lt61_c27 ;
  wire \u2_Display/lt61_c29 ;
  wire \u2_Display/lt61_c3 ;
  wire \u2_Display/lt61_c31 ;
  wire \u2_Display/lt61_c5 ;
  wire \u2_Display/lt61_c7 ;
  wire \u2_Display/lt61_c9 ;
  wire \u2_Display/lt62_c1 ;
  wire \u2_Display/lt62_c11 ;
  wire \u2_Display/lt62_c13 ;
  wire \u2_Display/lt62_c15 ;
  wire \u2_Display/lt62_c17 ;
  wire \u2_Display/lt62_c19 ;
  wire \u2_Display/lt62_c21 ;
  wire \u2_Display/lt62_c23 ;
  wire \u2_Display/lt62_c25 ;
  wire \u2_Display/lt62_c27 ;
  wire \u2_Display/lt62_c29 ;
  wire \u2_Display/lt62_c3 ;
  wire \u2_Display/lt62_c31 ;
  wire \u2_Display/lt62_c5 ;
  wire \u2_Display/lt62_c7 ;
  wire \u2_Display/lt62_c9 ;
  wire \u2_Display/lt63_c1 ;
  wire \u2_Display/lt63_c11 ;
  wire \u2_Display/lt63_c13 ;
  wire \u2_Display/lt63_c15 ;
  wire \u2_Display/lt63_c17 ;
  wire \u2_Display/lt63_c19 ;
  wire \u2_Display/lt63_c21 ;
  wire \u2_Display/lt63_c23 ;
  wire \u2_Display/lt63_c25 ;
  wire \u2_Display/lt63_c27 ;
  wire \u2_Display/lt63_c29 ;
  wire \u2_Display/lt63_c3 ;
  wire \u2_Display/lt63_c31 ;
  wire \u2_Display/lt63_c5 ;
  wire \u2_Display/lt63_c7 ;
  wire \u2_Display/lt63_c9 ;
  wire \u2_Display/lt64_c1 ;
  wire \u2_Display/lt64_c11 ;
  wire \u2_Display/lt64_c13 ;
  wire \u2_Display/lt64_c15 ;
  wire \u2_Display/lt64_c17 ;
  wire \u2_Display/lt64_c19 ;
  wire \u2_Display/lt64_c21 ;
  wire \u2_Display/lt64_c23 ;
  wire \u2_Display/lt64_c25 ;
  wire \u2_Display/lt64_c27 ;
  wire \u2_Display/lt64_c29 ;
  wire \u2_Display/lt64_c3 ;
  wire \u2_Display/lt64_c31 ;
  wire \u2_Display/lt64_c5 ;
  wire \u2_Display/lt64_c7 ;
  wire \u2_Display/lt64_c9 ;
  wire \u2_Display/lt65_c1 ;
  wire \u2_Display/lt65_c11 ;
  wire \u2_Display/lt65_c13 ;
  wire \u2_Display/lt65_c15 ;
  wire \u2_Display/lt65_c17 ;
  wire \u2_Display/lt65_c19 ;
  wire \u2_Display/lt65_c21 ;
  wire \u2_Display/lt65_c23 ;
  wire \u2_Display/lt65_c25 ;
  wire \u2_Display/lt65_c27 ;
  wire \u2_Display/lt65_c29 ;
  wire \u2_Display/lt65_c3 ;
  wire \u2_Display/lt65_c31 ;
  wire \u2_Display/lt65_c5 ;
  wire \u2_Display/lt65_c7 ;
  wire \u2_Display/lt65_c9 ;
  wire \u2_Display/lt66_c1 ;
  wire \u2_Display/lt66_c11 ;
  wire \u2_Display/lt66_c13 ;
  wire \u2_Display/lt66_c15 ;
  wire \u2_Display/lt66_c17 ;
  wire \u2_Display/lt66_c19 ;
  wire \u2_Display/lt66_c21 ;
  wire \u2_Display/lt66_c23 ;
  wire \u2_Display/lt66_c25 ;
  wire \u2_Display/lt66_c27 ;
  wire \u2_Display/lt66_c29 ;
  wire \u2_Display/lt66_c3 ;
  wire \u2_Display/lt66_c31 ;
  wire \u2_Display/lt66_c5 ;
  wire \u2_Display/lt66_c7 ;
  wire \u2_Display/lt66_c9 ;
  wire \u2_Display/lt67_c1 ;
  wire \u2_Display/lt67_c11 ;
  wire \u2_Display/lt67_c13 ;
  wire \u2_Display/lt67_c15 ;
  wire \u2_Display/lt67_c17 ;
  wire \u2_Display/lt67_c19 ;
  wire \u2_Display/lt67_c21 ;
  wire \u2_Display/lt67_c23 ;
  wire \u2_Display/lt67_c25 ;
  wire \u2_Display/lt67_c27 ;
  wire \u2_Display/lt67_c29 ;
  wire \u2_Display/lt67_c3 ;
  wire \u2_Display/lt67_c31 ;
  wire \u2_Display/lt67_c5 ;
  wire \u2_Display/lt67_c7 ;
  wire \u2_Display/lt67_c9 ;
  wire \u2_Display/lt68_c1 ;
  wire \u2_Display/lt68_c11 ;
  wire \u2_Display/lt68_c13 ;
  wire \u2_Display/lt68_c15 ;
  wire \u2_Display/lt68_c17 ;
  wire \u2_Display/lt68_c19 ;
  wire \u2_Display/lt68_c21 ;
  wire \u2_Display/lt68_c23 ;
  wire \u2_Display/lt68_c25 ;
  wire \u2_Display/lt68_c27 ;
  wire \u2_Display/lt68_c29 ;
  wire \u2_Display/lt68_c3 ;
  wire \u2_Display/lt68_c31 ;
  wire \u2_Display/lt68_c5 ;
  wire \u2_Display/lt68_c7 ;
  wire \u2_Display/lt68_c9 ;
  wire \u2_Display/lt69_c1 ;
  wire \u2_Display/lt69_c11 ;
  wire \u2_Display/lt69_c13 ;
  wire \u2_Display/lt69_c15 ;
  wire \u2_Display/lt69_c17 ;
  wire \u2_Display/lt69_c19 ;
  wire \u2_Display/lt69_c21 ;
  wire \u2_Display/lt69_c23 ;
  wire \u2_Display/lt69_c25 ;
  wire \u2_Display/lt69_c27 ;
  wire \u2_Display/lt69_c29 ;
  wire \u2_Display/lt69_c3 ;
  wire \u2_Display/lt69_c31 ;
  wire \u2_Display/lt69_c5 ;
  wire \u2_Display/lt69_c7 ;
  wire \u2_Display/lt69_c9 ;
  wire \u2_Display/lt6_2_c1 ;
  wire \u2_Display/lt6_2_c11 ;
  wire \u2_Display/lt6_2_c3 ;
  wire \u2_Display/lt6_2_c5 ;
  wire \u2_Display/lt6_2_c7 ;
  wire \u2_Display/lt6_2_c9 ;
  wire \u2_Display/lt70_c1 ;
  wire \u2_Display/lt70_c11 ;
  wire \u2_Display/lt70_c13 ;
  wire \u2_Display/lt70_c15 ;
  wire \u2_Display/lt70_c17 ;
  wire \u2_Display/lt70_c19 ;
  wire \u2_Display/lt70_c21 ;
  wire \u2_Display/lt70_c23 ;
  wire \u2_Display/lt70_c25 ;
  wire \u2_Display/lt70_c27 ;
  wire \u2_Display/lt70_c29 ;
  wire \u2_Display/lt70_c3 ;
  wire \u2_Display/lt70_c31 ;
  wire \u2_Display/lt70_c5 ;
  wire \u2_Display/lt70_c7 ;
  wire \u2_Display/lt70_c9 ;
  wire \u2_Display/lt71_c1 ;
  wire \u2_Display/lt71_c11 ;
  wire \u2_Display/lt71_c13 ;
  wire \u2_Display/lt71_c15 ;
  wire \u2_Display/lt71_c17 ;
  wire \u2_Display/lt71_c19 ;
  wire \u2_Display/lt71_c21 ;
  wire \u2_Display/lt71_c23 ;
  wire \u2_Display/lt71_c25 ;
  wire \u2_Display/lt71_c27 ;
  wire \u2_Display/lt71_c29 ;
  wire \u2_Display/lt71_c3 ;
  wire \u2_Display/lt71_c31 ;
  wire \u2_Display/lt71_c5 ;
  wire \u2_Display/lt71_c7 ;
  wire \u2_Display/lt71_c9 ;
  wire \u2_Display/lt72_c1 ;
  wire \u2_Display/lt72_c11 ;
  wire \u2_Display/lt72_c13 ;
  wire \u2_Display/lt72_c15 ;
  wire \u2_Display/lt72_c17 ;
  wire \u2_Display/lt72_c19 ;
  wire \u2_Display/lt72_c21 ;
  wire \u2_Display/lt72_c23 ;
  wire \u2_Display/lt72_c25 ;
  wire \u2_Display/lt72_c27 ;
  wire \u2_Display/lt72_c29 ;
  wire \u2_Display/lt72_c3 ;
  wire \u2_Display/lt72_c31 ;
  wire \u2_Display/lt72_c5 ;
  wire \u2_Display/lt72_c7 ;
  wire \u2_Display/lt72_c9 ;
  wire \u2_Display/lt73_c1 ;
  wire \u2_Display/lt73_c11 ;
  wire \u2_Display/lt73_c13 ;
  wire \u2_Display/lt73_c15 ;
  wire \u2_Display/lt73_c17 ;
  wire \u2_Display/lt73_c19 ;
  wire \u2_Display/lt73_c21 ;
  wire \u2_Display/lt73_c23 ;
  wire \u2_Display/lt73_c25 ;
  wire \u2_Display/lt73_c27 ;
  wire \u2_Display/lt73_c29 ;
  wire \u2_Display/lt73_c3 ;
  wire \u2_Display/lt73_c31 ;
  wire \u2_Display/lt73_c5 ;
  wire \u2_Display/lt73_c7 ;
  wire \u2_Display/lt73_c9 ;
  wire \u2_Display/lt74_c1 ;
  wire \u2_Display/lt74_c11 ;
  wire \u2_Display/lt74_c13 ;
  wire \u2_Display/lt74_c15 ;
  wire \u2_Display/lt74_c17 ;
  wire \u2_Display/lt74_c19 ;
  wire \u2_Display/lt74_c21 ;
  wire \u2_Display/lt74_c23 ;
  wire \u2_Display/lt74_c25 ;
  wire \u2_Display/lt74_c27 ;
  wire \u2_Display/lt74_c29 ;
  wire \u2_Display/lt74_c3 ;
  wire \u2_Display/lt74_c31 ;
  wire \u2_Display/lt74_c5 ;
  wire \u2_Display/lt74_c7 ;
  wire \u2_Display/lt74_c9 ;
  wire \u2_Display/lt75_c1 ;
  wire \u2_Display/lt75_c11 ;
  wire \u2_Display/lt75_c13 ;
  wire \u2_Display/lt75_c15 ;
  wire \u2_Display/lt75_c17 ;
  wire \u2_Display/lt75_c19 ;
  wire \u2_Display/lt75_c21 ;
  wire \u2_Display/lt75_c23 ;
  wire \u2_Display/lt75_c25 ;
  wire \u2_Display/lt75_c27 ;
  wire \u2_Display/lt75_c29 ;
  wire \u2_Display/lt75_c3 ;
  wire \u2_Display/lt75_c31 ;
  wire \u2_Display/lt75_c5 ;
  wire \u2_Display/lt75_c7 ;
  wire \u2_Display/lt75_c9 ;
  wire \u2_Display/lt76_c1 ;
  wire \u2_Display/lt76_c11 ;
  wire \u2_Display/lt76_c13 ;
  wire \u2_Display/lt76_c15 ;
  wire \u2_Display/lt76_c17 ;
  wire \u2_Display/lt76_c19 ;
  wire \u2_Display/lt76_c21 ;
  wire \u2_Display/lt76_c23 ;
  wire \u2_Display/lt76_c25 ;
  wire \u2_Display/lt76_c27 ;
  wire \u2_Display/lt76_c29 ;
  wire \u2_Display/lt76_c3 ;
  wire \u2_Display/lt76_c31 ;
  wire \u2_Display/lt76_c5 ;
  wire \u2_Display/lt76_c7 ;
  wire \u2_Display/lt76_c9 ;
  wire \u2_Display/lt77_c1 ;
  wire \u2_Display/lt77_c11 ;
  wire \u2_Display/lt77_c13 ;
  wire \u2_Display/lt77_c15 ;
  wire \u2_Display/lt77_c17 ;
  wire \u2_Display/lt77_c19 ;
  wire \u2_Display/lt77_c21 ;
  wire \u2_Display/lt77_c23 ;
  wire \u2_Display/lt77_c25 ;
  wire \u2_Display/lt77_c27 ;
  wire \u2_Display/lt77_c29 ;
  wire \u2_Display/lt77_c3 ;
  wire \u2_Display/lt77_c31 ;
  wire \u2_Display/lt77_c5 ;
  wire \u2_Display/lt77_c7 ;
  wire \u2_Display/lt77_c9 ;
  wire \u2_Display/lt7_2_c1 ;
  wire \u2_Display/lt7_2_c11 ;
  wire \u2_Display/lt7_2_c13 ;
  wire \u2_Display/lt7_2_c3 ;
  wire \u2_Display/lt7_2_c5 ;
  wire \u2_Display/lt7_2_c7 ;
  wire \u2_Display/lt7_2_c9 ;
  wire \u2_Display/lt88_c1 ;
  wire \u2_Display/lt88_c11 ;
  wire \u2_Display/lt88_c13 ;
  wire \u2_Display/lt88_c15 ;
  wire \u2_Display/lt88_c17 ;
  wire \u2_Display/lt88_c19 ;
  wire \u2_Display/lt88_c21 ;
  wire \u2_Display/lt88_c23 ;
  wire \u2_Display/lt88_c25 ;
  wire \u2_Display/lt88_c27 ;
  wire \u2_Display/lt88_c29 ;
  wire \u2_Display/lt88_c3 ;
  wire \u2_Display/lt88_c31 ;
  wire \u2_Display/lt88_c5 ;
  wire \u2_Display/lt88_c7 ;
  wire \u2_Display/lt88_c9 ;
  wire \u2_Display/lt89_c1 ;
  wire \u2_Display/lt89_c11 ;
  wire \u2_Display/lt89_c13 ;
  wire \u2_Display/lt89_c15 ;
  wire \u2_Display/lt89_c17 ;
  wire \u2_Display/lt89_c19 ;
  wire \u2_Display/lt89_c21 ;
  wire \u2_Display/lt89_c23 ;
  wire \u2_Display/lt89_c25 ;
  wire \u2_Display/lt89_c27 ;
  wire \u2_Display/lt89_c29 ;
  wire \u2_Display/lt89_c3 ;
  wire \u2_Display/lt89_c31 ;
  wire \u2_Display/lt89_c5 ;
  wire \u2_Display/lt89_c7 ;
  wire \u2_Display/lt89_c9 ;
  wire \u2_Display/lt8_2_c1 ;
  wire \u2_Display/lt8_2_c11 ;
  wire \u2_Display/lt8_2_c3 ;
  wire \u2_Display/lt8_2_c5 ;
  wire \u2_Display/lt8_2_c7 ;
  wire \u2_Display/lt8_2_c9 ;
  wire \u2_Display/lt90_c1 ;
  wire \u2_Display/lt90_c11 ;
  wire \u2_Display/lt90_c13 ;
  wire \u2_Display/lt90_c15 ;
  wire \u2_Display/lt90_c17 ;
  wire \u2_Display/lt90_c19 ;
  wire \u2_Display/lt90_c21 ;
  wire \u2_Display/lt90_c23 ;
  wire \u2_Display/lt90_c25 ;
  wire \u2_Display/lt90_c27 ;
  wire \u2_Display/lt90_c29 ;
  wire \u2_Display/lt90_c3 ;
  wire \u2_Display/lt90_c31 ;
  wire \u2_Display/lt90_c5 ;
  wire \u2_Display/lt90_c7 ;
  wire \u2_Display/lt90_c9 ;
  wire \u2_Display/lt91_c1 ;
  wire \u2_Display/lt91_c11 ;
  wire \u2_Display/lt91_c13 ;
  wire \u2_Display/lt91_c15 ;
  wire \u2_Display/lt91_c17 ;
  wire \u2_Display/lt91_c19 ;
  wire \u2_Display/lt91_c21 ;
  wire \u2_Display/lt91_c23 ;
  wire \u2_Display/lt91_c25 ;
  wire \u2_Display/lt91_c27 ;
  wire \u2_Display/lt91_c29 ;
  wire \u2_Display/lt91_c3 ;
  wire \u2_Display/lt91_c31 ;
  wire \u2_Display/lt91_c5 ;
  wire \u2_Display/lt91_c7 ;
  wire \u2_Display/lt91_c9 ;
  wire \u2_Display/lt92_c1 ;
  wire \u2_Display/lt92_c11 ;
  wire \u2_Display/lt92_c13 ;
  wire \u2_Display/lt92_c15 ;
  wire \u2_Display/lt92_c17 ;
  wire \u2_Display/lt92_c19 ;
  wire \u2_Display/lt92_c21 ;
  wire \u2_Display/lt92_c23 ;
  wire \u2_Display/lt92_c25 ;
  wire \u2_Display/lt92_c27 ;
  wire \u2_Display/lt92_c29 ;
  wire \u2_Display/lt92_c3 ;
  wire \u2_Display/lt92_c31 ;
  wire \u2_Display/lt92_c5 ;
  wire \u2_Display/lt92_c7 ;
  wire \u2_Display/lt92_c9 ;
  wire \u2_Display/lt93_c1 ;
  wire \u2_Display/lt93_c11 ;
  wire \u2_Display/lt93_c13 ;
  wire \u2_Display/lt93_c15 ;
  wire \u2_Display/lt93_c17 ;
  wire \u2_Display/lt93_c19 ;
  wire \u2_Display/lt93_c21 ;
  wire \u2_Display/lt93_c23 ;
  wire \u2_Display/lt93_c25 ;
  wire \u2_Display/lt93_c27 ;
  wire \u2_Display/lt93_c29 ;
  wire \u2_Display/lt93_c3 ;
  wire \u2_Display/lt93_c31 ;
  wire \u2_Display/lt93_c5 ;
  wire \u2_Display/lt93_c7 ;
  wire \u2_Display/lt93_c9 ;
  wire \u2_Display/lt94_c1 ;
  wire \u2_Display/lt94_c11 ;
  wire \u2_Display/lt94_c13 ;
  wire \u2_Display/lt94_c15 ;
  wire \u2_Display/lt94_c17 ;
  wire \u2_Display/lt94_c19 ;
  wire \u2_Display/lt94_c21 ;
  wire \u2_Display/lt94_c23 ;
  wire \u2_Display/lt94_c25 ;
  wire \u2_Display/lt94_c27 ;
  wire \u2_Display/lt94_c29 ;
  wire \u2_Display/lt94_c3 ;
  wire \u2_Display/lt94_c31 ;
  wire \u2_Display/lt94_c5 ;
  wire \u2_Display/lt94_c7 ;
  wire \u2_Display/lt94_c9 ;
  wire \u2_Display/lt95_c1 ;
  wire \u2_Display/lt95_c11 ;
  wire \u2_Display/lt95_c13 ;
  wire \u2_Display/lt95_c15 ;
  wire \u2_Display/lt95_c17 ;
  wire \u2_Display/lt95_c19 ;
  wire \u2_Display/lt95_c21 ;
  wire \u2_Display/lt95_c23 ;
  wire \u2_Display/lt95_c25 ;
  wire \u2_Display/lt95_c27 ;
  wire \u2_Display/lt95_c29 ;
  wire \u2_Display/lt95_c3 ;
  wire \u2_Display/lt95_c31 ;
  wire \u2_Display/lt95_c5 ;
  wire \u2_Display/lt95_c7 ;
  wire \u2_Display/lt95_c9 ;
  wire \u2_Display/lt96_c1 ;
  wire \u2_Display/lt96_c11 ;
  wire \u2_Display/lt96_c13 ;
  wire \u2_Display/lt96_c15 ;
  wire \u2_Display/lt96_c17 ;
  wire \u2_Display/lt96_c19 ;
  wire \u2_Display/lt96_c21 ;
  wire \u2_Display/lt96_c23 ;
  wire \u2_Display/lt96_c25 ;
  wire \u2_Display/lt96_c27 ;
  wire \u2_Display/lt96_c29 ;
  wire \u2_Display/lt96_c3 ;
  wire \u2_Display/lt96_c31 ;
  wire \u2_Display/lt96_c5 ;
  wire \u2_Display/lt96_c7 ;
  wire \u2_Display/lt96_c9 ;
  wire \u2_Display/lt97_c1 ;
  wire \u2_Display/lt97_c11 ;
  wire \u2_Display/lt97_c13 ;
  wire \u2_Display/lt97_c15 ;
  wire \u2_Display/lt97_c17 ;
  wire \u2_Display/lt97_c19 ;
  wire \u2_Display/lt97_c21 ;
  wire \u2_Display/lt97_c23 ;
  wire \u2_Display/lt97_c25 ;
  wire \u2_Display/lt97_c27 ;
  wire \u2_Display/lt97_c29 ;
  wire \u2_Display/lt97_c3 ;
  wire \u2_Display/lt97_c31 ;
  wire \u2_Display/lt97_c5 ;
  wire \u2_Display/lt97_c7 ;
  wire \u2_Display/lt97_c9 ;
  wire \u2_Display/lt98_c1 ;
  wire \u2_Display/lt98_c11 ;
  wire \u2_Display/lt98_c13 ;
  wire \u2_Display/lt98_c15 ;
  wire \u2_Display/lt98_c17 ;
  wire \u2_Display/lt98_c19 ;
  wire \u2_Display/lt98_c21 ;
  wire \u2_Display/lt98_c23 ;
  wire \u2_Display/lt98_c25 ;
  wire \u2_Display/lt98_c27 ;
  wire \u2_Display/lt98_c29 ;
  wire \u2_Display/lt98_c3 ;
  wire \u2_Display/lt98_c31 ;
  wire \u2_Display/lt98_c5 ;
  wire \u2_Display/lt98_c7 ;
  wire \u2_Display/lt98_c9 ;
  wire \u2_Display/lt99_c1 ;
  wire \u2_Display/lt99_c11 ;
  wire \u2_Display/lt99_c13 ;
  wire \u2_Display/lt99_c15 ;
  wire \u2_Display/lt99_c17 ;
  wire \u2_Display/lt99_c19 ;
  wire \u2_Display/lt99_c21 ;
  wire \u2_Display/lt99_c23 ;
  wire \u2_Display/lt99_c25 ;
  wire \u2_Display/lt99_c27 ;
  wire \u2_Display/lt99_c29 ;
  wire \u2_Display/lt99_c3 ;
  wire \u2_Display/lt99_c31 ;
  wire \u2_Display/lt99_c5 ;
  wire \u2_Display/lt99_c7 ;
  wire \u2_Display/lt99_c9 ;
  wire \u2_Display/lt9_2_c1 ;
  wire \u2_Display/lt9_2_c11 ;
  wire \u2_Display/lt9_2_c13 ;
  wire \u2_Display/lt9_2_c3 ;
  wire \u2_Display/lt9_2_c5 ;
  wire \u2_Display/lt9_2_c7 ;
  wire \u2_Display/lt9_2_c9 ;
  wire \u2_Display/mux11_b0_sel_is_0_o ;
  wire \u2_Display/mux19_b0_sel_is_0_o ;
  wire \u2_Display/mux21_b0_sel_is_0_o ;
  wire \u2_Display/mux5_b0_sel_is_0_o ;
  wire \u2_Display/n100 ;
  wire \u2_Display/n1000 ;
  wire \u2_Display/n1001 ;
  wire \u2_Display/n1002 ;
  wire \u2_Display/n1003 ;
  wire \u2_Display/n1004 ;
  wire \u2_Display/n1005 ;
  wire \u2_Display/n1006 ;
  wire \u2_Display/n1007 ;
  wire \u2_Display/n1008 ;
  wire \u2_Display/n1009 ;
  wire \u2_Display/n1010 ;
  wire \u2_Display/n1011 ;
  wire \u2_Display/n1012 ;
  wire \u2_Display/n1015 ;
  wire \u2_Display/n1016 ;
  wire \u2_Display/n1017 ;
  wire \u2_Display/n1018 ;
  wire \u2_Display/n1019 ;
  wire \u2_Display/n1020 ;
  wire \u2_Display/n1021 ;
  wire \u2_Display/n1022 ;
  wire \u2_Display/n1023 ;
  wire \u2_Display/n1024 ;
  wire \u2_Display/n1025 ;
  wire \u2_Display/n1026 ;
  wire \u2_Display/n1027 ;
  wire \u2_Display/n1028 ;
  wire \u2_Display/n1029 ;
  wire \u2_Display/n103 ;
  wire \u2_Display/n1030 ;
  wire \u2_Display/n1031 ;
  wire \u2_Display/n1032 ;
  wire \u2_Display/n1033 ;
  wire \u2_Display/n1034 ;
  wire \u2_Display/n1035 ;
  wire \u2_Display/n1036 ;
  wire \u2_Display/n1037 ;
  wire \u2_Display/n1038 ;
  wire \u2_Display/n1039 ;
  wire \u2_Display/n104 ;
  wire \u2_Display/n1040 ;
  wire \u2_Display/n1041 ;
  wire \u2_Display/n1042 ;
  wire \u2_Display/n1043 ;
  wire \u2_Display/n1044 ;
  wire \u2_Display/n1045 ;
  wire \u2_Display/n1046 ;
  wire \u2_Display/n1047 ;
  wire \u2_Display/n1050 ;
  wire \u2_Display/n1051 ;
  wire \u2_Display/n1052 ;
  wire \u2_Display/n1053 ;
  wire \u2_Display/n1054 ;
  wire \u2_Display/n1055 ;
  wire \u2_Display/n1056 ;
  wire \u2_Display/n1057 ;
  wire \u2_Display/n1058 ;
  wire \u2_Display/n1059 ;
  wire \u2_Display/n1060 ;
  wire \u2_Display/n1061 ;
  wire \u2_Display/n1062 ;
  wire \u2_Display/n1063 ;
  wire \u2_Display/n1064 ;
  wire \u2_Display/n1065 ;
  wire \u2_Display/n1066 ;
  wire \u2_Display/n1067 ;
  wire \u2_Display/n1068 ;
  wire \u2_Display/n1069 ;
  wire \u2_Display/n1070 ;
  wire \u2_Display/n1071 ;
  wire \u2_Display/n1072 ;
  wire \u2_Display/n1073 ;
  wire \u2_Display/n1074 ;
  wire \u2_Display/n1075 ;
  wire \u2_Display/n1076 ;
  wire \u2_Display/n1077 ;
  wire \u2_Display/n1078 ;
  wire \u2_Display/n1079 ;
  wire \u2_Display/n1080 ;
  wire \u2_Display/n1081 ;
  wire \u2_Display/n1082 ;
  wire \u2_Display/n1085 ;
  wire \u2_Display/n1086 ;
  wire \u2_Display/n1087 ;
  wire \u2_Display/n1088 ;
  wire \u2_Display/n1089 ;
  wire \u2_Display/n1090 ;
  wire \u2_Display/n1091 ;
  wire \u2_Display/n1092 ;
  wire \u2_Display/n1093 ;
  wire \u2_Display/n1094 ;
  wire \u2_Display/n1095 ;
  wire \u2_Display/n1096 ;
  wire \u2_Display/n1097 ;
  wire \u2_Display/n1098 ;
  wire \u2_Display/n1099 ;
  wire \u2_Display/n1100 ;
  wire \u2_Display/n1101 ;
  wire \u2_Display/n1102 ;
  wire \u2_Display/n1103 ;
  wire \u2_Display/n1104 ;
  wire \u2_Display/n1105 ;
  wire \u2_Display/n1106 ;
  wire \u2_Display/n1107 ;
  wire \u2_Display/n1108 ;
  wire \u2_Display/n1109 ;
  wire \u2_Display/n1110 ;
  wire \u2_Display/n1111 ;
  wire \u2_Display/n1112 ;
  wire \u2_Display/n1113 ;
  wire \u2_Display/n1114 ;
  wire \u2_Display/n1115 ;
  wire \u2_Display/n1116 ;
  wire \u2_Display/n1117 ;
  wire \u2_Display/n1120 ;
  wire \u2_Display/n1121 ;
  wire \u2_Display/n1122 ;
  wire \u2_Display/n1123 ;
  wire \u2_Display/n1124 ;
  wire \u2_Display/n1125 ;
  wire \u2_Display/n1126 ;
  wire \u2_Display/n1127 ;
  wire \u2_Display/n1128 ;
  wire \u2_Display/n1129 ;
  wire \u2_Display/n1130 ;
  wire \u2_Display/n1131 ;
  wire \u2_Display/n1132 ;
  wire \u2_Display/n1133 ;
  wire \u2_Display/n1134 ;
  wire \u2_Display/n1135 ;
  wire \u2_Display/n1136 ;
  wire \u2_Display/n1137 ;
  wire \u2_Display/n1138 ;
  wire \u2_Display/n1139 ;
  wire \u2_Display/n1140 ;
  wire \u2_Display/n1141 ;
  wire \u2_Display/n1142 ;
  wire \u2_Display/n1143 ;
  wire \u2_Display/n1144 ;
  wire \u2_Display/n1145 ;
  wire \u2_Display/n1146 ;
  wire \u2_Display/n1147 ;
  wire \u2_Display/n1148 ;
  wire \u2_Display/n1149 ;
  wire \u2_Display/n1150 ;
  wire \u2_Display/n1151 ;
  wire \u2_Display/n1152 ;
  wire \u2_Display/n1155 ;
  wire \u2_Display/n1156 ;
  wire \u2_Display/n1157 ;
  wire \u2_Display/n1158 ;
  wire \u2_Display/n1159 ;
  wire \u2_Display/n1160 ;
  wire \u2_Display/n1161 ;
  wire \u2_Display/n1162 ;
  wire \u2_Display/n1163 ;
  wire \u2_Display/n1164 ;
  wire \u2_Display/n1165 ;
  wire \u2_Display/n1166 ;
  wire \u2_Display/n1167 ;
  wire \u2_Display/n1168 ;
  wire \u2_Display/n1169 ;
  wire \u2_Display/n1170 ;
  wire \u2_Display/n1171 ;
  wire \u2_Display/n1172 ;
  wire \u2_Display/n1173 ;
  wire \u2_Display/n1174 ;
  wire \u2_Display/n1175 ;
  wire \u2_Display/n1176 ;
  wire \u2_Display/n1177 ;
  wire \u2_Display/n1178 ;
  wire \u2_Display/n1179 ;
  wire \u2_Display/n1180 ;
  wire \u2_Display/n1181 ;
  wire \u2_Display/n1182 ;
  wire \u2_Display/n1183 ;
  wire \u2_Display/n1184 ;
  wire \u2_Display/n1185 ;
  wire \u2_Display/n1186 ;
  wire \u2_Display/n1187 ;
  wire \u2_Display/n136 ;
  wire \u2_Display/n138 ;
  wire \u2_Display/n141 ;
  wire \u2_Display/n144 ;
  wire \u2_Display/n145 ;
  wire \u2_Display/n1540 ;
  wire \u2_Display/n1543 ;
  wire \u2_Display/n1544 ;
  wire \u2_Display/n1545 ;
  wire \u2_Display/n1546 ;
  wire \u2_Display/n1547 ;
  wire \u2_Display/n1548 ;
  wire \u2_Display/n1549 ;
  wire \u2_Display/n1550 ;
  wire \u2_Display/n1551 ;
  wire \u2_Display/n1552 ;
  wire \u2_Display/n1553 ;
  wire \u2_Display/n1554 ;
  wire \u2_Display/n1555 ;
  wire \u2_Display/n1556 ;
  wire \u2_Display/n1557 ;
  wire \u2_Display/n1558 ;
  wire \u2_Display/n1559 ;
  wire \u2_Display/n1560 ;
  wire \u2_Display/n1561 ;
  wire \u2_Display/n1562 ;
  wire \u2_Display/n1563 ;
  wire \u2_Display/n1564 ;
  wire \u2_Display/n1565 ;
  wire \u2_Display/n1566 ;
  wire \u2_Display/n1567 ;
  wire \u2_Display/n1568 ;
  wire \u2_Display/n1569 ;
  wire \u2_Display/n1570 ;
  wire \u2_Display/n1571 ;
  wire \u2_Display/n1572 ;
  wire \u2_Display/n1573 ;
  wire \u2_Display/n1574 ;
  wire \u2_Display/n1575 ;
  wire \u2_Display/n1578 ;
  wire \u2_Display/n1579 ;
  wire \u2_Display/n1580 ;
  wire \u2_Display/n1581 ;
  wire \u2_Display/n1582 ;
  wire \u2_Display/n1583 ;
  wire \u2_Display/n1584 ;
  wire \u2_Display/n1585 ;
  wire \u2_Display/n1586 ;
  wire \u2_Display/n1587 ;
  wire \u2_Display/n1588 ;
  wire \u2_Display/n1589 ;
  wire \u2_Display/n1590 ;
  wire \u2_Display/n1591 ;
  wire \u2_Display/n1592 ;
  wire \u2_Display/n1593 ;
  wire \u2_Display/n1594 ;
  wire \u2_Display/n1595 ;
  wire \u2_Display/n1596 ;
  wire \u2_Display/n1597 ;
  wire \u2_Display/n1598 ;
  wire \u2_Display/n1599 ;
  wire \u2_Display/n1600 ;
  wire \u2_Display/n1601 ;
  wire \u2_Display/n1602 ;
  wire \u2_Display/n1603 ;
  wire \u2_Display/n1604 ;
  wire \u2_Display/n1605 ;
  wire \u2_Display/n1606 ;
  wire \u2_Display/n1607 ;
  wire \u2_Display/n1608 ;
  wire \u2_Display/n1609 ;
  wire \u2_Display/n1610 ;
  wire \u2_Display/n1613 ;
  wire \u2_Display/n1614 ;
  wire \u2_Display/n1615 ;
  wire \u2_Display/n1616 ;
  wire \u2_Display/n1617 ;
  wire \u2_Display/n1618 ;
  wire \u2_Display/n1619 ;
  wire \u2_Display/n1620 ;
  wire \u2_Display/n1621 ;
  wire \u2_Display/n1622 ;
  wire \u2_Display/n1623 ;
  wire \u2_Display/n1624 ;
  wire \u2_Display/n1625 ;
  wire \u2_Display/n1626 ;
  wire \u2_Display/n1627 ;
  wire \u2_Display/n1628 ;
  wire \u2_Display/n1629 ;
  wire \u2_Display/n1630 ;
  wire \u2_Display/n1631 ;
  wire \u2_Display/n1632 ;
  wire \u2_Display/n1633 ;
  wire \u2_Display/n1634 ;
  wire \u2_Display/n1635 ;
  wire \u2_Display/n1636 ;
  wire \u2_Display/n1637 ;
  wire \u2_Display/n1638 ;
  wire \u2_Display/n1639 ;
  wire \u2_Display/n1640 ;
  wire \u2_Display/n1641 ;
  wire \u2_Display/n1642 ;
  wire \u2_Display/n1643 ;
  wire \u2_Display/n1644 ;
  wire \u2_Display/n1645 ;
  wire \u2_Display/n1648 ;
  wire \u2_Display/n1649 ;
  wire \u2_Display/n1650 ;
  wire \u2_Display/n1651 ;
  wire \u2_Display/n1652 ;
  wire \u2_Display/n1653 ;
  wire \u2_Display/n1654 ;
  wire \u2_Display/n1655 ;
  wire \u2_Display/n1656 ;
  wire \u2_Display/n1657 ;
  wire \u2_Display/n1658 ;
  wire \u2_Display/n1659 ;
  wire \u2_Display/n1660 ;
  wire \u2_Display/n1661 ;
  wire \u2_Display/n1662 ;
  wire \u2_Display/n1663 ;
  wire \u2_Display/n1664 ;
  wire \u2_Display/n1665 ;
  wire \u2_Display/n1666 ;
  wire \u2_Display/n1667 ;
  wire \u2_Display/n1668 ;
  wire \u2_Display/n1669 ;
  wire \u2_Display/n1670 ;
  wire \u2_Display/n1671 ;
  wire \u2_Display/n1672 ;
  wire \u2_Display/n1673 ;
  wire \u2_Display/n1674 ;
  wire \u2_Display/n1675 ;
  wire \u2_Display/n1676 ;
  wire \u2_Display/n1677 ;
  wire \u2_Display/n1678 ;
  wire \u2_Display/n1679 ;
  wire \u2_Display/n1680 ;
  wire \u2_Display/n1683 ;
  wire \u2_Display/n1684 ;
  wire \u2_Display/n1685 ;
  wire \u2_Display/n1686 ;
  wire \u2_Display/n1687 ;
  wire \u2_Display/n1688 ;
  wire \u2_Display/n1689 ;
  wire \u2_Display/n1690 ;
  wire \u2_Display/n1691 ;
  wire \u2_Display/n1692 ;
  wire \u2_Display/n1693 ;
  wire \u2_Display/n1694 ;
  wire \u2_Display/n1695 ;
  wire \u2_Display/n1696 ;
  wire \u2_Display/n1697 ;
  wire \u2_Display/n1698 ;
  wire \u2_Display/n1699 ;
  wire \u2_Display/n1700 ;
  wire \u2_Display/n1701 ;
  wire \u2_Display/n1702 ;
  wire \u2_Display/n1703 ;
  wire \u2_Display/n1704 ;
  wire \u2_Display/n1705 ;
  wire \u2_Display/n1706 ;
  wire \u2_Display/n1707 ;
  wire \u2_Display/n1708 ;
  wire \u2_Display/n1709 ;
  wire \u2_Display/n1710 ;
  wire \u2_Display/n1711 ;
  wire \u2_Display/n1712 ;
  wire \u2_Display/n1713 ;
  wire \u2_Display/n1714 ;
  wire \u2_Display/n1715 ;
  wire \u2_Display/n1718 ;
  wire \u2_Display/n1719 ;
  wire \u2_Display/n1720 ;
  wire \u2_Display/n1721 ;
  wire \u2_Display/n1722 ;
  wire \u2_Display/n1723 ;
  wire \u2_Display/n1724 ;
  wire \u2_Display/n1725 ;
  wire \u2_Display/n1726 ;
  wire \u2_Display/n1727 ;
  wire \u2_Display/n1728 ;
  wire \u2_Display/n1729 ;
  wire \u2_Display/n1730 ;
  wire \u2_Display/n1731 ;
  wire \u2_Display/n1732 ;
  wire \u2_Display/n1733 ;
  wire \u2_Display/n1734 ;
  wire \u2_Display/n1735 ;
  wire \u2_Display/n1736 ;
  wire \u2_Display/n1737 ;
  wire \u2_Display/n1738 ;
  wire \u2_Display/n1739 ;
  wire \u2_Display/n1740 ;
  wire \u2_Display/n1741 ;
  wire \u2_Display/n1742 ;
  wire \u2_Display/n1743 ;
  wire \u2_Display/n1744 ;
  wire \u2_Display/n1745 ;
  wire \u2_Display/n1746 ;
  wire \u2_Display/n1747 ;
  wire \u2_Display/n1748 ;
  wire \u2_Display/n1749 ;
  wire \u2_Display/n1750 ;
  wire \u2_Display/n1753 ;
  wire \u2_Display/n1754 ;
  wire \u2_Display/n1755 ;
  wire \u2_Display/n1756 ;
  wire \u2_Display/n1757 ;
  wire \u2_Display/n1758 ;
  wire \u2_Display/n1759 ;
  wire \u2_Display/n1760 ;
  wire \u2_Display/n1761 ;
  wire \u2_Display/n1762 ;
  wire \u2_Display/n1763 ;
  wire \u2_Display/n1764 ;
  wire \u2_Display/n1765 ;
  wire \u2_Display/n1766 ;
  wire \u2_Display/n1767 ;
  wire \u2_Display/n1768 ;
  wire \u2_Display/n1769 ;
  wire \u2_Display/n1770 ;
  wire \u2_Display/n1771 ;
  wire \u2_Display/n1772 ;
  wire \u2_Display/n1773 ;
  wire \u2_Display/n1774 ;
  wire \u2_Display/n1775 ;
  wire \u2_Display/n1776 ;
  wire \u2_Display/n1777 ;
  wire \u2_Display/n1778 ;
  wire \u2_Display/n1779 ;
  wire \u2_Display/n1780 ;
  wire \u2_Display/n1781 ;
  wire \u2_Display/n1782 ;
  wire \u2_Display/n1783 ;
  wire \u2_Display/n1784 ;
  wire \u2_Display/n1785 ;
  wire \u2_Display/n1788 ;
  wire \u2_Display/n1789 ;
  wire \u2_Display/n1790 ;
  wire \u2_Display/n1791 ;
  wire \u2_Display/n1792 ;
  wire \u2_Display/n1793 ;
  wire \u2_Display/n1794 ;
  wire \u2_Display/n1795 ;
  wire \u2_Display/n1796 ;
  wire \u2_Display/n1797 ;
  wire \u2_Display/n1798 ;
  wire \u2_Display/n1799 ;
  wire \u2_Display/n1800 ;
  wire \u2_Display/n1801 ;
  wire \u2_Display/n1802 ;
  wire \u2_Display/n1803 ;
  wire \u2_Display/n1804 ;
  wire \u2_Display/n1805 ;
  wire \u2_Display/n1806 ;
  wire \u2_Display/n1807 ;
  wire \u2_Display/n1808 ;
  wire \u2_Display/n1809 ;
  wire \u2_Display/n1810 ;
  wire \u2_Display/n1811 ;
  wire \u2_Display/n1812 ;
  wire \u2_Display/n1813 ;
  wire \u2_Display/n1814 ;
  wire \u2_Display/n1815 ;
  wire \u2_Display/n1816 ;
  wire \u2_Display/n1817 ;
  wire \u2_Display/n1818 ;
  wire \u2_Display/n1819 ;
  wire \u2_Display/n1820 ;
  wire \u2_Display/n1823 ;
  wire \u2_Display/n1824 ;
  wire \u2_Display/n1825 ;
  wire \u2_Display/n1826 ;
  wire \u2_Display/n1827 ;
  wire \u2_Display/n1828 ;
  wire \u2_Display/n1829 ;
  wire \u2_Display/n1830 ;
  wire \u2_Display/n1831 ;
  wire \u2_Display/n1832 ;
  wire \u2_Display/n1833 ;
  wire \u2_Display/n1834 ;
  wire \u2_Display/n1835 ;
  wire \u2_Display/n1836 ;
  wire \u2_Display/n1837 ;
  wire \u2_Display/n1838 ;
  wire \u2_Display/n1839 ;
  wire \u2_Display/n1840 ;
  wire \u2_Display/n1841 ;
  wire \u2_Display/n1842 ;
  wire \u2_Display/n1843 ;
  wire \u2_Display/n1844 ;
  wire \u2_Display/n1845 ;
  wire \u2_Display/n1846 ;
  wire \u2_Display/n1847 ;
  wire \u2_Display/n1848 ;
  wire \u2_Display/n1849 ;
  wire \u2_Display/n1850 ;
  wire \u2_Display/n1851 ;
  wire \u2_Display/n1852 ;
  wire \u2_Display/n1853 ;
  wire \u2_Display/n1854 ;
  wire \u2_Display/n1855 ;
  wire \u2_Display/n1858 ;
  wire \u2_Display/n1859 ;
  wire \u2_Display/n1860 ;
  wire \u2_Display/n1861 ;
  wire \u2_Display/n1862 ;
  wire \u2_Display/n1863 ;
  wire \u2_Display/n1864 ;
  wire \u2_Display/n1865 ;
  wire \u2_Display/n1866 ;
  wire \u2_Display/n1867 ;
  wire \u2_Display/n1868 ;
  wire \u2_Display/n1869 ;
  wire \u2_Display/n1870 ;
  wire \u2_Display/n1871 ;
  wire \u2_Display/n1872 ;
  wire \u2_Display/n1873 ;
  wire \u2_Display/n1874 ;
  wire \u2_Display/n1875 ;
  wire \u2_Display/n1876 ;
  wire \u2_Display/n1877 ;
  wire \u2_Display/n1878 ;
  wire \u2_Display/n1879 ;
  wire \u2_Display/n1880 ;
  wire \u2_Display/n1881 ;
  wire \u2_Display/n1882 ;
  wire \u2_Display/n1883 ;
  wire \u2_Display/n1884 ;
  wire \u2_Display/n1885 ;
  wire \u2_Display/n1886 ;
  wire \u2_Display/n1887 ;
  wire \u2_Display/n1888 ;
  wire \u2_Display/n1889 ;
  wire \u2_Display/n1890 ;
  wire \u2_Display/n1893 ;
  wire \u2_Display/n1894 ;
  wire \u2_Display/n1895 ;
  wire \u2_Display/n1896 ;
  wire \u2_Display/n1897 ;
  wire \u2_Display/n1898 ;
  wire \u2_Display/n1899 ;
  wire \u2_Display/n1900 ;
  wire \u2_Display/n1901 ;
  wire \u2_Display/n1902 ;
  wire \u2_Display/n1903 ;
  wire \u2_Display/n1904 ;
  wire \u2_Display/n1905 ;
  wire \u2_Display/n1906 ;
  wire \u2_Display/n1907 ;
  wire \u2_Display/n1908 ;
  wire \u2_Display/n1909 ;
  wire \u2_Display/n1910 ;
  wire \u2_Display/n1911 ;
  wire \u2_Display/n1912 ;
  wire \u2_Display/n1913 ;
  wire \u2_Display/n1914 ;
  wire \u2_Display/n1915 ;
  wire \u2_Display/n1916 ;
  wire \u2_Display/n1917 ;
  wire \u2_Display/n1918 ;
  wire \u2_Display/n1919 ;
  wire \u2_Display/n1920 ;
  wire \u2_Display/n1921 ;
  wire \u2_Display/n1922 ;
  wire \u2_Display/n1923 ;
  wire \u2_Display/n1924 ;
  wire \u2_Display/n1925 ;
  wire \u2_Display/n1928 ;
  wire \u2_Display/n1929 ;
  wire \u2_Display/n1930 ;
  wire \u2_Display/n1931 ;
  wire \u2_Display/n1932 ;
  wire \u2_Display/n1933 ;
  wire \u2_Display/n1934 ;
  wire \u2_Display/n1935 ;
  wire \u2_Display/n1936 ;
  wire \u2_Display/n1937 ;
  wire \u2_Display/n1938 ;
  wire \u2_Display/n1939 ;
  wire \u2_Display/n1940 ;
  wire \u2_Display/n1941 ;
  wire \u2_Display/n1942 ;
  wire \u2_Display/n1943 ;
  wire \u2_Display/n1944 ;
  wire \u2_Display/n1945 ;
  wire \u2_Display/n1946 ;
  wire \u2_Display/n1947 ;
  wire \u2_Display/n1948 ;
  wire \u2_Display/n1949 ;
  wire \u2_Display/n1950 ;
  wire \u2_Display/n1951 ;
  wire \u2_Display/n1952 ;
  wire \u2_Display/n1953 ;
  wire \u2_Display/n1954 ;
  wire \u2_Display/n1955 ;
  wire \u2_Display/n1956 ;
  wire \u2_Display/n1957 ;
  wire \u2_Display/n1958 ;
  wire \u2_Display/n1959 ;
  wire \u2_Display/n1960 ;
  wire \u2_Display/n1963 ;
  wire \u2_Display/n1964 ;
  wire \u2_Display/n1965 ;
  wire \u2_Display/n1966 ;
  wire \u2_Display/n1967 ;
  wire \u2_Display/n1968 ;
  wire \u2_Display/n1969 ;
  wire \u2_Display/n1970 ;
  wire \u2_Display/n1971 ;
  wire \u2_Display/n1972 ;
  wire \u2_Display/n1973 ;
  wire \u2_Display/n1974 ;
  wire \u2_Display/n1975 ;
  wire \u2_Display/n1976 ;
  wire \u2_Display/n1977 ;
  wire \u2_Display/n1978 ;
  wire \u2_Display/n1979 ;
  wire \u2_Display/n1980 ;
  wire \u2_Display/n1981 ;
  wire \u2_Display/n1982 ;
  wire \u2_Display/n1983 ;
  wire \u2_Display/n1984 ;
  wire \u2_Display/n1985 ;
  wire \u2_Display/n1986 ;
  wire \u2_Display/n1987 ;
  wire \u2_Display/n1988 ;
  wire \u2_Display/n1989 ;
  wire \u2_Display/n1990 ;
  wire \u2_Display/n1991 ;
  wire \u2_Display/n1992 ;
  wire \u2_Display/n1993 ;
  wire \u2_Display/n1994 ;
  wire \u2_Display/n1995 ;
  wire \u2_Display/n1998 ;
  wire \u2_Display/n1999 ;
  wire \u2_Display/n2000 ;
  wire \u2_Display/n2001 ;
  wire \u2_Display/n2002 ;
  wire \u2_Display/n2003 ;
  wire \u2_Display/n2004 ;
  wire \u2_Display/n2005 ;
  wire \u2_Display/n2006 ;
  wire \u2_Display/n2007 ;
  wire \u2_Display/n2008 ;
  wire \u2_Display/n2009 ;
  wire \u2_Display/n2010 ;
  wire \u2_Display/n2011 ;
  wire \u2_Display/n2012 ;
  wire \u2_Display/n2013 ;
  wire \u2_Display/n2014 ;
  wire \u2_Display/n2015 ;
  wire \u2_Display/n2016 ;
  wire \u2_Display/n2017 ;
  wire \u2_Display/n2018 ;
  wire \u2_Display/n2019 ;
  wire \u2_Display/n2020 ;
  wire \u2_Display/n2021 ;
  wire \u2_Display/n2022 ;
  wire \u2_Display/n2023 ;
  wire \u2_Display/n2024 ;
  wire \u2_Display/n2025 ;
  wire \u2_Display/n2026 ;
  wire \u2_Display/n2027 ;
  wire \u2_Display/n2028 ;
  wire \u2_Display/n2029 ;
  wire \u2_Display/n2030 ;
  wire \u2_Display/n2033 ;
  wire \u2_Display/n2034 ;
  wire \u2_Display/n2035 ;
  wire \u2_Display/n2036 ;
  wire \u2_Display/n2037 ;
  wire \u2_Display/n2038 ;
  wire \u2_Display/n2039 ;
  wire \u2_Display/n2040 ;
  wire \u2_Display/n2041 ;
  wire \u2_Display/n2042 ;
  wire \u2_Display/n2043 ;
  wire \u2_Display/n2044 ;
  wire \u2_Display/n2045 ;
  wire \u2_Display/n2046 ;
  wire \u2_Display/n2047 ;
  wire \u2_Display/n2048 ;
  wire \u2_Display/n2049 ;
  wire \u2_Display/n2050 ;
  wire \u2_Display/n2051 ;
  wire \u2_Display/n2052 ;
  wire \u2_Display/n2053 ;
  wire \u2_Display/n2054 ;
  wire \u2_Display/n2055 ;
  wire \u2_Display/n2056 ;
  wire \u2_Display/n2057 ;
  wire \u2_Display/n2058 ;
  wire \u2_Display/n2059 ;
  wire \u2_Display/n2060 ;
  wire \u2_Display/n2061 ;
  wire \u2_Display/n2062 ;
  wire \u2_Display/n2063 ;
  wire \u2_Display/n2064 ;
  wire \u2_Display/n2065 ;
  wire \u2_Display/n2068 ;
  wire \u2_Display/n2069 ;
  wire \u2_Display/n2070 ;
  wire \u2_Display/n2071 ;
  wire \u2_Display/n2072 ;
  wire \u2_Display/n2073 ;
  wire \u2_Display/n2074 ;
  wire \u2_Display/n2075 ;
  wire \u2_Display/n2076 ;
  wire \u2_Display/n2077 ;
  wire \u2_Display/n2078 ;
  wire \u2_Display/n2079 ;
  wire \u2_Display/n2080 ;
  wire \u2_Display/n2081 ;
  wire \u2_Display/n2082 ;
  wire \u2_Display/n2083 ;
  wire \u2_Display/n2084 ;
  wire \u2_Display/n2085 ;
  wire \u2_Display/n2086 ;
  wire \u2_Display/n2087 ;
  wire \u2_Display/n2088 ;
  wire \u2_Display/n2089 ;
  wire \u2_Display/n2090 ;
  wire \u2_Display/n2091 ;
  wire \u2_Display/n2092 ;
  wire \u2_Display/n2093 ;
  wire \u2_Display/n2094 ;
  wire \u2_Display/n2095 ;
  wire \u2_Display/n2096 ;
  wire \u2_Display/n2097 ;
  wire \u2_Display/n2098 ;
  wire \u2_Display/n2099 ;
  wire \u2_Display/n2100 ;
  wire \u2_Display/n2103 ;
  wire \u2_Display/n2104 ;
  wire \u2_Display/n2105 ;
  wire \u2_Display/n2106 ;
  wire \u2_Display/n2107 ;
  wire \u2_Display/n2108 ;
  wire \u2_Display/n2109 ;
  wire \u2_Display/n2110 ;
  wire \u2_Display/n2111 ;
  wire \u2_Display/n2112 ;
  wire \u2_Display/n2113 ;
  wire \u2_Display/n2114 ;
  wire \u2_Display/n2115 ;
  wire \u2_Display/n2116 ;
  wire \u2_Display/n2117 ;
  wire \u2_Display/n2118 ;
  wire \u2_Display/n2119 ;
  wire \u2_Display/n2120 ;
  wire \u2_Display/n2121 ;
  wire \u2_Display/n2122 ;
  wire \u2_Display/n2123 ;
  wire \u2_Display/n2124 ;
  wire \u2_Display/n2125 ;
  wire \u2_Display/n2126 ;
  wire \u2_Display/n2127 ;
  wire \u2_Display/n2128 ;
  wire \u2_Display/n2129 ;
  wire \u2_Display/n2130 ;
  wire \u2_Display/n2131 ;
  wire \u2_Display/n2132 ;
  wire \u2_Display/n2133 ;
  wire \u2_Display/n2134 ;
  wire \u2_Display/n2135 ;
  wire \u2_Display/n2138 ;
  wire \u2_Display/n2139 ;
  wire \u2_Display/n2140 ;
  wire \u2_Display/n2141 ;
  wire \u2_Display/n2142 ;
  wire \u2_Display/n2143 ;
  wire \u2_Display/n2144 ;
  wire \u2_Display/n2145 ;
  wire \u2_Display/n2146 ;
  wire \u2_Display/n2147 ;
  wire \u2_Display/n2148 ;
  wire \u2_Display/n2149 ;
  wire \u2_Display/n2150 ;
  wire \u2_Display/n2151 ;
  wire \u2_Display/n2152 ;
  wire \u2_Display/n2153 ;
  wire \u2_Display/n2154 ;
  wire \u2_Display/n2155 ;
  wire \u2_Display/n2156 ;
  wire \u2_Display/n2157 ;
  wire \u2_Display/n2158 ;
  wire \u2_Display/n2159 ;
  wire \u2_Display/n2160 ;
  wire \u2_Display/n2161 ;
  wire \u2_Display/n2162 ;
  wire \u2_Display/n2163 ;
  wire \u2_Display/n2164 ;
  wire \u2_Display/n2165 ;
  wire \u2_Display/n2166 ;
  wire \u2_Display/n2167 ;
  wire \u2_Display/n2168 ;
  wire \u2_Display/n2169 ;
  wire \u2_Display/n2170 ;
  wire \u2_Display/n2173 ;
  wire \u2_Display/n2174 ;
  wire \u2_Display/n2175 ;
  wire \u2_Display/n2176 ;
  wire \u2_Display/n2177 ;
  wire \u2_Display/n2178 ;
  wire \u2_Display/n2179 ;
  wire \u2_Display/n2180 ;
  wire \u2_Display/n2181 ;
  wire \u2_Display/n2182 ;
  wire \u2_Display/n2183 ;
  wire \u2_Display/n2184 ;
  wire \u2_Display/n2185 ;
  wire \u2_Display/n2186 ;
  wire \u2_Display/n2187 ;
  wire \u2_Display/n2188 ;
  wire \u2_Display/n2189 ;
  wire \u2_Display/n2190 ;
  wire \u2_Display/n2191 ;
  wire \u2_Display/n2192 ;
  wire \u2_Display/n2193 ;
  wire \u2_Display/n2194 ;
  wire \u2_Display/n2195 ;
  wire \u2_Display/n2196 ;
  wire \u2_Display/n2197 ;
  wire \u2_Display/n2198 ;
  wire \u2_Display/n2199 ;
  wire \u2_Display/n2200 ;
  wire \u2_Display/n2201 ;
  wire \u2_Display/n2202 ;
  wire \u2_Display/n2203 ;
  wire \u2_Display/n2204 ;
  wire \u2_Display/n2205 ;
  wire \u2_Display/n2208 ;
  wire \u2_Display/n2209 ;
  wire \u2_Display/n2210 ;
  wire \u2_Display/n2211 ;
  wire \u2_Display/n2212 ;
  wire \u2_Display/n2213 ;
  wire \u2_Display/n2214 ;
  wire \u2_Display/n2215 ;
  wire \u2_Display/n2216 ;
  wire \u2_Display/n2217 ;
  wire \u2_Display/n2218 ;
  wire \u2_Display/n2219 ;
  wire \u2_Display/n2220 ;
  wire \u2_Display/n2221 ;
  wire \u2_Display/n2222 ;
  wire \u2_Display/n2223 ;
  wire \u2_Display/n2224 ;
  wire \u2_Display/n2225 ;
  wire \u2_Display/n2226 ;
  wire \u2_Display/n2227 ;
  wire \u2_Display/n2228 ;
  wire \u2_Display/n2229 ;
  wire \u2_Display/n2230 ;
  wire \u2_Display/n2231 ;
  wire \u2_Display/n2232 ;
  wire \u2_Display/n2233 ;
  wire \u2_Display/n2234 ;
  wire \u2_Display/n2235 ;
  wire \u2_Display/n2236 ;
  wire \u2_Display/n2237 ;
  wire \u2_Display/n2238 ;
  wire \u2_Display/n2239 ;
  wire \u2_Display/n2240 ;
  wire \u2_Display/n2243 ;
  wire \u2_Display/n2244 ;
  wire \u2_Display/n2245 ;
  wire \u2_Display/n2246 ;
  wire \u2_Display/n2247 ;
  wire \u2_Display/n2248 ;
  wire \u2_Display/n2249 ;
  wire \u2_Display/n2250 ;
  wire \u2_Display/n2251 ;
  wire \u2_Display/n2252 ;
  wire \u2_Display/n2253 ;
  wire \u2_Display/n2254 ;
  wire \u2_Display/n2255 ;
  wire \u2_Display/n2256 ;
  wire \u2_Display/n2257 ;
  wire \u2_Display/n2258 ;
  wire \u2_Display/n2259 ;
  wire \u2_Display/n2260 ;
  wire \u2_Display/n2261 ;
  wire \u2_Display/n2262 ;
  wire \u2_Display/n2263 ;
  wire \u2_Display/n2264 ;
  wire \u2_Display/n2265 ;
  wire \u2_Display/n2266 ;
  wire \u2_Display/n2267 ;
  wire \u2_Display/n2268 ;
  wire \u2_Display/n2269 ;
  wire \u2_Display/n2270 ;
  wire \u2_Display/n2271 ;
  wire \u2_Display/n2272 ;
  wire \u2_Display/n2273 ;
  wire \u2_Display/n2274 ;
  wire \u2_Display/n2275 ;
  wire \u2_Display/n2278 ;
  wire \u2_Display/n2279 ;
  wire \u2_Display/n2280 ;
  wire \u2_Display/n2281 ;
  wire \u2_Display/n2282 ;
  wire \u2_Display/n2283 ;
  wire \u2_Display/n2284 ;
  wire \u2_Display/n2285 ;
  wire \u2_Display/n2286 ;
  wire \u2_Display/n2287 ;
  wire \u2_Display/n2288 ;
  wire \u2_Display/n2289 ;
  wire \u2_Display/n2290 ;
  wire \u2_Display/n2291 ;
  wire \u2_Display/n2292 ;
  wire \u2_Display/n2293 ;
  wire \u2_Display/n2294 ;
  wire \u2_Display/n2295 ;
  wire \u2_Display/n2296 ;
  wire \u2_Display/n2297 ;
  wire \u2_Display/n2298 ;
  wire \u2_Display/n2299 ;
  wire \u2_Display/n2300 ;
  wire \u2_Display/n2301 ;
  wire \u2_Display/n2302 ;
  wire \u2_Display/n2303 ;
  wire \u2_Display/n2304 ;
  wire \u2_Display/n2305 ;
  wire \u2_Display/n2306 ;
  wire \u2_Display/n2307 ;
  wire \u2_Display/n2308 ;
  wire \u2_Display/n2309 ;
  wire \u2_Display/n2310 ;
  wire \u2_Display/n2663 ;
  wire \u2_Display/n2666 ;
  wire \u2_Display/n2667 ;
  wire \u2_Display/n2668 ;
  wire \u2_Display/n2669 ;
  wire \u2_Display/n2670 ;
  wire \u2_Display/n2671 ;
  wire \u2_Display/n2672 ;
  wire \u2_Display/n2673 ;
  wire \u2_Display/n2674 ;
  wire \u2_Display/n2675 ;
  wire \u2_Display/n2676 ;
  wire \u2_Display/n2677 ;
  wire \u2_Display/n2678 ;
  wire \u2_Display/n2679 ;
  wire \u2_Display/n2680 ;
  wire \u2_Display/n2681 ;
  wire \u2_Display/n2682 ;
  wire \u2_Display/n2683 ;
  wire \u2_Display/n2684 ;
  wire \u2_Display/n2685 ;
  wire \u2_Display/n2686 ;
  wire \u2_Display/n2687 ;
  wire \u2_Display/n2688 ;
  wire \u2_Display/n2689 ;
  wire \u2_Display/n2690 ;
  wire \u2_Display/n2691 ;
  wire \u2_Display/n2692 ;
  wire \u2_Display/n2693 ;
  wire \u2_Display/n2694 ;
  wire \u2_Display/n2695 ;
  wire \u2_Display/n2696 ;
  wire \u2_Display/n2697 ;
  wire \u2_Display/n2698 ;
  wire \u2_Display/n2701 ;
  wire \u2_Display/n2702 ;
  wire \u2_Display/n2703 ;
  wire \u2_Display/n2704 ;
  wire \u2_Display/n2705 ;
  wire \u2_Display/n2706 ;
  wire \u2_Display/n2707 ;
  wire \u2_Display/n2708 ;
  wire \u2_Display/n2709 ;
  wire \u2_Display/n2710 ;
  wire \u2_Display/n2711 ;
  wire \u2_Display/n2712 ;
  wire \u2_Display/n2713 ;
  wire \u2_Display/n2714 ;
  wire \u2_Display/n2715 ;
  wire \u2_Display/n2716 ;
  wire \u2_Display/n2717 ;
  wire \u2_Display/n2718 ;
  wire \u2_Display/n2719 ;
  wire \u2_Display/n2720 ;
  wire \u2_Display/n2721 ;
  wire \u2_Display/n2722 ;
  wire \u2_Display/n2723 ;
  wire \u2_Display/n2724 ;
  wire \u2_Display/n2725 ;
  wire \u2_Display/n2726 ;
  wire \u2_Display/n2727 ;
  wire \u2_Display/n2728 ;
  wire \u2_Display/n2729 ;
  wire \u2_Display/n2730 ;
  wire \u2_Display/n2731 ;
  wire \u2_Display/n2732 ;
  wire \u2_Display/n2733 ;
  wire \u2_Display/n2736 ;
  wire \u2_Display/n2737 ;
  wire \u2_Display/n2738 ;
  wire \u2_Display/n2739 ;
  wire \u2_Display/n2740 ;
  wire \u2_Display/n2741 ;
  wire \u2_Display/n2742 ;
  wire \u2_Display/n2743 ;
  wire \u2_Display/n2744 ;
  wire \u2_Display/n2745 ;
  wire \u2_Display/n2746 ;
  wire \u2_Display/n2747 ;
  wire \u2_Display/n2748 ;
  wire \u2_Display/n2749 ;
  wire \u2_Display/n2750 ;
  wire \u2_Display/n2751 ;
  wire \u2_Display/n2752 ;
  wire \u2_Display/n2753 ;
  wire \u2_Display/n2754 ;
  wire \u2_Display/n2755 ;
  wire \u2_Display/n2756 ;
  wire \u2_Display/n2757 ;
  wire \u2_Display/n2758 ;
  wire \u2_Display/n2759 ;
  wire \u2_Display/n2760 ;
  wire \u2_Display/n2761 ;
  wire \u2_Display/n2762 ;
  wire \u2_Display/n2763 ;
  wire \u2_Display/n2764 ;
  wire \u2_Display/n2765 ;
  wire \u2_Display/n2766 ;
  wire \u2_Display/n2767 ;
  wire \u2_Display/n2768 ;
  wire \u2_Display/n2771 ;
  wire \u2_Display/n2772 ;
  wire \u2_Display/n2773 ;
  wire \u2_Display/n2774 ;
  wire \u2_Display/n2775 ;
  wire \u2_Display/n2776 ;
  wire \u2_Display/n2777 ;
  wire \u2_Display/n2778 ;
  wire \u2_Display/n2779 ;
  wire \u2_Display/n2780 ;
  wire \u2_Display/n2781 ;
  wire \u2_Display/n2782 ;
  wire \u2_Display/n2783 ;
  wire \u2_Display/n2784 ;
  wire \u2_Display/n2785 ;
  wire \u2_Display/n2786 ;
  wire \u2_Display/n2787 ;
  wire \u2_Display/n2788 ;
  wire \u2_Display/n2789 ;
  wire \u2_Display/n2790 ;
  wire \u2_Display/n2791 ;
  wire \u2_Display/n2792 ;
  wire \u2_Display/n2793 ;
  wire \u2_Display/n2794 ;
  wire \u2_Display/n2795 ;
  wire \u2_Display/n2796 ;
  wire \u2_Display/n2797 ;
  wire \u2_Display/n2798 ;
  wire \u2_Display/n2799 ;
  wire \u2_Display/n2800 ;
  wire \u2_Display/n2801 ;
  wire \u2_Display/n2802 ;
  wire \u2_Display/n2803 ;
  wire \u2_Display/n2806 ;
  wire \u2_Display/n2807 ;
  wire \u2_Display/n2808 ;
  wire \u2_Display/n2809 ;
  wire \u2_Display/n2810 ;
  wire \u2_Display/n2811 ;
  wire \u2_Display/n2812 ;
  wire \u2_Display/n2813 ;
  wire \u2_Display/n2814 ;
  wire \u2_Display/n2815 ;
  wire \u2_Display/n2816 ;
  wire \u2_Display/n2817 ;
  wire \u2_Display/n2818 ;
  wire \u2_Display/n2819 ;
  wire \u2_Display/n2820 ;
  wire \u2_Display/n2821 ;
  wire \u2_Display/n2822 ;
  wire \u2_Display/n2823 ;
  wire \u2_Display/n2824 ;
  wire \u2_Display/n2825 ;
  wire \u2_Display/n2826 ;
  wire \u2_Display/n2827 ;
  wire \u2_Display/n2828 ;
  wire \u2_Display/n2829 ;
  wire \u2_Display/n2830 ;
  wire \u2_Display/n2831 ;
  wire \u2_Display/n2832 ;
  wire \u2_Display/n2833 ;
  wire \u2_Display/n2834 ;
  wire \u2_Display/n2835 ;
  wire \u2_Display/n2836 ;
  wire \u2_Display/n2837 ;
  wire \u2_Display/n2838 ;
  wire \u2_Display/n2841 ;
  wire \u2_Display/n2842 ;
  wire \u2_Display/n2843 ;
  wire \u2_Display/n2844 ;
  wire \u2_Display/n2845 ;
  wire \u2_Display/n2846 ;
  wire \u2_Display/n2847 ;
  wire \u2_Display/n2848 ;
  wire \u2_Display/n2849 ;
  wire \u2_Display/n2850 ;
  wire \u2_Display/n2851 ;
  wire \u2_Display/n2852 ;
  wire \u2_Display/n2853 ;
  wire \u2_Display/n2854 ;
  wire \u2_Display/n2855 ;
  wire \u2_Display/n2856 ;
  wire \u2_Display/n2857 ;
  wire \u2_Display/n2858 ;
  wire \u2_Display/n2859 ;
  wire \u2_Display/n2860 ;
  wire \u2_Display/n2861 ;
  wire \u2_Display/n2862 ;
  wire \u2_Display/n2863 ;
  wire \u2_Display/n2864 ;
  wire \u2_Display/n2865 ;
  wire \u2_Display/n2866 ;
  wire \u2_Display/n2867 ;
  wire \u2_Display/n2868 ;
  wire \u2_Display/n2869 ;
  wire \u2_Display/n2870 ;
  wire \u2_Display/n2871 ;
  wire \u2_Display/n2872 ;
  wire \u2_Display/n2873 ;
  wire \u2_Display/n2876 ;
  wire \u2_Display/n2877 ;
  wire \u2_Display/n2878 ;
  wire \u2_Display/n2879 ;
  wire \u2_Display/n2880 ;
  wire \u2_Display/n2881 ;
  wire \u2_Display/n2882 ;
  wire \u2_Display/n2883 ;
  wire \u2_Display/n2884 ;
  wire \u2_Display/n2885 ;
  wire \u2_Display/n2886 ;
  wire \u2_Display/n2887 ;
  wire \u2_Display/n2888 ;
  wire \u2_Display/n2889 ;
  wire \u2_Display/n2890 ;
  wire \u2_Display/n2891 ;
  wire \u2_Display/n2892 ;
  wire \u2_Display/n2893 ;
  wire \u2_Display/n2894 ;
  wire \u2_Display/n2895 ;
  wire \u2_Display/n2896 ;
  wire \u2_Display/n2897 ;
  wire \u2_Display/n2898 ;
  wire \u2_Display/n2899 ;
  wire \u2_Display/n2900 ;
  wire \u2_Display/n2901 ;
  wire \u2_Display/n2902 ;
  wire \u2_Display/n2903 ;
  wire \u2_Display/n2904 ;
  wire \u2_Display/n2905 ;
  wire \u2_Display/n2906 ;
  wire \u2_Display/n2907 ;
  wire \u2_Display/n2908 ;
  wire \u2_Display/n2911 ;
  wire \u2_Display/n2912 ;
  wire \u2_Display/n2913 ;
  wire \u2_Display/n2914 ;
  wire \u2_Display/n2915 ;
  wire \u2_Display/n2916 ;
  wire \u2_Display/n2917 ;
  wire \u2_Display/n2918 ;
  wire \u2_Display/n2919 ;
  wire \u2_Display/n2920 ;
  wire \u2_Display/n2921 ;
  wire \u2_Display/n2922 ;
  wire \u2_Display/n2923 ;
  wire \u2_Display/n2924 ;
  wire \u2_Display/n2925 ;
  wire \u2_Display/n2926 ;
  wire \u2_Display/n2927 ;
  wire \u2_Display/n2928 ;
  wire \u2_Display/n2929 ;
  wire \u2_Display/n2930 ;
  wire \u2_Display/n2931 ;
  wire \u2_Display/n2932 ;
  wire \u2_Display/n2933 ;
  wire \u2_Display/n2934 ;
  wire \u2_Display/n2935 ;
  wire \u2_Display/n2936 ;
  wire \u2_Display/n2937 ;
  wire \u2_Display/n2938 ;
  wire \u2_Display/n2939 ;
  wire \u2_Display/n2940 ;
  wire \u2_Display/n2941 ;
  wire \u2_Display/n2942 ;
  wire \u2_Display/n2943 ;
  wire \u2_Display/n2946 ;
  wire \u2_Display/n2947 ;
  wire \u2_Display/n2948 ;
  wire \u2_Display/n2949 ;
  wire \u2_Display/n2950 ;
  wire \u2_Display/n2951 ;
  wire \u2_Display/n2952 ;
  wire \u2_Display/n2953 ;
  wire \u2_Display/n2954 ;
  wire \u2_Display/n2955 ;
  wire \u2_Display/n2956 ;
  wire \u2_Display/n2957 ;
  wire \u2_Display/n2958 ;
  wire \u2_Display/n2959 ;
  wire \u2_Display/n2960 ;
  wire \u2_Display/n2961 ;
  wire \u2_Display/n2962 ;
  wire \u2_Display/n2963 ;
  wire \u2_Display/n2964 ;
  wire \u2_Display/n2965 ;
  wire \u2_Display/n2966 ;
  wire \u2_Display/n2967 ;
  wire \u2_Display/n2968 ;
  wire \u2_Display/n2969 ;
  wire \u2_Display/n2970 ;
  wire \u2_Display/n2971 ;
  wire \u2_Display/n2972 ;
  wire \u2_Display/n2973 ;
  wire \u2_Display/n2974 ;
  wire \u2_Display/n2975 ;
  wire \u2_Display/n2976 ;
  wire \u2_Display/n2977 ;
  wire \u2_Display/n2978 ;
  wire \u2_Display/n2981 ;
  wire \u2_Display/n2982 ;
  wire \u2_Display/n2983 ;
  wire \u2_Display/n2984 ;
  wire \u2_Display/n2985 ;
  wire \u2_Display/n2986 ;
  wire \u2_Display/n2987 ;
  wire \u2_Display/n2988 ;
  wire \u2_Display/n2989 ;
  wire \u2_Display/n2990 ;
  wire \u2_Display/n2991 ;
  wire \u2_Display/n2992 ;
  wire \u2_Display/n2993 ;
  wire \u2_Display/n2994 ;
  wire \u2_Display/n2995 ;
  wire \u2_Display/n2996 ;
  wire \u2_Display/n2997 ;
  wire \u2_Display/n2998 ;
  wire \u2_Display/n2999 ;
  wire \u2_Display/n3000 ;
  wire \u2_Display/n3001 ;
  wire \u2_Display/n3002 ;
  wire \u2_Display/n3003 ;
  wire \u2_Display/n3004 ;
  wire \u2_Display/n3005 ;
  wire \u2_Display/n3006 ;
  wire \u2_Display/n3007 ;
  wire \u2_Display/n3008 ;
  wire \u2_Display/n3009 ;
  wire \u2_Display/n3010 ;
  wire \u2_Display/n3011 ;
  wire \u2_Display/n3012 ;
  wire \u2_Display/n3013 ;
  wire \u2_Display/n3016 ;
  wire \u2_Display/n3017 ;
  wire \u2_Display/n3018 ;
  wire \u2_Display/n3019 ;
  wire \u2_Display/n3020 ;
  wire \u2_Display/n3021 ;
  wire \u2_Display/n3022 ;
  wire \u2_Display/n3023 ;
  wire \u2_Display/n3024 ;
  wire \u2_Display/n3025 ;
  wire \u2_Display/n3026 ;
  wire \u2_Display/n3027 ;
  wire \u2_Display/n3028 ;
  wire \u2_Display/n3029 ;
  wire \u2_Display/n3030 ;
  wire \u2_Display/n3031 ;
  wire \u2_Display/n3032 ;
  wire \u2_Display/n3033 ;
  wire \u2_Display/n3034 ;
  wire \u2_Display/n3035 ;
  wire \u2_Display/n3036 ;
  wire \u2_Display/n3037 ;
  wire \u2_Display/n3038 ;
  wire \u2_Display/n3039 ;
  wire \u2_Display/n3040 ;
  wire \u2_Display/n3041 ;
  wire \u2_Display/n3042 ;
  wire \u2_Display/n3043 ;
  wire \u2_Display/n3044 ;
  wire \u2_Display/n3045 ;
  wire \u2_Display/n3046 ;
  wire \u2_Display/n3047 ;
  wire \u2_Display/n3048 ;
  wire \u2_Display/n3051 ;
  wire \u2_Display/n3052 ;
  wire \u2_Display/n3053 ;
  wire \u2_Display/n3054 ;
  wire \u2_Display/n3055 ;
  wire \u2_Display/n3056 ;
  wire \u2_Display/n3057 ;
  wire \u2_Display/n3058 ;
  wire \u2_Display/n3059 ;
  wire \u2_Display/n3060 ;
  wire \u2_Display/n3061 ;
  wire \u2_Display/n3062 ;
  wire \u2_Display/n3063 ;
  wire \u2_Display/n3064 ;
  wire \u2_Display/n3065 ;
  wire \u2_Display/n3066 ;
  wire \u2_Display/n3067 ;
  wire \u2_Display/n3068 ;
  wire \u2_Display/n3069 ;
  wire \u2_Display/n3070 ;
  wire \u2_Display/n3071 ;
  wire \u2_Display/n3072 ;
  wire \u2_Display/n3073 ;
  wire \u2_Display/n3074 ;
  wire \u2_Display/n3075 ;
  wire \u2_Display/n3076 ;
  wire \u2_Display/n3077 ;
  wire \u2_Display/n3078 ;
  wire \u2_Display/n3079 ;
  wire \u2_Display/n3080 ;
  wire \u2_Display/n3081 ;
  wire \u2_Display/n3082 ;
  wire \u2_Display/n3083 ;
  wire \u2_Display/n3086 ;
  wire \u2_Display/n3087 ;
  wire \u2_Display/n3088 ;
  wire \u2_Display/n3089 ;
  wire \u2_Display/n3090 ;
  wire \u2_Display/n3091 ;
  wire \u2_Display/n3092 ;
  wire \u2_Display/n3093 ;
  wire \u2_Display/n3094 ;
  wire \u2_Display/n3095 ;
  wire \u2_Display/n3096 ;
  wire \u2_Display/n3097 ;
  wire \u2_Display/n3098 ;
  wire \u2_Display/n3099 ;
  wire \u2_Display/n3100 ;
  wire \u2_Display/n3101 ;
  wire \u2_Display/n3102 ;
  wire \u2_Display/n3103 ;
  wire \u2_Display/n3104 ;
  wire \u2_Display/n3105 ;
  wire \u2_Display/n3106 ;
  wire \u2_Display/n3107 ;
  wire \u2_Display/n3108 ;
  wire \u2_Display/n3109 ;
  wire \u2_Display/n3110 ;
  wire \u2_Display/n3111 ;
  wire \u2_Display/n3112 ;
  wire \u2_Display/n3113 ;
  wire \u2_Display/n3114 ;
  wire \u2_Display/n3115 ;
  wire \u2_Display/n3116 ;
  wire \u2_Display/n3117 ;
  wire \u2_Display/n3118 ;
  wire \u2_Display/n3121 ;
  wire \u2_Display/n3122 ;
  wire \u2_Display/n3123 ;
  wire \u2_Display/n3124 ;
  wire \u2_Display/n3125 ;
  wire \u2_Display/n3126 ;
  wire \u2_Display/n3127 ;
  wire \u2_Display/n3128 ;
  wire \u2_Display/n3129 ;
  wire \u2_Display/n3130 ;
  wire \u2_Display/n3131 ;
  wire \u2_Display/n3132 ;
  wire \u2_Display/n3133 ;
  wire \u2_Display/n3134 ;
  wire \u2_Display/n3135 ;
  wire \u2_Display/n3136 ;
  wire \u2_Display/n3137 ;
  wire \u2_Display/n3138 ;
  wire \u2_Display/n3139 ;
  wire \u2_Display/n3140 ;
  wire \u2_Display/n3141 ;
  wire \u2_Display/n3142 ;
  wire \u2_Display/n3143 ;
  wire \u2_Display/n3144 ;
  wire \u2_Display/n3145 ;
  wire \u2_Display/n3146 ;
  wire \u2_Display/n3147 ;
  wire \u2_Display/n3148 ;
  wire \u2_Display/n3149 ;
  wire \u2_Display/n3150 ;
  wire \u2_Display/n3151 ;
  wire \u2_Display/n3152 ;
  wire \u2_Display/n3153 ;
  wire \u2_Display/n3156 ;
  wire \u2_Display/n3157 ;
  wire \u2_Display/n3158 ;
  wire \u2_Display/n3159 ;
  wire \u2_Display/n3160 ;
  wire \u2_Display/n3161 ;
  wire \u2_Display/n3162 ;
  wire \u2_Display/n3163 ;
  wire \u2_Display/n3164 ;
  wire \u2_Display/n3165 ;
  wire \u2_Display/n3166 ;
  wire \u2_Display/n3167 ;
  wire \u2_Display/n3168 ;
  wire \u2_Display/n3169 ;
  wire \u2_Display/n3170 ;
  wire \u2_Display/n3171 ;
  wire \u2_Display/n3172 ;
  wire \u2_Display/n3173 ;
  wire \u2_Display/n3174 ;
  wire \u2_Display/n3175 ;
  wire \u2_Display/n3176 ;
  wire \u2_Display/n3177 ;
  wire \u2_Display/n3178 ;
  wire \u2_Display/n3179 ;
  wire \u2_Display/n3180 ;
  wire \u2_Display/n3181 ;
  wire \u2_Display/n3182 ;
  wire \u2_Display/n3183 ;
  wire \u2_Display/n3184 ;
  wire \u2_Display/n3185 ;
  wire \u2_Display/n3186 ;
  wire \u2_Display/n3187 ;
  wire \u2_Display/n3188 ;
  wire \u2_Display/n3191 ;
  wire \u2_Display/n3192 ;
  wire \u2_Display/n3193 ;
  wire \u2_Display/n3194 ;
  wire \u2_Display/n3195 ;
  wire \u2_Display/n3196 ;
  wire \u2_Display/n3197 ;
  wire \u2_Display/n3198 ;
  wire \u2_Display/n3199 ;
  wire \u2_Display/n3200 ;
  wire \u2_Display/n3201 ;
  wire \u2_Display/n3202 ;
  wire \u2_Display/n3203 ;
  wire \u2_Display/n3204 ;
  wire \u2_Display/n3205 ;
  wire \u2_Display/n3206 ;
  wire \u2_Display/n3207 ;
  wire \u2_Display/n3208 ;
  wire \u2_Display/n3209 ;
  wire \u2_Display/n3210 ;
  wire \u2_Display/n3211 ;
  wire \u2_Display/n3212 ;
  wire \u2_Display/n3213 ;
  wire \u2_Display/n3214 ;
  wire \u2_Display/n3215 ;
  wire \u2_Display/n3216 ;
  wire \u2_Display/n3217 ;
  wire \u2_Display/n3218 ;
  wire \u2_Display/n3219 ;
  wire \u2_Display/n3220 ;
  wire \u2_Display/n3221 ;
  wire \u2_Display/n3222 ;
  wire \u2_Display/n3223 ;
  wire \u2_Display/n3226 ;
  wire \u2_Display/n3227 ;
  wire \u2_Display/n3228 ;
  wire \u2_Display/n3229 ;
  wire \u2_Display/n3230 ;
  wire \u2_Display/n3231 ;
  wire \u2_Display/n3232 ;
  wire \u2_Display/n3233 ;
  wire \u2_Display/n3234 ;
  wire \u2_Display/n3235 ;
  wire \u2_Display/n3236 ;
  wire \u2_Display/n3237 ;
  wire \u2_Display/n3238 ;
  wire \u2_Display/n3239 ;
  wire \u2_Display/n3240 ;
  wire \u2_Display/n3241 ;
  wire \u2_Display/n3242 ;
  wire \u2_Display/n3243 ;
  wire \u2_Display/n3244 ;
  wire \u2_Display/n3245 ;
  wire \u2_Display/n3246 ;
  wire \u2_Display/n3247 ;
  wire \u2_Display/n3248 ;
  wire \u2_Display/n3249 ;
  wire \u2_Display/n3250 ;
  wire \u2_Display/n3251 ;
  wire \u2_Display/n3252 ;
  wire \u2_Display/n3253 ;
  wire \u2_Display/n3254 ;
  wire \u2_Display/n3255 ;
  wire \u2_Display/n3256 ;
  wire \u2_Display/n3257 ;
  wire \u2_Display/n3258 ;
  wire \u2_Display/n3261 ;
  wire \u2_Display/n3262 ;
  wire \u2_Display/n3263 ;
  wire \u2_Display/n3264 ;
  wire \u2_Display/n3265 ;
  wire \u2_Display/n3266 ;
  wire \u2_Display/n3267 ;
  wire \u2_Display/n3268 ;
  wire \u2_Display/n3269 ;
  wire \u2_Display/n3270 ;
  wire \u2_Display/n3271 ;
  wire \u2_Display/n3272 ;
  wire \u2_Display/n3273 ;
  wire \u2_Display/n3274 ;
  wire \u2_Display/n3275 ;
  wire \u2_Display/n3276 ;
  wire \u2_Display/n3277 ;
  wire \u2_Display/n3278 ;
  wire \u2_Display/n3279 ;
  wire \u2_Display/n3280 ;
  wire \u2_Display/n3281 ;
  wire \u2_Display/n3282 ;
  wire \u2_Display/n3283 ;
  wire \u2_Display/n3284 ;
  wire \u2_Display/n3285 ;
  wire \u2_Display/n3286 ;
  wire \u2_Display/n3287 ;
  wire \u2_Display/n3288 ;
  wire \u2_Display/n3289 ;
  wire \u2_Display/n3290 ;
  wire \u2_Display/n3291 ;
  wire \u2_Display/n3292 ;
  wire \u2_Display/n3293 ;
  wire \u2_Display/n3296 ;
  wire \u2_Display/n3297 ;
  wire \u2_Display/n3298 ;
  wire \u2_Display/n3299 ;
  wire \u2_Display/n3300 ;
  wire \u2_Display/n3301 ;
  wire \u2_Display/n3302 ;
  wire \u2_Display/n3303 ;
  wire \u2_Display/n3304 ;
  wire \u2_Display/n3305 ;
  wire \u2_Display/n3306 ;
  wire \u2_Display/n3307 ;
  wire \u2_Display/n3308 ;
  wire \u2_Display/n3309 ;
  wire \u2_Display/n3310 ;
  wire \u2_Display/n3311 ;
  wire \u2_Display/n3312 ;
  wire \u2_Display/n3313 ;
  wire \u2_Display/n3314 ;
  wire \u2_Display/n3315 ;
  wire \u2_Display/n3316 ;
  wire \u2_Display/n3317 ;
  wire \u2_Display/n3318 ;
  wire \u2_Display/n3319 ;
  wire \u2_Display/n3320 ;
  wire \u2_Display/n3321 ;
  wire \u2_Display/n3322 ;
  wire \u2_Display/n3323 ;
  wire \u2_Display/n3324 ;
  wire \u2_Display/n3325 ;
  wire \u2_Display/n3326 ;
  wire \u2_Display/n3327 ;
  wire \u2_Display/n3328 ;
  wire \u2_Display/n3331 ;
  wire \u2_Display/n3332 ;
  wire \u2_Display/n3333 ;
  wire \u2_Display/n3334 ;
  wire \u2_Display/n3335 ;
  wire \u2_Display/n3336 ;
  wire \u2_Display/n3337 ;
  wire \u2_Display/n3338 ;
  wire \u2_Display/n3339 ;
  wire \u2_Display/n3340 ;
  wire \u2_Display/n3341 ;
  wire \u2_Display/n3342 ;
  wire \u2_Display/n3343 ;
  wire \u2_Display/n3344 ;
  wire \u2_Display/n3345 ;
  wire \u2_Display/n3346 ;
  wire \u2_Display/n3347 ;
  wire \u2_Display/n3348 ;
  wire \u2_Display/n3349 ;
  wire \u2_Display/n3350 ;
  wire \u2_Display/n3351 ;
  wire \u2_Display/n3352 ;
  wire \u2_Display/n3353 ;
  wire \u2_Display/n3354 ;
  wire \u2_Display/n3355 ;
  wire \u2_Display/n3356 ;
  wire \u2_Display/n3357 ;
  wire \u2_Display/n3358 ;
  wire \u2_Display/n3359 ;
  wire \u2_Display/n3360 ;
  wire \u2_Display/n3361 ;
  wire \u2_Display/n3362 ;
  wire \u2_Display/n3363 ;
  wire \u2_Display/n3366 ;
  wire \u2_Display/n3367 ;
  wire \u2_Display/n3368 ;
  wire \u2_Display/n3369 ;
  wire \u2_Display/n3370 ;
  wire \u2_Display/n3371 ;
  wire \u2_Display/n3372 ;
  wire \u2_Display/n3373 ;
  wire \u2_Display/n3374 ;
  wire \u2_Display/n3375 ;
  wire \u2_Display/n3376 ;
  wire \u2_Display/n3377 ;
  wire \u2_Display/n3378 ;
  wire \u2_Display/n3379 ;
  wire \u2_Display/n3380 ;
  wire \u2_Display/n3381 ;
  wire \u2_Display/n3382 ;
  wire \u2_Display/n3383 ;
  wire \u2_Display/n3384 ;
  wire \u2_Display/n3385 ;
  wire \u2_Display/n3386 ;
  wire \u2_Display/n3387 ;
  wire \u2_Display/n3388 ;
  wire \u2_Display/n3389 ;
  wire \u2_Display/n3390 ;
  wire \u2_Display/n3391 ;
  wire \u2_Display/n3392 ;
  wire \u2_Display/n3393 ;
  wire \u2_Display/n3394 ;
  wire \u2_Display/n3395 ;
  wire \u2_Display/n3396 ;
  wire \u2_Display/n3397 ;
  wire \u2_Display/n3398 ;
  wire \u2_Display/n3401 ;
  wire \u2_Display/n3402 ;
  wire \u2_Display/n3403 ;
  wire \u2_Display/n3404 ;
  wire \u2_Display/n3405 ;
  wire \u2_Display/n3406 ;
  wire \u2_Display/n3407 ;
  wire \u2_Display/n3408 ;
  wire \u2_Display/n3409 ;
  wire \u2_Display/n3410 ;
  wire \u2_Display/n3411 ;
  wire \u2_Display/n3412 ;
  wire \u2_Display/n3413 ;
  wire \u2_Display/n3414 ;
  wire \u2_Display/n3415 ;
  wire \u2_Display/n3416 ;
  wire \u2_Display/n3417 ;
  wire \u2_Display/n3418 ;
  wire \u2_Display/n3419 ;
  wire \u2_Display/n3420 ;
  wire \u2_Display/n3421 ;
  wire \u2_Display/n3422 ;
  wire \u2_Display/n3423 ;
  wire \u2_Display/n3424 ;
  wire \u2_Display/n3425 ;
  wire \u2_Display/n3426 ;
  wire \u2_Display/n3427 ;
  wire \u2_Display/n3428 ;
  wire \u2_Display/n3429 ;
  wire \u2_Display/n3430 ;
  wire \u2_Display/n3431 ;
  wire \u2_Display/n3432 ;
  wire \u2_Display/n3433 ;
  wire \u2_Display/n35 ;
  wire \u2_Display/n36 ;
  wire \u2_Display/n3786 ;
  wire \u2_Display/n3789 ;
  wire \u2_Display/n3790 ;
  wire \u2_Display/n3791 ;
  wire \u2_Display/n3792 ;
  wire \u2_Display/n3793 ;
  wire \u2_Display/n3794 ;
  wire \u2_Display/n3795 ;
  wire \u2_Display/n3796 ;
  wire \u2_Display/n3797 ;
  wire \u2_Display/n3798 ;
  wire \u2_Display/n3799 ;
  wire \u2_Display/n3800 ;
  wire \u2_Display/n3801 ;
  wire \u2_Display/n3802 ;
  wire \u2_Display/n3803 ;
  wire \u2_Display/n3804 ;
  wire \u2_Display/n3805 ;
  wire \u2_Display/n3806 ;
  wire \u2_Display/n3807 ;
  wire \u2_Display/n3808 ;
  wire \u2_Display/n3809 ;
  wire \u2_Display/n3810 ;
  wire \u2_Display/n3811 ;
  wire \u2_Display/n3812 ;
  wire \u2_Display/n3813 ;
  wire \u2_Display/n3814 ;
  wire \u2_Display/n3815 ;
  wire \u2_Display/n3816 ;
  wire \u2_Display/n3817 ;
  wire \u2_Display/n3818 ;
  wire \u2_Display/n3819 ;
  wire \u2_Display/n3820 ;
  wire \u2_Display/n3821 ;
  wire \u2_Display/n3824 ;
  wire \u2_Display/n3825 ;
  wire \u2_Display/n3826 ;
  wire \u2_Display/n3827 ;
  wire \u2_Display/n3828 ;
  wire \u2_Display/n3829 ;
  wire \u2_Display/n3830 ;
  wire \u2_Display/n3831 ;
  wire \u2_Display/n3832 ;
  wire \u2_Display/n3833 ;
  wire \u2_Display/n3834 ;
  wire \u2_Display/n3835 ;
  wire \u2_Display/n3836 ;
  wire \u2_Display/n3837 ;
  wire \u2_Display/n3838 ;
  wire \u2_Display/n3839 ;
  wire \u2_Display/n3840 ;
  wire \u2_Display/n3841 ;
  wire \u2_Display/n3842 ;
  wire \u2_Display/n3843 ;
  wire \u2_Display/n3844 ;
  wire \u2_Display/n3845 ;
  wire \u2_Display/n3846 ;
  wire \u2_Display/n3847 ;
  wire \u2_Display/n3848 ;
  wire \u2_Display/n3849 ;
  wire \u2_Display/n3850 ;
  wire \u2_Display/n3851 ;
  wire \u2_Display/n3852 ;
  wire \u2_Display/n3853 ;
  wire \u2_Display/n3854 ;
  wire \u2_Display/n3855 ;
  wire \u2_Display/n3856 ;
  wire \u2_Display/n3859 ;
  wire \u2_Display/n3860 ;
  wire \u2_Display/n3861 ;
  wire \u2_Display/n3862 ;
  wire \u2_Display/n3863 ;
  wire \u2_Display/n3864 ;
  wire \u2_Display/n3865 ;
  wire \u2_Display/n3866 ;
  wire \u2_Display/n3867 ;
  wire \u2_Display/n3868 ;
  wire \u2_Display/n3869 ;
  wire \u2_Display/n3870 ;
  wire \u2_Display/n3871 ;
  wire \u2_Display/n3872 ;
  wire \u2_Display/n3873 ;
  wire \u2_Display/n3874 ;
  wire \u2_Display/n3875 ;
  wire \u2_Display/n3876 ;
  wire \u2_Display/n3877 ;
  wire \u2_Display/n3878 ;
  wire \u2_Display/n3879 ;
  wire \u2_Display/n3880 ;
  wire \u2_Display/n3881 ;
  wire \u2_Display/n3882 ;
  wire \u2_Display/n3883 ;
  wire \u2_Display/n3884 ;
  wire \u2_Display/n3885 ;
  wire \u2_Display/n3886 ;
  wire \u2_Display/n3887 ;
  wire \u2_Display/n3888 ;
  wire \u2_Display/n3889 ;
  wire \u2_Display/n3890 ;
  wire \u2_Display/n3891 ;
  wire \u2_Display/n3894 ;
  wire \u2_Display/n3895 ;
  wire \u2_Display/n3896 ;
  wire \u2_Display/n3897 ;
  wire \u2_Display/n3898 ;
  wire \u2_Display/n3899 ;
  wire \u2_Display/n3900 ;
  wire \u2_Display/n3901 ;
  wire \u2_Display/n3902 ;
  wire \u2_Display/n3903 ;
  wire \u2_Display/n3904 ;
  wire \u2_Display/n3905 ;
  wire \u2_Display/n3906 ;
  wire \u2_Display/n3907 ;
  wire \u2_Display/n3908 ;
  wire \u2_Display/n3909 ;
  wire \u2_Display/n3910 ;
  wire \u2_Display/n3911 ;
  wire \u2_Display/n3912 ;
  wire \u2_Display/n3913 ;
  wire \u2_Display/n3914 ;
  wire \u2_Display/n3915 ;
  wire \u2_Display/n3916 ;
  wire \u2_Display/n3917 ;
  wire \u2_Display/n3918 ;
  wire \u2_Display/n3919 ;
  wire \u2_Display/n3920 ;
  wire \u2_Display/n3921 ;
  wire \u2_Display/n3922 ;
  wire \u2_Display/n3923 ;
  wire \u2_Display/n3924 ;
  wire \u2_Display/n3925 ;
  wire \u2_Display/n3926 ;
  wire \u2_Display/n3929 ;
  wire \u2_Display/n3930 ;
  wire \u2_Display/n3931 ;
  wire \u2_Display/n3932 ;
  wire \u2_Display/n3933 ;
  wire \u2_Display/n3934 ;
  wire \u2_Display/n3935 ;
  wire \u2_Display/n3936 ;
  wire \u2_Display/n3937 ;
  wire \u2_Display/n3938 ;
  wire \u2_Display/n3939 ;
  wire \u2_Display/n3940 ;
  wire \u2_Display/n3941 ;
  wire \u2_Display/n3942 ;
  wire \u2_Display/n3943 ;
  wire \u2_Display/n3944 ;
  wire \u2_Display/n3945 ;
  wire \u2_Display/n3946 ;
  wire \u2_Display/n3947 ;
  wire \u2_Display/n3948 ;
  wire \u2_Display/n3949 ;
  wire \u2_Display/n3950 ;
  wire \u2_Display/n3951 ;
  wire \u2_Display/n3952 ;
  wire \u2_Display/n3953 ;
  wire \u2_Display/n3954 ;
  wire \u2_Display/n3955 ;
  wire \u2_Display/n3956 ;
  wire \u2_Display/n3957 ;
  wire \u2_Display/n3958 ;
  wire \u2_Display/n3959 ;
  wire \u2_Display/n3960 ;
  wire \u2_Display/n3961 ;
  wire \u2_Display/n3964 ;
  wire \u2_Display/n3965 ;
  wire \u2_Display/n3966 ;
  wire \u2_Display/n3967 ;
  wire \u2_Display/n3968 ;
  wire \u2_Display/n3969 ;
  wire \u2_Display/n3970 ;
  wire \u2_Display/n3971 ;
  wire \u2_Display/n3972 ;
  wire \u2_Display/n3973 ;
  wire \u2_Display/n3974 ;
  wire \u2_Display/n3975 ;
  wire \u2_Display/n3976 ;
  wire \u2_Display/n3977 ;
  wire \u2_Display/n3978 ;
  wire \u2_Display/n3979 ;
  wire \u2_Display/n3980 ;
  wire \u2_Display/n3981 ;
  wire \u2_Display/n3982 ;
  wire \u2_Display/n3983 ;
  wire \u2_Display/n3984 ;
  wire \u2_Display/n3985 ;
  wire \u2_Display/n3986 ;
  wire \u2_Display/n3987 ;
  wire \u2_Display/n3988 ;
  wire \u2_Display/n3989 ;
  wire \u2_Display/n3990 ;
  wire \u2_Display/n3991 ;
  wire \u2_Display/n3992 ;
  wire \u2_Display/n3993 ;
  wire \u2_Display/n3994 ;
  wire \u2_Display/n3995 ;
  wire \u2_Display/n3996 ;
  wire \u2_Display/n3999 ;
  wire \u2_Display/n4000 ;
  wire \u2_Display/n4001 ;
  wire \u2_Display/n4002 ;
  wire \u2_Display/n4003 ;
  wire \u2_Display/n4004 ;
  wire \u2_Display/n4005 ;
  wire \u2_Display/n4006 ;
  wire \u2_Display/n4007 ;
  wire \u2_Display/n4008 ;
  wire \u2_Display/n4009 ;
  wire \u2_Display/n4010 ;
  wire \u2_Display/n4011 ;
  wire \u2_Display/n4012 ;
  wire \u2_Display/n4013 ;
  wire \u2_Display/n4014 ;
  wire \u2_Display/n4015 ;
  wire \u2_Display/n4016 ;
  wire \u2_Display/n4017 ;
  wire \u2_Display/n4018 ;
  wire \u2_Display/n4019 ;
  wire \u2_Display/n4020 ;
  wire \u2_Display/n4021 ;
  wire \u2_Display/n4022 ;
  wire \u2_Display/n4023 ;
  wire \u2_Display/n4024 ;
  wire \u2_Display/n4025 ;
  wire \u2_Display/n4026 ;
  wire \u2_Display/n4027 ;
  wire \u2_Display/n4028 ;
  wire \u2_Display/n4029 ;
  wire \u2_Display/n4030 ;
  wire \u2_Display/n4031 ;
  wire \u2_Display/n4034 ;
  wire \u2_Display/n4035 ;
  wire \u2_Display/n4036 ;
  wire \u2_Display/n4037 ;
  wire \u2_Display/n4038 ;
  wire \u2_Display/n4039 ;
  wire \u2_Display/n4040 ;
  wire \u2_Display/n4041 ;
  wire \u2_Display/n4042 ;
  wire \u2_Display/n4043 ;
  wire \u2_Display/n4044 ;
  wire \u2_Display/n4045 ;
  wire \u2_Display/n4046 ;
  wire \u2_Display/n4047 ;
  wire \u2_Display/n4048 ;
  wire \u2_Display/n4049 ;
  wire \u2_Display/n4050 ;
  wire \u2_Display/n4051 ;
  wire \u2_Display/n4052 ;
  wire \u2_Display/n4053 ;
  wire \u2_Display/n4054 ;
  wire \u2_Display/n4055 ;
  wire \u2_Display/n4056 ;
  wire \u2_Display/n4057 ;
  wire \u2_Display/n4058 ;
  wire \u2_Display/n4059 ;
  wire \u2_Display/n4060 ;
  wire \u2_Display/n4061 ;
  wire \u2_Display/n4062 ;
  wire \u2_Display/n4063 ;
  wire \u2_Display/n4064 ;
  wire \u2_Display/n4065 ;
  wire \u2_Display/n4066 ;
  wire \u2_Display/n4069 ;
  wire \u2_Display/n4070 ;
  wire \u2_Display/n4071 ;
  wire \u2_Display/n4072 ;
  wire \u2_Display/n4073 ;
  wire \u2_Display/n4074 ;
  wire \u2_Display/n4075 ;
  wire \u2_Display/n4076 ;
  wire \u2_Display/n4077 ;
  wire \u2_Display/n4078 ;
  wire \u2_Display/n4079 ;
  wire \u2_Display/n4080 ;
  wire \u2_Display/n4081 ;
  wire \u2_Display/n4082 ;
  wire \u2_Display/n4083 ;
  wire \u2_Display/n4084 ;
  wire \u2_Display/n4085 ;
  wire \u2_Display/n4086 ;
  wire \u2_Display/n4087 ;
  wire \u2_Display/n4088 ;
  wire \u2_Display/n4089 ;
  wire \u2_Display/n4090 ;
  wire \u2_Display/n4091 ;
  wire \u2_Display/n4092 ;
  wire \u2_Display/n4093 ;
  wire \u2_Display/n4094 ;
  wire \u2_Display/n4095 ;
  wire \u2_Display/n4096 ;
  wire \u2_Display/n4097 ;
  wire \u2_Display/n4098 ;
  wire \u2_Display/n4099 ;
  wire \u2_Display/n4100 ;
  wire \u2_Display/n4101 ;
  wire \u2_Display/n4104 ;
  wire \u2_Display/n4105 ;
  wire \u2_Display/n4106 ;
  wire \u2_Display/n4107 ;
  wire \u2_Display/n4108 ;
  wire \u2_Display/n4109 ;
  wire \u2_Display/n4110 ;
  wire \u2_Display/n4111 ;
  wire \u2_Display/n4112 ;
  wire \u2_Display/n4113 ;
  wire \u2_Display/n4114 ;
  wire \u2_Display/n4115 ;
  wire \u2_Display/n4116 ;
  wire \u2_Display/n4117 ;
  wire \u2_Display/n4118 ;
  wire \u2_Display/n4119 ;
  wire \u2_Display/n4120 ;
  wire \u2_Display/n4121 ;
  wire \u2_Display/n4122 ;
  wire \u2_Display/n4123 ;
  wire \u2_Display/n4124 ;
  wire \u2_Display/n4125 ;
  wire \u2_Display/n4126 ;
  wire \u2_Display/n4127 ;
  wire \u2_Display/n4128 ;
  wire \u2_Display/n4129 ;
  wire \u2_Display/n4130 ;
  wire \u2_Display/n4131 ;
  wire \u2_Display/n4132 ;
  wire \u2_Display/n4133 ;
  wire \u2_Display/n4134 ;
  wire \u2_Display/n4135 ;
  wire \u2_Display/n4136 ;
  wire \u2_Display/n4139 ;
  wire \u2_Display/n4140 ;
  wire \u2_Display/n4141 ;
  wire \u2_Display/n4142 ;
  wire \u2_Display/n4143 ;
  wire \u2_Display/n4144 ;
  wire \u2_Display/n4145 ;
  wire \u2_Display/n4146 ;
  wire \u2_Display/n4147 ;
  wire \u2_Display/n4148 ;
  wire \u2_Display/n4149 ;
  wire \u2_Display/n4150 ;
  wire \u2_Display/n4151 ;
  wire \u2_Display/n4152 ;
  wire \u2_Display/n4153 ;
  wire \u2_Display/n4154 ;
  wire \u2_Display/n4155 ;
  wire \u2_Display/n4156 ;
  wire \u2_Display/n4157 ;
  wire \u2_Display/n4158 ;
  wire \u2_Display/n4159 ;
  wire \u2_Display/n4160 ;
  wire \u2_Display/n4161 ;
  wire \u2_Display/n4162 ;
  wire \u2_Display/n4163 ;
  wire \u2_Display/n4164 ;
  wire \u2_Display/n4165 ;
  wire \u2_Display/n4166 ;
  wire \u2_Display/n4167 ;
  wire \u2_Display/n4168 ;
  wire \u2_Display/n4169 ;
  wire \u2_Display/n417 ;
  wire \u2_Display/n4170 ;
  wire \u2_Display/n4171 ;
  wire \u2_Display/n4174 ;
  wire \u2_Display/n4175 ;
  wire \u2_Display/n4176 ;
  wire \u2_Display/n4177 ;
  wire \u2_Display/n4178 ;
  wire \u2_Display/n4179 ;
  wire \u2_Display/n4180 ;
  wire \u2_Display/n4181 ;
  wire \u2_Display/n4182 ;
  wire \u2_Display/n4183 ;
  wire \u2_Display/n4184 ;
  wire \u2_Display/n4185 ;
  wire \u2_Display/n4186 ;
  wire \u2_Display/n4187 ;
  wire \u2_Display/n4188 ;
  wire \u2_Display/n4189 ;
  wire \u2_Display/n4190 ;
  wire \u2_Display/n4191 ;
  wire \u2_Display/n4192 ;
  wire \u2_Display/n4193 ;
  wire \u2_Display/n4194 ;
  wire \u2_Display/n4195 ;
  wire \u2_Display/n4196 ;
  wire \u2_Display/n4197 ;
  wire \u2_Display/n4198 ;
  wire \u2_Display/n4199 ;
  wire \u2_Display/n420 ;
  wire \u2_Display/n4200 ;
  wire \u2_Display/n4201 ;
  wire \u2_Display/n4202 ;
  wire \u2_Display/n4203 ;
  wire \u2_Display/n4204 ;
  wire \u2_Display/n4205 ;
  wire \u2_Display/n4206 ;
  wire \u2_Display/n4209 ;
  wire \u2_Display/n421 ;
  wire \u2_Display/n4210 ;
  wire \u2_Display/n4211 ;
  wire \u2_Display/n4212 ;
  wire \u2_Display/n4213 ;
  wire \u2_Display/n4214 ;
  wire \u2_Display/n4215 ;
  wire \u2_Display/n4216 ;
  wire \u2_Display/n4217 ;
  wire \u2_Display/n4218 ;
  wire \u2_Display/n4219 ;
  wire \u2_Display/n422 ;
  wire \u2_Display/n4220 ;
  wire \u2_Display/n4221 ;
  wire \u2_Display/n4222 ;
  wire \u2_Display/n4223 ;
  wire \u2_Display/n4224 ;
  wire \u2_Display/n4225 ;
  wire \u2_Display/n4226 ;
  wire \u2_Display/n4227 ;
  wire \u2_Display/n4228 ;
  wire \u2_Display/n4229 ;
  wire \u2_Display/n423 ;
  wire \u2_Display/n4230 ;
  wire \u2_Display/n4231 ;
  wire \u2_Display/n4232 ;
  wire \u2_Display/n4233 ;
  wire \u2_Display/n4234 ;
  wire \u2_Display/n4235 ;
  wire \u2_Display/n4236 ;
  wire \u2_Display/n4237 ;
  wire \u2_Display/n4238 ;
  wire \u2_Display/n4239 ;
  wire \u2_Display/n424 ;
  wire \u2_Display/n4240 ;
  wire \u2_Display/n4241 ;
  wire \u2_Display/n4244 ;
  wire \u2_Display/n4245 ;
  wire \u2_Display/n4246 ;
  wire \u2_Display/n4247 ;
  wire \u2_Display/n4248 ;
  wire \u2_Display/n4249 ;
  wire \u2_Display/n425 ;
  wire \u2_Display/n4250 ;
  wire \u2_Display/n4251 ;
  wire \u2_Display/n4252 ;
  wire \u2_Display/n4253 ;
  wire \u2_Display/n4254 ;
  wire \u2_Display/n4255 ;
  wire \u2_Display/n4256 ;
  wire \u2_Display/n4257 ;
  wire \u2_Display/n4258 ;
  wire \u2_Display/n4259 ;
  wire \u2_Display/n426 ;
  wire \u2_Display/n4260 ;
  wire \u2_Display/n4261 ;
  wire \u2_Display/n4262 ;
  wire \u2_Display/n4263 ;
  wire \u2_Display/n4264 ;
  wire \u2_Display/n4265 ;
  wire \u2_Display/n4266 ;
  wire \u2_Display/n4267 ;
  wire \u2_Display/n4268 ;
  wire \u2_Display/n4269 ;
  wire \u2_Display/n427 ;
  wire \u2_Display/n4270 ;
  wire \u2_Display/n4271 ;
  wire \u2_Display/n4272 ;
  wire \u2_Display/n4273 ;
  wire \u2_Display/n4274 ;
  wire \u2_Display/n4275 ;
  wire \u2_Display/n4276 ;
  wire \u2_Display/n4279 ;
  wire \u2_Display/n428 ;
  wire \u2_Display/n4280 ;
  wire \u2_Display/n4281 ;
  wire \u2_Display/n4282 ;
  wire \u2_Display/n4283 ;
  wire \u2_Display/n4284 ;
  wire \u2_Display/n4285 ;
  wire \u2_Display/n4286 ;
  wire \u2_Display/n4287 ;
  wire \u2_Display/n4288 ;
  wire \u2_Display/n4289 ;
  wire \u2_Display/n429 ;
  wire \u2_Display/n4290 ;
  wire \u2_Display/n4291 ;
  wire \u2_Display/n4292 ;
  wire \u2_Display/n4293 ;
  wire \u2_Display/n4294 ;
  wire \u2_Display/n4295 ;
  wire \u2_Display/n4296 ;
  wire \u2_Display/n4297 ;
  wire \u2_Display/n4298 ;
  wire \u2_Display/n4299 ;
  wire \u2_Display/n430 ;
  wire \u2_Display/n4300 ;
  wire \u2_Display/n4301 ;
  wire \u2_Display/n4302 ;
  wire \u2_Display/n4303 ;
  wire \u2_Display/n4304 ;
  wire \u2_Display/n4305 ;
  wire \u2_Display/n4306 ;
  wire \u2_Display/n4307 ;
  wire \u2_Display/n4308 ;
  wire \u2_Display/n4309 ;
  wire \u2_Display/n431 ;
  wire \u2_Display/n4310 ;
  wire \u2_Display/n4311 ;
  wire \u2_Display/n4314 ;
  wire \u2_Display/n4315 ;
  wire \u2_Display/n4316 ;
  wire \u2_Display/n4317 ;
  wire \u2_Display/n4318 ;
  wire \u2_Display/n4319 ;
  wire \u2_Display/n432 ;
  wire \u2_Display/n4320 ;
  wire \u2_Display/n4321 ;
  wire \u2_Display/n4322 ;
  wire \u2_Display/n4323 ;
  wire \u2_Display/n4324 ;
  wire \u2_Display/n4325 ;
  wire \u2_Display/n4326 ;
  wire \u2_Display/n4327 ;
  wire \u2_Display/n4328 ;
  wire \u2_Display/n4329 ;
  wire \u2_Display/n433 ;
  wire \u2_Display/n4330 ;
  wire \u2_Display/n4331 ;
  wire \u2_Display/n4332 ;
  wire \u2_Display/n4333 ;
  wire \u2_Display/n4334 ;
  wire \u2_Display/n4335 ;
  wire \u2_Display/n4336 ;
  wire \u2_Display/n4337 ;
  wire \u2_Display/n4338 ;
  wire \u2_Display/n4339 ;
  wire \u2_Display/n434 ;
  wire \u2_Display/n4340 ;
  wire \u2_Display/n4341 ;
  wire \u2_Display/n4342 ;
  wire \u2_Display/n4343 ;
  wire \u2_Display/n4344 ;
  wire \u2_Display/n4345 ;
  wire \u2_Display/n4346 ;
  wire \u2_Display/n4349 ;
  wire \u2_Display/n435 ;
  wire \u2_Display/n4350 ;
  wire \u2_Display/n4351 ;
  wire \u2_Display/n4352 ;
  wire \u2_Display/n4353 ;
  wire \u2_Display/n4354 ;
  wire \u2_Display/n4355 ;
  wire \u2_Display/n4356 ;
  wire \u2_Display/n4357 ;
  wire \u2_Display/n4358 ;
  wire \u2_Display/n4359 ;
  wire \u2_Display/n436 ;
  wire \u2_Display/n4360 ;
  wire \u2_Display/n4361 ;
  wire \u2_Display/n4362 ;
  wire \u2_Display/n4363 ;
  wire \u2_Display/n4364 ;
  wire \u2_Display/n4365 ;
  wire \u2_Display/n4366 ;
  wire \u2_Display/n4367 ;
  wire \u2_Display/n4368 ;
  wire \u2_Display/n4369 ;
  wire \u2_Display/n437 ;
  wire \u2_Display/n4370 ;
  wire \u2_Display/n4371 ;
  wire \u2_Display/n4372 ;
  wire \u2_Display/n4373 ;
  wire \u2_Display/n4374 ;
  wire \u2_Display/n4375 ;
  wire \u2_Display/n4376 ;
  wire \u2_Display/n4377 ;
  wire \u2_Display/n4378 ;
  wire \u2_Display/n4379 ;
  wire \u2_Display/n438 ;
  wire \u2_Display/n4380 ;
  wire \u2_Display/n4381 ;
  wire \u2_Display/n4384 ;
  wire \u2_Display/n4385 ;
  wire \u2_Display/n4386 ;
  wire \u2_Display/n4387 ;
  wire \u2_Display/n4388 ;
  wire \u2_Display/n4389 ;
  wire \u2_Display/n439 ;
  wire \u2_Display/n4390 ;
  wire \u2_Display/n4391 ;
  wire \u2_Display/n4392 ;
  wire \u2_Display/n4393 ;
  wire \u2_Display/n4394 ;
  wire \u2_Display/n4395 ;
  wire \u2_Display/n4396 ;
  wire \u2_Display/n4397 ;
  wire \u2_Display/n4398 ;
  wire \u2_Display/n4399 ;
  wire \u2_Display/n44 ;
  wire \u2_Display/n440 ;
  wire \u2_Display/n4400 ;
  wire \u2_Display/n4401 ;
  wire \u2_Display/n4402 ;
  wire \u2_Display/n4403 ;
  wire \u2_Display/n4404 ;
  wire \u2_Display/n4405 ;
  wire \u2_Display/n4406 ;
  wire \u2_Display/n4407 ;
  wire \u2_Display/n4408 ;
  wire \u2_Display/n4409 ;
  wire \u2_Display/n441 ;
  wire \u2_Display/n4410 ;
  wire \u2_Display/n4411 ;
  wire \u2_Display/n4412 ;
  wire \u2_Display/n4413 ;
  wire \u2_Display/n4414 ;
  wire \u2_Display/n4415 ;
  wire \u2_Display/n4416 ;
  wire \u2_Display/n4419 ;
  wire \u2_Display/n442 ;
  wire \u2_Display/n4420 ;
  wire \u2_Display/n4421 ;
  wire \u2_Display/n4422 ;
  wire \u2_Display/n4423 ;
  wire \u2_Display/n4424 ;
  wire \u2_Display/n4425 ;
  wire \u2_Display/n4426 ;
  wire \u2_Display/n4427 ;
  wire \u2_Display/n4428 ;
  wire \u2_Display/n4429 ;
  wire \u2_Display/n443 ;
  wire \u2_Display/n4430 ;
  wire \u2_Display/n4431 ;
  wire \u2_Display/n4432 ;
  wire \u2_Display/n4433 ;
  wire \u2_Display/n4434 ;
  wire \u2_Display/n4435 ;
  wire \u2_Display/n4436 ;
  wire \u2_Display/n4437 ;
  wire \u2_Display/n4438 ;
  wire \u2_Display/n4439 ;
  wire \u2_Display/n444 ;
  wire \u2_Display/n4440 ;
  wire \u2_Display/n4441 ;
  wire \u2_Display/n4442 ;
  wire \u2_Display/n4443 ;
  wire \u2_Display/n4444 ;
  wire \u2_Display/n4445 ;
  wire \u2_Display/n4446 ;
  wire \u2_Display/n4447 ;
  wire \u2_Display/n4448 ;
  wire \u2_Display/n4449 ;
  wire \u2_Display/n445 ;
  wire \u2_Display/n4450 ;
  wire \u2_Display/n4451 ;
  wire \u2_Display/n4454 ;
  wire \u2_Display/n4455 ;
  wire \u2_Display/n4456 ;
  wire \u2_Display/n4457 ;
  wire \u2_Display/n4458 ;
  wire \u2_Display/n4459 ;
  wire \u2_Display/n446 ;
  wire \u2_Display/n4460 ;
  wire \u2_Display/n4461 ;
  wire \u2_Display/n4462 ;
  wire \u2_Display/n4463 ;
  wire \u2_Display/n4464 ;
  wire \u2_Display/n4465 ;
  wire \u2_Display/n4466 ;
  wire \u2_Display/n4467 ;
  wire \u2_Display/n4468 ;
  wire \u2_Display/n4469 ;
  wire \u2_Display/n447 ;
  wire \u2_Display/n4470 ;
  wire \u2_Display/n4471 ;
  wire \u2_Display/n4472 ;
  wire \u2_Display/n4473 ;
  wire \u2_Display/n4474 ;
  wire \u2_Display/n4475 ;
  wire \u2_Display/n4476 ;
  wire \u2_Display/n4477 ;
  wire \u2_Display/n4478 ;
  wire \u2_Display/n4479 ;
  wire \u2_Display/n448 ;
  wire \u2_Display/n4480 ;
  wire \u2_Display/n4481 ;
  wire \u2_Display/n4482 ;
  wire \u2_Display/n4483 ;
  wire \u2_Display/n4484 ;
  wire \u2_Display/n4485 ;
  wire \u2_Display/n4486 ;
  wire \u2_Display/n4489 ;
  wire \u2_Display/n449 ;
  wire \u2_Display/n4490 ;
  wire \u2_Display/n4491 ;
  wire \u2_Display/n4492 ;
  wire \u2_Display/n4493 ;
  wire \u2_Display/n4494 ;
  wire \u2_Display/n4495 ;
  wire \u2_Display/n4496 ;
  wire \u2_Display/n4497 ;
  wire \u2_Display/n4498 ;
  wire \u2_Display/n4499 ;
  wire \u2_Display/n45 ;
  wire \u2_Display/n450 ;
  wire \u2_Display/n4500 ;
  wire \u2_Display/n4501 ;
  wire \u2_Display/n4502 ;
  wire \u2_Display/n4503 ;
  wire \u2_Display/n4504 ;
  wire \u2_Display/n4505 ;
  wire \u2_Display/n4506 ;
  wire \u2_Display/n4507 ;
  wire \u2_Display/n4508 ;
  wire \u2_Display/n4509 ;
  wire \u2_Display/n451 ;
  wire \u2_Display/n4510 ;
  wire \u2_Display/n4511 ;
  wire \u2_Display/n4512 ;
  wire \u2_Display/n4513 ;
  wire \u2_Display/n4514 ;
  wire \u2_Display/n4515 ;
  wire \u2_Display/n4516 ;
  wire \u2_Display/n4517 ;
  wire \u2_Display/n4518 ;
  wire \u2_Display/n4519 ;
  wire \u2_Display/n452 ;
  wire \u2_Display/n4520 ;
  wire \u2_Display/n4521 ;
  wire \u2_Display/n4524 ;
  wire \u2_Display/n4525 ;
  wire \u2_Display/n4526 ;
  wire \u2_Display/n4527 ;
  wire \u2_Display/n4528 ;
  wire \u2_Display/n4529 ;
  wire \u2_Display/n4530 ;
  wire \u2_Display/n4531 ;
  wire \u2_Display/n4532 ;
  wire \u2_Display/n4533 ;
  wire \u2_Display/n4534 ;
  wire \u2_Display/n4535 ;
  wire \u2_Display/n4536 ;
  wire \u2_Display/n4537 ;
  wire \u2_Display/n4538 ;
  wire \u2_Display/n4539 ;
  wire \u2_Display/n4540 ;
  wire \u2_Display/n4541 ;
  wire \u2_Display/n4542 ;
  wire \u2_Display/n4543 ;
  wire \u2_Display/n4544 ;
  wire \u2_Display/n4545 ;
  wire \u2_Display/n4546 ;
  wire \u2_Display/n4547 ;
  wire \u2_Display/n4548 ;
  wire \u2_Display/n4549 ;
  wire \u2_Display/n455 ;
  wire \u2_Display/n4550 ;
  wire \u2_Display/n4551 ;
  wire \u2_Display/n4552 ;
  wire \u2_Display/n4553 ;
  wire \u2_Display/n4554 ;
  wire \u2_Display/n4555 ;
  wire \u2_Display/n4556 ;
  wire \u2_Display/n456 ;
  wire \u2_Display/n457 ;
  wire \u2_Display/n458 ;
  wire \u2_Display/n459 ;
  wire \u2_Display/n460 ;
  wire \u2_Display/n461 ;
  wire \u2_Display/n462 ;
  wire \u2_Display/n463 ;
  wire \u2_Display/n464 ;
  wire \u2_Display/n465 ;
  wire \u2_Display/n466 ;
  wire \u2_Display/n467 ;
  wire \u2_Display/n468 ;
  wire \u2_Display/n469 ;
  wire \u2_Display/n470 ;
  wire \u2_Display/n471 ;
  wire \u2_Display/n472 ;
  wire \u2_Display/n473 ;
  wire \u2_Display/n474 ;
  wire \u2_Display/n475 ;
  wire \u2_Display/n476 ;
  wire \u2_Display/n477 ;
  wire \u2_Display/n478 ;
  wire \u2_Display/n479 ;
  wire \u2_Display/n48 ;
  wire \u2_Display/n480 ;
  wire \u2_Display/n481 ;
  wire \u2_Display/n482 ;
  wire \u2_Display/n483 ;
  wire \u2_Display/n484 ;
  wire \u2_Display/n485 ;
  wire \u2_Display/n486 ;
  wire \u2_Display/n487 ;
  wire \u2_Display/n490 ;
  wire \u2_Display/n4909 ;
  wire \u2_Display/n491 ;
  wire \u2_Display/n492 ;
  wire \u2_Display/n493 ;
  wire \u2_Display/n494 ;
  wire \u2_Display/n4944 ;
  wire \u2_Display/n495 ;
  wire \u2_Display/n496 ;
  wire \u2_Display/n497 ;
  wire \u2_Display/n4979 ;
  wire \u2_Display/n498 ;
  wire \u2_Display/n499 ;
  wire \u2_Display/n50 ;
  wire \u2_Display/n500 ;
  wire \u2_Display/n501 ;
  wire \u2_Display/n5014 ;
  wire \u2_Display/n502 ;
  wire \u2_Display/n503 ;
  wire \u2_Display/n504 ;
  wire \u2_Display/n5049 ;
  wire \u2_Display/n505 ;
  wire \u2_Display/n506 ;
  wire \u2_Display/n507 ;
  wire \u2_Display/n508 ;
  wire \u2_Display/n5084 ;
  wire \u2_Display/n509 ;
  wire \u2_Display/n51 ;
  wire \u2_Display/n510 ;
  wire \u2_Display/n511 ;
  wire \u2_Display/n5119 ;
  wire \u2_Display/n512 ;
  wire \u2_Display/n513 ;
  wire \u2_Display/n514 ;
  wire \u2_Display/n515 ;
  wire \u2_Display/n5154 ;
  wire \u2_Display/n516 ;
  wire \u2_Display/n517 ;
  wire \u2_Display/n518 ;
  wire \u2_Display/n5189 ;
  wire \u2_Display/n519 ;
  wire \u2_Display/n5196 ;
  wire \u2_Display/n5197 ;
  wire \u2_Display/n5198 ;
  wire \u2_Display/n5199 ;
  wire \u2_Display/n520 ;
  wire \u2_Display/n5200 ;
  wire \u2_Display/n5201 ;
  wire \u2_Display/n5202 ;
  wire \u2_Display/n5203 ;
  wire \u2_Display/n5204 ;
  wire \u2_Display/n5205 ;
  wire \u2_Display/n5206 ;
  wire \u2_Display/n5207 ;
  wire \u2_Display/n5208 ;
  wire \u2_Display/n5209 ;
  wire \u2_Display/n521 ;
  wire \u2_Display/n5210 ;
  wire \u2_Display/n5211 ;
  wire \u2_Display/n5212 ;
  wire \u2_Display/n5213 ;
  wire \u2_Display/n5214 ;
  wire \u2_Display/n5215 ;
  wire \u2_Display/n5216 ;
  wire \u2_Display/n5217 ;
  wire \u2_Display/n5218 ;
  wire \u2_Display/n5219 ;
  wire \u2_Display/n522 ;
  wire \u2_Display/n5220 ;
  wire \u2_Display/n5221 ;
  wire \u2_Display/n5222 ;
  wire \u2_Display/n5223 ;
  wire \u2_Display/n5224 ;
  wire \u2_Display/n5227 ;
  wire \u2_Display/n5228 ;
  wire \u2_Display/n5229 ;
  wire \u2_Display/n5230 ;
  wire \u2_Display/n5231 ;
  wire \u2_Display/n5232 ;
  wire \u2_Display/n5233 ;
  wire \u2_Display/n5234 ;
  wire \u2_Display/n5235 ;
  wire \u2_Display/n5236 ;
  wire \u2_Display/n5237 ;
  wire \u2_Display/n5238 ;
  wire \u2_Display/n5239 ;
  wire \u2_Display/n5240 ;
  wire \u2_Display/n5241 ;
  wire \u2_Display/n5242 ;
  wire \u2_Display/n5243 ;
  wire \u2_Display/n5244 ;
  wire \u2_Display/n5245 ;
  wire \u2_Display/n5246 ;
  wire \u2_Display/n5247 ;
  wire \u2_Display/n5248 ;
  wire \u2_Display/n5249 ;
  wire \u2_Display/n525 ;
  wire \u2_Display/n5250 ;
  wire \u2_Display/n5251 ;
  wire \u2_Display/n5252 ;
  wire \u2_Display/n5253 ;
  wire \u2_Display/n5254 ;
  wire \u2_Display/n5255 ;
  wire \u2_Display/n5256 ;
  wire \u2_Display/n5257 ;
  wire \u2_Display/n5258 ;
  wire \u2_Display/n5259 ;
  wire \u2_Display/n526 ;
  wire \u2_Display/n5262 ;
  wire \u2_Display/n5263 ;
  wire \u2_Display/n5264 ;
  wire \u2_Display/n5265 ;
  wire \u2_Display/n5266 ;
  wire \u2_Display/n5267 ;
  wire \u2_Display/n5268 ;
  wire \u2_Display/n5269 ;
  wire \u2_Display/n527 ;
  wire \u2_Display/n5270 ;
  wire \u2_Display/n5271 ;
  wire \u2_Display/n5272 ;
  wire \u2_Display/n5273 ;
  wire \u2_Display/n5274 ;
  wire \u2_Display/n5275 ;
  wire \u2_Display/n5276 ;
  wire \u2_Display/n5277 ;
  wire \u2_Display/n5278 ;
  wire \u2_Display/n5279 ;
  wire \u2_Display/n528 ;
  wire \u2_Display/n5280 ;
  wire \u2_Display/n5281 ;
  wire \u2_Display/n5282 ;
  wire \u2_Display/n5283 ;
  wire \u2_Display/n5284 ;
  wire \u2_Display/n5285 ;
  wire \u2_Display/n5286 ;
  wire \u2_Display/n5287 ;
  wire \u2_Display/n5288 ;
  wire \u2_Display/n5289 ;
  wire \u2_Display/n529 ;
  wire \u2_Display/n5290 ;
  wire \u2_Display/n5291 ;
  wire \u2_Display/n5292 ;
  wire \u2_Display/n5293 ;
  wire \u2_Display/n5294 ;
  wire \u2_Display/n5297 ;
  wire \u2_Display/n5298 ;
  wire \u2_Display/n5299 ;
  wire \u2_Display/n530 ;
  wire \u2_Display/n5300 ;
  wire \u2_Display/n5301 ;
  wire \u2_Display/n5302 ;
  wire \u2_Display/n5303 ;
  wire \u2_Display/n5304 ;
  wire \u2_Display/n5305 ;
  wire \u2_Display/n5306 ;
  wire \u2_Display/n5307 ;
  wire \u2_Display/n5308 ;
  wire \u2_Display/n5309 ;
  wire \u2_Display/n531 ;
  wire \u2_Display/n5310 ;
  wire \u2_Display/n5311 ;
  wire \u2_Display/n5312 ;
  wire \u2_Display/n5313 ;
  wire \u2_Display/n5314 ;
  wire \u2_Display/n5315 ;
  wire \u2_Display/n5316 ;
  wire \u2_Display/n5317 ;
  wire \u2_Display/n5318 ;
  wire \u2_Display/n5319 ;
  wire \u2_Display/n532 ;
  wire \u2_Display/n5320 ;
  wire \u2_Display/n5321 ;
  wire \u2_Display/n5322 ;
  wire \u2_Display/n5323 ;
  wire \u2_Display/n5324 ;
  wire \u2_Display/n5325 ;
  wire \u2_Display/n5326 ;
  wire \u2_Display/n5327 ;
  wire \u2_Display/n5328 ;
  wire \u2_Display/n5329 ;
  wire \u2_Display/n533 ;
  wire \u2_Display/n5332 ;
  wire \u2_Display/n5333 ;
  wire \u2_Display/n5334 ;
  wire \u2_Display/n5335 ;
  wire \u2_Display/n5336 ;
  wire \u2_Display/n5337 ;
  wire \u2_Display/n5338 ;
  wire \u2_Display/n5339 ;
  wire \u2_Display/n534 ;
  wire \u2_Display/n5340 ;
  wire \u2_Display/n5341 ;
  wire \u2_Display/n5342 ;
  wire \u2_Display/n5343 ;
  wire \u2_Display/n5344 ;
  wire \u2_Display/n5345 ;
  wire \u2_Display/n5346 ;
  wire \u2_Display/n5347 ;
  wire \u2_Display/n5348 ;
  wire \u2_Display/n5349 ;
  wire \u2_Display/n535 ;
  wire \u2_Display/n5350 ;
  wire \u2_Display/n5351 ;
  wire \u2_Display/n5352 ;
  wire \u2_Display/n5353 ;
  wire \u2_Display/n5354 ;
  wire \u2_Display/n5355 ;
  wire \u2_Display/n5356 ;
  wire \u2_Display/n5357 ;
  wire \u2_Display/n5358 ;
  wire \u2_Display/n5359 ;
  wire \u2_Display/n536 ;
  wire \u2_Display/n5360 ;
  wire \u2_Display/n5361 ;
  wire \u2_Display/n5362 ;
  wire \u2_Display/n5363 ;
  wire \u2_Display/n5364 ;
  wire \u2_Display/n5367 ;
  wire \u2_Display/n5368 ;
  wire \u2_Display/n5369 ;
  wire \u2_Display/n537 ;
  wire \u2_Display/n5370 ;
  wire \u2_Display/n5371 ;
  wire \u2_Display/n5372 ;
  wire \u2_Display/n5373 ;
  wire \u2_Display/n5374 ;
  wire \u2_Display/n5375 ;
  wire \u2_Display/n5376 ;
  wire \u2_Display/n5377 ;
  wire \u2_Display/n5378 ;
  wire \u2_Display/n5379 ;
  wire \u2_Display/n538 ;
  wire \u2_Display/n5380 ;
  wire \u2_Display/n5381 ;
  wire \u2_Display/n5382 ;
  wire \u2_Display/n5383 ;
  wire \u2_Display/n5384 ;
  wire \u2_Display/n5385 ;
  wire \u2_Display/n5386 ;
  wire \u2_Display/n5387 ;
  wire \u2_Display/n5388 ;
  wire \u2_Display/n5389 ;
  wire \u2_Display/n539 ;
  wire \u2_Display/n5390 ;
  wire \u2_Display/n5391 ;
  wire \u2_Display/n5392 ;
  wire \u2_Display/n5393 ;
  wire \u2_Display/n5394 ;
  wire \u2_Display/n5395 ;
  wire \u2_Display/n5396 ;
  wire \u2_Display/n5397 ;
  wire \u2_Display/n5398 ;
  wire \u2_Display/n5399 ;
  wire \u2_Display/n540 ;
  wire \u2_Display/n5402 ;
  wire \u2_Display/n5403 ;
  wire \u2_Display/n5404 ;
  wire \u2_Display/n5405 ;
  wire \u2_Display/n5406 ;
  wire \u2_Display/n5407 ;
  wire \u2_Display/n5408 ;
  wire \u2_Display/n5409 ;
  wire \u2_Display/n541 ;
  wire \u2_Display/n5410 ;
  wire \u2_Display/n5411 ;
  wire \u2_Display/n5412 ;
  wire \u2_Display/n5413 ;
  wire \u2_Display/n5414 ;
  wire \u2_Display/n5415 ;
  wire \u2_Display/n5416 ;
  wire \u2_Display/n5417 ;
  wire \u2_Display/n5418 ;
  wire \u2_Display/n5419 ;
  wire \u2_Display/n542 ;
  wire \u2_Display/n5420 ;
  wire \u2_Display/n5421 ;
  wire \u2_Display/n5422 ;
  wire \u2_Display/n5423 ;
  wire \u2_Display/n5424 ;
  wire \u2_Display/n5425 ;
  wire \u2_Display/n5426 ;
  wire \u2_Display/n5427 ;
  wire \u2_Display/n5428 ;
  wire \u2_Display/n5429 ;
  wire \u2_Display/n543 ;
  wire \u2_Display/n5430 ;
  wire \u2_Display/n5431 ;
  wire \u2_Display/n5432 ;
  wire \u2_Display/n5433 ;
  wire \u2_Display/n5434 ;
  wire \u2_Display/n5437 ;
  wire \u2_Display/n5438 ;
  wire \u2_Display/n5439 ;
  wire \u2_Display/n544 ;
  wire \u2_Display/n5440 ;
  wire \u2_Display/n5441 ;
  wire \u2_Display/n5442 ;
  wire \u2_Display/n5443 ;
  wire \u2_Display/n5444 ;
  wire \u2_Display/n5445 ;
  wire \u2_Display/n5446 ;
  wire \u2_Display/n5447 ;
  wire \u2_Display/n5448 ;
  wire \u2_Display/n5449 ;
  wire \u2_Display/n545 ;
  wire \u2_Display/n5450 ;
  wire \u2_Display/n5451 ;
  wire \u2_Display/n5452 ;
  wire \u2_Display/n5453 ;
  wire \u2_Display/n5454 ;
  wire \u2_Display/n5455 ;
  wire \u2_Display/n5456 ;
  wire \u2_Display/n5457 ;
  wire \u2_Display/n5458 ;
  wire \u2_Display/n5459 ;
  wire \u2_Display/n546 ;
  wire \u2_Display/n5460 ;
  wire \u2_Display/n5461 ;
  wire \u2_Display/n5462 ;
  wire \u2_Display/n5463 ;
  wire \u2_Display/n5464 ;
  wire \u2_Display/n5465 ;
  wire \u2_Display/n5466 ;
  wire \u2_Display/n5467 ;
  wire \u2_Display/n5468 ;
  wire \u2_Display/n5469 ;
  wire \u2_Display/n547 ;
  wire \u2_Display/n5472 ;
  wire \u2_Display/n5473 ;
  wire \u2_Display/n5474 ;
  wire \u2_Display/n5475 ;
  wire \u2_Display/n5476 ;
  wire \u2_Display/n5477 ;
  wire \u2_Display/n5478 ;
  wire \u2_Display/n5479 ;
  wire \u2_Display/n548 ;
  wire \u2_Display/n5480 ;
  wire \u2_Display/n5481 ;
  wire \u2_Display/n5482 ;
  wire \u2_Display/n5483 ;
  wire \u2_Display/n5484 ;
  wire \u2_Display/n5485 ;
  wire \u2_Display/n5486 ;
  wire \u2_Display/n5487 ;
  wire \u2_Display/n5488 ;
  wire \u2_Display/n5489 ;
  wire \u2_Display/n549 ;
  wire \u2_Display/n5490 ;
  wire \u2_Display/n5491 ;
  wire \u2_Display/n5492 ;
  wire \u2_Display/n5493 ;
  wire \u2_Display/n5494 ;
  wire \u2_Display/n5495 ;
  wire \u2_Display/n5496 ;
  wire \u2_Display/n5497 ;
  wire \u2_Display/n5498 ;
  wire \u2_Display/n5499 ;
  wire \u2_Display/n550 ;
  wire \u2_Display/n5500 ;
  wire \u2_Display/n5501 ;
  wire \u2_Display/n5502 ;
  wire \u2_Display/n5503 ;
  wire \u2_Display/n5504 ;
  wire \u2_Display/n5507 ;
  wire \u2_Display/n5508 ;
  wire \u2_Display/n5509 ;
  wire \u2_Display/n551 ;
  wire \u2_Display/n5510 ;
  wire \u2_Display/n5511 ;
  wire \u2_Display/n5512 ;
  wire \u2_Display/n5513 ;
  wire \u2_Display/n5514 ;
  wire \u2_Display/n5515 ;
  wire \u2_Display/n5516 ;
  wire \u2_Display/n5517 ;
  wire \u2_Display/n5518 ;
  wire \u2_Display/n5519 ;
  wire \u2_Display/n552 ;
  wire \u2_Display/n5520 ;
  wire \u2_Display/n5521 ;
  wire \u2_Display/n5522 ;
  wire \u2_Display/n5523 ;
  wire \u2_Display/n5524 ;
  wire \u2_Display/n5525 ;
  wire \u2_Display/n5526 ;
  wire \u2_Display/n5527 ;
  wire \u2_Display/n5528 ;
  wire \u2_Display/n5529 ;
  wire \u2_Display/n553 ;
  wire \u2_Display/n5530 ;
  wire \u2_Display/n5531 ;
  wire \u2_Display/n5532 ;
  wire \u2_Display/n5533 ;
  wire \u2_Display/n5534 ;
  wire \u2_Display/n5535 ;
  wire \u2_Display/n5536 ;
  wire \u2_Display/n5537 ;
  wire \u2_Display/n5538 ;
  wire \u2_Display/n5539 ;
  wire \u2_Display/n554 ;
  wire \u2_Display/n5542 ;
  wire \u2_Display/n5543 ;
  wire \u2_Display/n5544 ;
  wire \u2_Display/n5545 ;
  wire \u2_Display/n5546 ;
  wire \u2_Display/n5547 ;
  wire \u2_Display/n5548 ;
  wire \u2_Display/n5549 ;
  wire \u2_Display/n555 ;
  wire \u2_Display/n5550 ;
  wire \u2_Display/n5551 ;
  wire \u2_Display/n5552 ;
  wire \u2_Display/n5553 ;
  wire \u2_Display/n5554 ;
  wire \u2_Display/n5555 ;
  wire \u2_Display/n5556 ;
  wire \u2_Display/n5557 ;
  wire \u2_Display/n5558 ;
  wire \u2_Display/n5559 ;
  wire \u2_Display/n556 ;
  wire \u2_Display/n5560 ;
  wire \u2_Display/n5561 ;
  wire \u2_Display/n5562 ;
  wire \u2_Display/n5563 ;
  wire \u2_Display/n5564 ;
  wire \u2_Display/n5565 ;
  wire \u2_Display/n5566 ;
  wire \u2_Display/n5567 ;
  wire \u2_Display/n5568 ;
  wire \u2_Display/n5569 ;
  wire \u2_Display/n557 ;
  wire \u2_Display/n5570 ;
  wire \u2_Display/n5571 ;
  wire \u2_Display/n5572 ;
  wire \u2_Display/n5573 ;
  wire \u2_Display/n5574 ;
  wire \u2_Display/n5577 ;
  wire \u2_Display/n5578 ;
  wire \u2_Display/n5579 ;
  wire \u2_Display/n5580 ;
  wire \u2_Display/n5581 ;
  wire \u2_Display/n5582 ;
  wire \u2_Display/n5583 ;
  wire \u2_Display/n5584 ;
  wire \u2_Display/n5585 ;
  wire \u2_Display/n5586 ;
  wire \u2_Display/n5587 ;
  wire \u2_Display/n5588 ;
  wire \u2_Display/n5589 ;
  wire \u2_Display/n5590 ;
  wire \u2_Display/n5591 ;
  wire \u2_Display/n5592 ;
  wire \u2_Display/n5593 ;
  wire \u2_Display/n5594 ;
  wire \u2_Display/n5595 ;
  wire \u2_Display/n5596 ;
  wire \u2_Display/n5597 ;
  wire \u2_Display/n5598 ;
  wire \u2_Display/n5599 ;
  wire \u2_Display/n560 ;
  wire \u2_Display/n5600 ;
  wire \u2_Display/n5601 ;
  wire \u2_Display/n5602 ;
  wire \u2_Display/n5603 ;
  wire \u2_Display/n5604 ;
  wire \u2_Display/n5605 ;
  wire \u2_Display/n5606 ;
  wire \u2_Display/n5607 ;
  wire \u2_Display/n5608 ;
  wire \u2_Display/n5609 ;
  wire \u2_Display/n561 ;
  wire \u2_Display/n5612 ;
  wire \u2_Display/n5613 ;
  wire \u2_Display/n5614 ;
  wire \u2_Display/n5615 ;
  wire \u2_Display/n5616 ;
  wire \u2_Display/n5617 ;
  wire \u2_Display/n5618 ;
  wire \u2_Display/n5619 ;
  wire \u2_Display/n562 ;
  wire \u2_Display/n5620 ;
  wire \u2_Display/n5621 ;
  wire \u2_Display/n5622 ;
  wire \u2_Display/n5623 ;
  wire \u2_Display/n5624 ;
  wire \u2_Display/n5625 ;
  wire \u2_Display/n5626 ;
  wire \u2_Display/n5627 ;
  wire \u2_Display/n5628 ;
  wire \u2_Display/n5629 ;
  wire \u2_Display/n563 ;
  wire \u2_Display/n5630 ;
  wire \u2_Display/n5631 ;
  wire \u2_Display/n5632 ;
  wire \u2_Display/n5633 ;
  wire \u2_Display/n5634 ;
  wire \u2_Display/n5635 ;
  wire \u2_Display/n5636 ;
  wire \u2_Display/n5637 ;
  wire \u2_Display/n5638 ;
  wire \u2_Display/n5639 ;
  wire \u2_Display/n564 ;
  wire \u2_Display/n5640 ;
  wire \u2_Display/n5641 ;
  wire \u2_Display/n5642 ;
  wire \u2_Display/n5643 ;
  wire \u2_Display/n5644 ;
  wire \u2_Display/n5647 ;
  wire \u2_Display/n5648 ;
  wire \u2_Display/n5649 ;
  wire \u2_Display/n565 ;
  wire \u2_Display/n5650 ;
  wire \u2_Display/n5651 ;
  wire \u2_Display/n5652 ;
  wire \u2_Display/n5653 ;
  wire \u2_Display/n5654 ;
  wire \u2_Display/n5655 ;
  wire \u2_Display/n5656 ;
  wire \u2_Display/n5657 ;
  wire \u2_Display/n5658 ;
  wire \u2_Display/n5659 ;
  wire \u2_Display/n566 ;
  wire \u2_Display/n5660 ;
  wire \u2_Display/n5661 ;
  wire \u2_Display/n5662 ;
  wire \u2_Display/n5663 ;
  wire \u2_Display/n5664 ;
  wire \u2_Display/n5665 ;
  wire \u2_Display/n5666 ;
  wire \u2_Display/n5667 ;
  wire \u2_Display/n5668 ;
  wire \u2_Display/n5669 ;
  wire \u2_Display/n567 ;
  wire \u2_Display/n5670 ;
  wire \u2_Display/n5671 ;
  wire \u2_Display/n5672 ;
  wire \u2_Display/n5673 ;
  wire \u2_Display/n5674 ;
  wire \u2_Display/n5675 ;
  wire \u2_Display/n5676 ;
  wire \u2_Display/n5677 ;
  wire \u2_Display/n5678 ;
  wire \u2_Display/n5679 ;
  wire \u2_Display/n568 ;
  wire \u2_Display/n569 ;
  wire \u2_Display/n570 ;
  wire \u2_Display/n571 ;
  wire \u2_Display/n572 ;
  wire \u2_Display/n573 ;
  wire \u2_Display/n574 ;
  wire \u2_Display/n575 ;
  wire \u2_Display/n576 ;
  wire \u2_Display/n577 ;
  wire \u2_Display/n578 ;
  wire \u2_Display/n579 ;
  wire \u2_Display/n580 ;
  wire \u2_Display/n581 ;
  wire \u2_Display/n582 ;
  wire \u2_Display/n583 ;
  wire \u2_Display/n584 ;
  wire \u2_Display/n585 ;
  wire \u2_Display/n586 ;
  wire \u2_Display/n587 ;
  wire \u2_Display/n588 ;
  wire \u2_Display/n589 ;
  wire \u2_Display/n590 ;
  wire \u2_Display/n591 ;
  wire \u2_Display/n592 ;
  wire \u2_Display/n595 ;
  wire \u2_Display/n596 ;
  wire \u2_Display/n597 ;
  wire \u2_Display/n598 ;
  wire \u2_Display/n599 ;
  wire \u2_Display/n600 ;
  wire \u2_Display/n601 ;
  wire \u2_Display/n602 ;
  wire \u2_Display/n603 ;
  wire \u2_Display/n604 ;
  wire \u2_Display/n605 ;
  wire \u2_Display/n606 ;
  wire \u2_Display/n607 ;
  wire \u2_Display/n6070 ;
  wire \u2_Display/n6071 ;
  wire \u2_Display/n6072 ;
  wire \u2_Display/n6073 ;
  wire \u2_Display/n6074 ;
  wire \u2_Display/n6075 ;
  wire \u2_Display/n6076 ;
  wire \u2_Display/n6077 ;
  wire \u2_Display/n6078 ;
  wire \u2_Display/n6079 ;
  wire \u2_Display/n608 ;
  wire \u2_Display/n6080 ;
  wire \u2_Display/n6081 ;
  wire \u2_Display/n6082 ;
  wire \u2_Display/n6083 ;
  wire \u2_Display/n6084 ;
  wire \u2_Display/n6085 ;
  wire \u2_Display/n6086 ;
  wire \u2_Display/n6087 ;
  wire \u2_Display/n6088 ;
  wire \u2_Display/n6089 ;
  wire \u2_Display/n609 ;
  wire \u2_Display/n6090 ;
  wire \u2_Display/n6091 ;
  wire \u2_Display/n6092 ;
  wire \u2_Display/n6093 ;
  wire \u2_Display/n6094 ;
  wire \u2_Display/n6095 ;
  wire \u2_Display/n6096 ;
  wire \u2_Display/n6097 ;
  wire \u2_Display/n6098 ;
  wire \u2_Display/n6099 ;
  wire \u2_Display/n610 ;
  wire \u2_Display/n6100 ;
  wire \u2_Display/n6101 ;
  wire \u2_Display/n6105 ;
  wire \u2_Display/n6106 ;
  wire \u2_Display/n6107 ;
  wire \u2_Display/n6108 ;
  wire \u2_Display/n6109 ;
  wire \u2_Display/n611 ;
  wire \u2_Display/n6110 ;
  wire \u2_Display/n6111 ;
  wire \u2_Display/n6112 ;
  wire \u2_Display/n6113 ;
  wire \u2_Display/n6114 ;
  wire \u2_Display/n6115 ;
  wire \u2_Display/n6116 ;
  wire \u2_Display/n6117 ;
  wire \u2_Display/n6118 ;
  wire \u2_Display/n6119 ;
  wire \u2_Display/n612 ;
  wire \u2_Display/n6120 ;
  wire \u2_Display/n6121 ;
  wire \u2_Display/n6122 ;
  wire \u2_Display/n6123 ;
  wire \u2_Display/n6124 ;
  wire \u2_Display/n6125 ;
  wire \u2_Display/n6126 ;
  wire \u2_Display/n6127 ;
  wire \u2_Display/n6128 ;
  wire \u2_Display/n6129 ;
  wire \u2_Display/n613 ;
  wire \u2_Display/n6130 ;
  wire \u2_Display/n6131 ;
  wire \u2_Display/n6132 ;
  wire \u2_Display/n6133 ;
  wire \u2_Display/n6134 ;
  wire \u2_Display/n6135 ;
  wire \u2_Display/n6136 ;
  wire \u2_Display/n614 ;
  wire \u2_Display/n6140 ;
  wire \u2_Display/n6141 ;
  wire \u2_Display/n6142 ;
  wire \u2_Display/n6143 ;
  wire \u2_Display/n6144 ;
  wire \u2_Display/n6145 ;
  wire \u2_Display/n6146 ;
  wire \u2_Display/n6147 ;
  wire \u2_Display/n6148 ;
  wire \u2_Display/n6149 ;
  wire \u2_Display/n615 ;
  wire \u2_Display/n6150 ;
  wire \u2_Display/n6151 ;
  wire \u2_Display/n6152 ;
  wire \u2_Display/n6153 ;
  wire \u2_Display/n6154 ;
  wire \u2_Display/n6155 ;
  wire \u2_Display/n6156 ;
  wire \u2_Display/n6157 ;
  wire \u2_Display/n6158 ;
  wire \u2_Display/n6159 ;
  wire \u2_Display/n616 ;
  wire \u2_Display/n6160 ;
  wire \u2_Display/n6161 ;
  wire \u2_Display/n6162 ;
  wire \u2_Display/n6163 ;
  wire \u2_Display/n6164 ;
  wire \u2_Display/n6165 ;
  wire \u2_Display/n6166 ;
  wire \u2_Display/n6167 ;
  wire \u2_Display/n6168 ;
  wire \u2_Display/n6169 ;
  wire \u2_Display/n617 ;
  wire \u2_Display/n6170 ;
  wire \u2_Display/n6171 ;
  wire \u2_Display/n6175 ;
  wire \u2_Display/n6176 ;
  wire \u2_Display/n6177 ;
  wire \u2_Display/n6178 ;
  wire \u2_Display/n6179 ;
  wire \u2_Display/n618 ;
  wire \u2_Display/n6180 ;
  wire \u2_Display/n6181 ;
  wire \u2_Display/n6182 ;
  wire \u2_Display/n6183 ;
  wire \u2_Display/n6184 ;
  wire \u2_Display/n6185 ;
  wire \u2_Display/n6186 ;
  wire \u2_Display/n6187 ;
  wire \u2_Display/n6188 ;
  wire \u2_Display/n6189 ;
  wire \u2_Display/n619 ;
  wire \u2_Display/n6190 ;
  wire \u2_Display/n6191 ;
  wire \u2_Display/n6192 ;
  wire \u2_Display/n6193 ;
  wire \u2_Display/n6194 ;
  wire \u2_Display/n6195 ;
  wire \u2_Display/n6196 ;
  wire \u2_Display/n6197 ;
  wire \u2_Display/n6198 ;
  wire \u2_Display/n6199 ;
  wire \u2_Display/n620 ;
  wire \u2_Display/n6200 ;
  wire \u2_Display/n6201 ;
  wire \u2_Display/n6202 ;
  wire \u2_Display/n6203 ;
  wire \u2_Display/n6204 ;
  wire \u2_Display/n6205 ;
  wire \u2_Display/n6206 ;
  wire \u2_Display/n621 ;
  wire \u2_Display/n6210 ;
  wire \u2_Display/n6211 ;
  wire \u2_Display/n6212 ;
  wire \u2_Display/n6213 ;
  wire \u2_Display/n6214 ;
  wire \u2_Display/n6215 ;
  wire \u2_Display/n6216 ;
  wire \u2_Display/n6217 ;
  wire \u2_Display/n6218 ;
  wire \u2_Display/n6219 ;
  wire \u2_Display/n622 ;
  wire \u2_Display/n6220 ;
  wire \u2_Display/n6221 ;
  wire \u2_Display/n6222 ;
  wire \u2_Display/n6223 ;
  wire \u2_Display/n6224 ;
  wire \u2_Display/n6225 ;
  wire \u2_Display/n6226 ;
  wire \u2_Display/n6227 ;
  wire \u2_Display/n6228 ;
  wire \u2_Display/n6229 ;
  wire \u2_Display/n623 ;
  wire \u2_Display/n6230 ;
  wire \u2_Display/n6231 ;
  wire \u2_Display/n6232 ;
  wire \u2_Display/n6233 ;
  wire \u2_Display/n6234 ;
  wire \u2_Display/n6235 ;
  wire \u2_Display/n6236 ;
  wire \u2_Display/n6237 ;
  wire \u2_Display/n6238 ;
  wire \u2_Display/n6239 ;
  wire \u2_Display/n624 ;
  wire \u2_Display/n6240 ;
  wire \u2_Display/n6241 ;
  wire \u2_Display/n6245 ;
  wire \u2_Display/n6246 ;
  wire \u2_Display/n6247 ;
  wire \u2_Display/n6248 ;
  wire \u2_Display/n6249 ;
  wire \u2_Display/n625 ;
  wire \u2_Display/n6250 ;
  wire \u2_Display/n6251 ;
  wire \u2_Display/n6252 ;
  wire \u2_Display/n6253 ;
  wire \u2_Display/n6254 ;
  wire \u2_Display/n6255 ;
  wire \u2_Display/n6256 ;
  wire \u2_Display/n6257 ;
  wire \u2_Display/n6258 ;
  wire \u2_Display/n6259 ;
  wire \u2_Display/n626 ;
  wire \u2_Display/n6260 ;
  wire \u2_Display/n6261 ;
  wire \u2_Display/n6262 ;
  wire \u2_Display/n6263 ;
  wire \u2_Display/n6264 ;
  wire \u2_Display/n6265 ;
  wire \u2_Display/n6266 ;
  wire \u2_Display/n6267 ;
  wire \u2_Display/n6268 ;
  wire \u2_Display/n6269 ;
  wire \u2_Display/n627 ;
  wire \u2_Display/n6270 ;
  wire \u2_Display/n6271 ;
  wire \u2_Display/n6272 ;
  wire \u2_Display/n6273 ;
  wire \u2_Display/n6274 ;
  wire \u2_Display/n6275 ;
  wire \u2_Display/n6276 ;
  wire \u2_Display/n6280 ;
  wire \u2_Display/n6281 ;
  wire \u2_Display/n6282 ;
  wire \u2_Display/n6283 ;
  wire \u2_Display/n6284 ;
  wire \u2_Display/n6285 ;
  wire \u2_Display/n6286 ;
  wire \u2_Display/n6287 ;
  wire \u2_Display/n6288 ;
  wire \u2_Display/n6289 ;
  wire \u2_Display/n6290 ;
  wire \u2_Display/n6291 ;
  wire \u2_Display/n6292 ;
  wire \u2_Display/n6293 ;
  wire \u2_Display/n6294 ;
  wire \u2_Display/n6295 ;
  wire \u2_Display/n6296 ;
  wire \u2_Display/n6297 ;
  wire \u2_Display/n6298 ;
  wire \u2_Display/n6299 ;
  wire \u2_Display/n630 ;
  wire \u2_Display/n6300 ;
  wire \u2_Display/n6301 ;
  wire \u2_Display/n6302 ;
  wire \u2_Display/n6303 ;
  wire \u2_Display/n6304 ;
  wire \u2_Display/n6305 ;
  wire \u2_Display/n6306 ;
  wire \u2_Display/n6307 ;
  wire \u2_Display/n6308 ;
  wire \u2_Display/n6309 ;
  wire \u2_Display/n631 ;
  wire \u2_Display/n6310 ;
  wire \u2_Display/n6311 ;
  wire \u2_Display/n6315 ;
  wire \u2_Display/n6316 ;
  wire \u2_Display/n6317 ;
  wire \u2_Display/n6318 ;
  wire \u2_Display/n6319 ;
  wire \u2_Display/n632 ;
  wire \u2_Display/n6320 ;
  wire \u2_Display/n6321 ;
  wire \u2_Display/n6322 ;
  wire \u2_Display/n6323 ;
  wire \u2_Display/n6324 ;
  wire \u2_Display/n6325 ;
  wire \u2_Display/n6326 ;
  wire \u2_Display/n6327 ;
  wire \u2_Display/n6328 ;
  wire \u2_Display/n6329 ;
  wire \u2_Display/n633 ;
  wire \u2_Display/n6330 ;
  wire \u2_Display/n6331 ;
  wire \u2_Display/n6332 ;
  wire \u2_Display/n6333 ;
  wire \u2_Display/n6334 ;
  wire \u2_Display/n6335 ;
  wire \u2_Display/n6336 ;
  wire \u2_Display/n6337 ;
  wire \u2_Display/n6338 ;
  wire \u2_Display/n6339 ;
  wire \u2_Display/n634 ;
  wire \u2_Display/n6340 ;
  wire \u2_Display/n6341 ;
  wire \u2_Display/n6342 ;
  wire \u2_Display/n6343 ;
  wire \u2_Display/n6344 ;
  wire \u2_Display/n6345 ;
  wire \u2_Display/n6346 ;
  wire \u2_Display/n635 ;
  wire \u2_Display/n6350 ;
  wire \u2_Display/n6351 ;
  wire \u2_Display/n6352 ;
  wire \u2_Display/n6353 ;
  wire \u2_Display/n636 ;
  wire \u2_Display/n637 ;
  wire \u2_Display/n638 ;
  wire \u2_Display/n639 ;
  wire \u2_Display/n640 ;
  wire \u2_Display/n641 ;
  wire \u2_Display/n642 ;
  wire \u2_Display/n643 ;
  wire \u2_Display/n644 ;
  wire \u2_Display/n645 ;
  wire \u2_Display/n646 ;
  wire \u2_Display/n647 ;
  wire \u2_Display/n648 ;
  wire \u2_Display/n649 ;
  wire \u2_Display/n650 ;
  wire \u2_Display/n651 ;
  wire \u2_Display/n652 ;
  wire \u2_Display/n653 ;
  wire \u2_Display/n654 ;
  wire \u2_Display/n655 ;
  wire \u2_Display/n656 ;
  wire \u2_Display/n657 ;
  wire \u2_Display/n658 ;
  wire \u2_Display/n659 ;
  wire \u2_Display/n660 ;
  wire \u2_Display/n661 ;
  wire \u2_Display/n662 ;
  wire \u2_Display/n665 ;
  wire \u2_Display/n666 ;
  wire \u2_Display/n667 ;
  wire \u2_Display/n668 ;
  wire \u2_Display/n669 ;
  wire \u2_Display/n670 ;
  wire \u2_Display/n671 ;
  wire \u2_Display/n672 ;
  wire \u2_Display/n673 ;
  wire \u2_Display/n674 ;
  wire \u2_Display/n675 ;
  wire \u2_Display/n676 ;
  wire \u2_Display/n677 ;
  wire \u2_Display/n678 ;
  wire \u2_Display/n679 ;
  wire \u2_Display/n680 ;
  wire \u2_Display/n681 ;
  wire \u2_Display/n682 ;
  wire \u2_Display/n683 ;
  wire \u2_Display/n684 ;
  wire \u2_Display/n685 ;
  wire \u2_Display/n686 ;
  wire \u2_Display/n687 ;
  wire \u2_Display/n688 ;
  wire \u2_Display/n689 ;
  wire \u2_Display/n690 ;
  wire \u2_Display/n691 ;
  wire \u2_Display/n692 ;
  wire \u2_Display/n693 ;
  wire \u2_Display/n694 ;
  wire \u2_Display/n695 ;
  wire \u2_Display/n696 ;
  wire \u2_Display/n697 ;
  wire \u2_Display/n700 ;
  wire \u2_Display/n701 ;
  wire \u2_Display/n702 ;
  wire \u2_Display/n703 ;
  wire \u2_Display/n704 ;
  wire \u2_Display/n705 ;
  wire \u2_Display/n706 ;
  wire \u2_Display/n707 ;
  wire \u2_Display/n708 ;
  wire \u2_Display/n709 ;
  wire \u2_Display/n710 ;
  wire \u2_Display/n711 ;
  wire \u2_Display/n712 ;
  wire \u2_Display/n713 ;
  wire \u2_Display/n714 ;
  wire \u2_Display/n715 ;
  wire \u2_Display/n716 ;
  wire \u2_Display/n717 ;
  wire \u2_Display/n718 ;
  wire \u2_Display/n719 ;
  wire \u2_Display/n720 ;
  wire \u2_Display/n721 ;
  wire \u2_Display/n722 ;
  wire \u2_Display/n723 ;
  wire \u2_Display/n724 ;
  wire \u2_Display/n725 ;
  wire \u2_Display/n726 ;
  wire \u2_Display/n727 ;
  wire \u2_Display/n728 ;
  wire \u2_Display/n729 ;
  wire \u2_Display/n730 ;
  wire \u2_Display/n731 ;
  wire \u2_Display/n732 ;
  wire \u2_Display/n735 ;
  wire \u2_Display/n736 ;
  wire \u2_Display/n737 ;
  wire \u2_Display/n738 ;
  wire \u2_Display/n739 ;
  wire \u2_Display/n740 ;
  wire \u2_Display/n741 ;
  wire \u2_Display/n742 ;
  wire \u2_Display/n743 ;
  wire \u2_Display/n744 ;
  wire \u2_Display/n745 ;
  wire \u2_Display/n746 ;
  wire \u2_Display/n747 ;
  wire \u2_Display/n748 ;
  wire \u2_Display/n749 ;
  wire \u2_Display/n750 ;
  wire \u2_Display/n751 ;
  wire \u2_Display/n752 ;
  wire \u2_Display/n753 ;
  wire \u2_Display/n754 ;
  wire \u2_Display/n755 ;
  wire \u2_Display/n756 ;
  wire \u2_Display/n757 ;
  wire \u2_Display/n758 ;
  wire \u2_Display/n759 ;
  wire \u2_Display/n760 ;
  wire \u2_Display/n761 ;
  wire \u2_Display/n762 ;
  wire \u2_Display/n763 ;
  wire \u2_Display/n764 ;
  wire \u2_Display/n765 ;
  wire \u2_Display/n766 ;
  wire \u2_Display/n767 ;
  wire \u2_Display/n770 ;
  wire \u2_Display/n771 ;
  wire \u2_Display/n772 ;
  wire \u2_Display/n773 ;
  wire \u2_Display/n774 ;
  wire \u2_Display/n775 ;
  wire \u2_Display/n776 ;
  wire \u2_Display/n777 ;
  wire \u2_Display/n778 ;
  wire \u2_Display/n779 ;
  wire \u2_Display/n780 ;
  wire \u2_Display/n781 ;
  wire \u2_Display/n782 ;
  wire \u2_Display/n783 ;
  wire \u2_Display/n784 ;
  wire \u2_Display/n785 ;
  wire \u2_Display/n786 ;
  wire \u2_Display/n787 ;
  wire \u2_Display/n788 ;
  wire \u2_Display/n789 ;
  wire \u2_Display/n790 ;
  wire \u2_Display/n791 ;
  wire \u2_Display/n792 ;
  wire \u2_Display/n793 ;
  wire \u2_Display/n794 ;
  wire \u2_Display/n795 ;
  wire \u2_Display/n796 ;
  wire \u2_Display/n797 ;
  wire \u2_Display/n798 ;
  wire \u2_Display/n799 ;
  wire \u2_Display/n800 ;
  wire \u2_Display/n801 ;
  wire \u2_Display/n802 ;
  wire \u2_Display/n805 ;
  wire \u2_Display/n806 ;
  wire \u2_Display/n807 ;
  wire \u2_Display/n808 ;
  wire \u2_Display/n809 ;
  wire \u2_Display/n810 ;
  wire \u2_Display/n811 ;
  wire \u2_Display/n812 ;
  wire \u2_Display/n813 ;
  wire \u2_Display/n814 ;
  wire \u2_Display/n815 ;
  wire \u2_Display/n816 ;
  wire \u2_Display/n817 ;
  wire \u2_Display/n818 ;
  wire \u2_Display/n819 ;
  wire \u2_Display/n820 ;
  wire \u2_Display/n821 ;
  wire \u2_Display/n822 ;
  wire \u2_Display/n823 ;
  wire \u2_Display/n824 ;
  wire \u2_Display/n825 ;
  wire \u2_Display/n826 ;
  wire \u2_Display/n827 ;
  wire \u2_Display/n828 ;
  wire \u2_Display/n829 ;
  wire \u2_Display/n830 ;
  wire \u2_Display/n831 ;
  wire \u2_Display/n832 ;
  wire \u2_Display/n833 ;
  wire \u2_Display/n834 ;
  wire \u2_Display/n835 ;
  wire \u2_Display/n836 ;
  wire \u2_Display/n837 ;
  wire \u2_Display/n840 ;
  wire \u2_Display/n841 ;
  wire \u2_Display/n842 ;
  wire \u2_Display/n843 ;
  wire \u2_Display/n844 ;
  wire \u2_Display/n845 ;
  wire \u2_Display/n846 ;
  wire \u2_Display/n847 ;
  wire \u2_Display/n848 ;
  wire \u2_Display/n849 ;
  wire \u2_Display/n850 ;
  wire \u2_Display/n851 ;
  wire \u2_Display/n852 ;
  wire \u2_Display/n853 ;
  wire \u2_Display/n854 ;
  wire \u2_Display/n855 ;
  wire \u2_Display/n856 ;
  wire \u2_Display/n857 ;
  wire \u2_Display/n858 ;
  wire \u2_Display/n859 ;
  wire \u2_Display/n860 ;
  wire \u2_Display/n861 ;
  wire \u2_Display/n862 ;
  wire \u2_Display/n863 ;
  wire \u2_Display/n864 ;
  wire \u2_Display/n865 ;
  wire \u2_Display/n866 ;
  wire \u2_Display/n867 ;
  wire \u2_Display/n868 ;
  wire \u2_Display/n869 ;
  wire \u2_Display/n870 ;
  wire \u2_Display/n871 ;
  wire \u2_Display/n872 ;
  wire \u2_Display/n875 ;
  wire \u2_Display/n876 ;
  wire \u2_Display/n877 ;
  wire \u2_Display/n878 ;
  wire \u2_Display/n879 ;
  wire \u2_Display/n880 ;
  wire \u2_Display/n881 ;
  wire \u2_Display/n882 ;
  wire \u2_Display/n883 ;
  wire \u2_Display/n884 ;
  wire \u2_Display/n885 ;
  wire \u2_Display/n886 ;
  wire \u2_Display/n887 ;
  wire \u2_Display/n888 ;
  wire \u2_Display/n889 ;
  wire \u2_Display/n890 ;
  wire \u2_Display/n891 ;
  wire \u2_Display/n892 ;
  wire \u2_Display/n893 ;
  wire \u2_Display/n894 ;
  wire \u2_Display/n895 ;
  wire \u2_Display/n896 ;
  wire \u2_Display/n897 ;
  wire \u2_Display/n898 ;
  wire \u2_Display/n899 ;
  wire \u2_Display/n900 ;
  wire \u2_Display/n901 ;
  wire \u2_Display/n902 ;
  wire \u2_Display/n903 ;
  wire \u2_Display/n904 ;
  wire \u2_Display/n905 ;
  wire \u2_Display/n906 ;
  wire \u2_Display/n907 ;
  wire \u2_Display/n910 ;
  wire \u2_Display/n911 ;
  wire \u2_Display/n912 ;
  wire \u2_Display/n913 ;
  wire \u2_Display/n914 ;
  wire \u2_Display/n915 ;
  wire \u2_Display/n916 ;
  wire \u2_Display/n917 ;
  wire \u2_Display/n918 ;
  wire \u2_Display/n919 ;
  wire \u2_Display/n920 ;
  wire \u2_Display/n921 ;
  wire \u2_Display/n922 ;
  wire \u2_Display/n923 ;
  wire \u2_Display/n924 ;
  wire \u2_Display/n925 ;
  wire \u2_Display/n926 ;
  wire \u2_Display/n927 ;
  wire \u2_Display/n928 ;
  wire \u2_Display/n929 ;
  wire \u2_Display/n930 ;
  wire \u2_Display/n931 ;
  wire \u2_Display/n932 ;
  wire \u2_Display/n933 ;
  wire \u2_Display/n934 ;
  wire \u2_Display/n935 ;
  wire \u2_Display/n936 ;
  wire \u2_Display/n937 ;
  wire \u2_Display/n938 ;
  wire \u2_Display/n939 ;
  wire \u2_Display/n940 ;
  wire \u2_Display/n941 ;
  wire \u2_Display/n942 ;
  wire \u2_Display/n945 ;
  wire \u2_Display/n946 ;
  wire \u2_Display/n947 ;
  wire \u2_Display/n948 ;
  wire \u2_Display/n949 ;
  wire \u2_Display/n95 ;
  wire \u2_Display/n950 ;
  wire \u2_Display/n951 ;
  wire \u2_Display/n952 ;
  wire \u2_Display/n953 ;
  wire \u2_Display/n954 ;
  wire \u2_Display/n955 ;
  wire \u2_Display/n956 ;
  wire \u2_Display/n957 ;
  wire \u2_Display/n958 ;
  wire \u2_Display/n959 ;
  wire \u2_Display/n960 ;
  wire \u2_Display/n961 ;
  wire \u2_Display/n962 ;
  wire \u2_Display/n963 ;
  wire \u2_Display/n964 ;
  wire \u2_Display/n965 ;
  wire \u2_Display/n966 ;
  wire \u2_Display/n967 ;
  wire \u2_Display/n968 ;
  wire \u2_Display/n969 ;
  wire \u2_Display/n97 ;
  wire \u2_Display/n970 ;
  wire \u2_Display/n971 ;
  wire \u2_Display/n972 ;
  wire \u2_Display/n973 ;
  wire \u2_Display/n974 ;
  wire \u2_Display/n975 ;
  wire \u2_Display/n976 ;
  wire \u2_Display/n977 ;
  wire \u2_Display/n980 ;
  wire \u2_Display/n981 ;
  wire \u2_Display/n982 ;
  wire \u2_Display/n983 ;
  wire \u2_Display/n984 ;
  wire \u2_Display/n985 ;
  wire \u2_Display/n986 ;
  wire \u2_Display/n987 ;
  wire \u2_Display/n988 ;
  wire \u2_Display/n989 ;
  wire \u2_Display/n990 ;
  wire \u2_Display/n991 ;
  wire \u2_Display/n992 ;
  wire \u2_Display/n993 ;
  wire \u2_Display/n994 ;
  wire \u2_Display/n995 ;
  wire \u2_Display/n996 ;
  wire \u2_Display/n997 ;
  wire \u2_Display/n998 ;
  wire \u2_Display/n999 ;
  wire \u2_Display/sub0_2/c11 ;
  wire \u2_Display/sub0_2/c3 ;
  wire \u2_Display/sub0_2/c7 ;
  wire \u2_Display/sub1_2/c3 ;
  wire \u2_Display/sub1_2/c7 ;
  wire \u2_Display/sub2_2/c3 ;
  wire \u2_Display/sub2_2/c7 ;
  wire \u2_Display/sub3_2/c11 ;
  wire \u2_Display/sub3_2/c3 ;
  wire \u2_Display/sub3_2/c7 ;
  wire vga_clk_pad;  // source/rtl/VGA_Demo.v(9)
  wire vga_de_pad;  // source/rtl/VGA_Demo.v(13)
  wire vga_hs_pad;  // source/rtl/VGA_Demo.v(10)
  wire vga_vs_pad;  // source/rtl/VGA_Demo.v(11)

  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1000 (
    .a(\u2_Display/n3925 ),
    .b(\u2_Display/n3928 [0]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3960 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1001 (
    .a(\u2_Display/n3924 ),
    .b(\u2_Display/n3928 [1]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3959 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1002 (
    .a(\u2_Display/n3923 ),
    .b(\u2_Display/n3928 [2]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3958 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1003 (
    .a(\u2_Display/n3922 ),
    .b(\u2_Display/n3928 [3]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3957 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1004 (
    .a(\u2_Display/n3921 ),
    .b(\u2_Display/n3928 [4]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3956 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1005 (
    .a(\u2_Display/n3920 ),
    .b(\u2_Display/n3928 [5]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3955 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1006 (
    .a(\u2_Display/n3919 ),
    .b(\u2_Display/n3928 [6]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3954 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1007 (
    .a(\u2_Display/n3918 ),
    .b(\u2_Display/n3928 [7]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3953 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1008 (
    .a(\u2_Display/n3917 ),
    .b(\u2_Display/n3928 [8]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3952 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1009 (
    .a(\u2_Display/n3916 ),
    .b(\u2_Display/n3928 [9]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3951 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1010 (
    .a(\u2_Display/n3915 ),
    .b(\u2_Display/n3928 [10]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3950 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1011 (
    .a(\u2_Display/n3914 ),
    .b(\u2_Display/n3928 [11]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3949 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1012 (
    .a(\u2_Display/n3913 ),
    .b(\u2_Display/n3928 [12]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3948 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1013 (
    .a(\u2_Display/n3912 ),
    .b(\u2_Display/n3928 [13]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3947 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1014 (
    .a(\u2_Display/n3911 ),
    .b(\u2_Display/n3928 [14]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3946 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1015 (
    .a(\u2_Display/n3910 ),
    .b(\u2_Display/n3928 [15]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3945 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1016 (
    .a(\u2_Display/n3909 ),
    .b(\u2_Display/n3928 [16]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3944 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1017 (
    .a(\u2_Display/n3908 ),
    .b(\u2_Display/n3928 [17]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3943 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1018 (
    .a(\u2_Display/n3907 ),
    .b(\u2_Display/n3928 [18]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3942 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1019 (
    .a(\u2_Display/n3906 ),
    .b(\u2_Display/n3928 [19]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3941 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1020 (
    .a(\u2_Display/n3905 ),
    .b(\u2_Display/n3928 [20]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3940 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1021 (
    .a(\u2_Display/n3904 ),
    .b(\u2_Display/n3928 [21]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3939 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1022 (
    .a(\u2_Display/n3903 ),
    .b(\u2_Display/n3928 [22]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3938 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1023 (
    .a(\u2_Display/n3902 ),
    .b(\u2_Display/n3928 [23]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3937 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1024 (
    .a(\u2_Display/n3901 ),
    .b(\u2_Display/n3928 [24]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3936 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1025 (
    .a(\u2_Display/n3900 ),
    .b(\u2_Display/n3928 [25]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3935 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1026 (
    .a(\u2_Display/n3899 ),
    .b(\u2_Display/n3928 [26]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3934 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1027 (
    .a(\u2_Display/n3898 ),
    .b(\u2_Display/n3928 [27]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3933 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1028 (
    .a(\u2_Display/n3897 ),
    .b(\u2_Display/n3928 [28]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3932 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1029 (
    .a(\u2_Display/n3896 ),
    .b(\u2_Display/n3928 [29]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3931 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1030 (
    .a(\u2_Display/n3895 ),
    .b(\u2_Display/n3928 [30]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3930 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1031 (
    .a(\u2_Display/n3894 ),
    .b(\u2_Display/n3928 [31]),
    .c(\u2_Display/n3926 ),
    .o(\u2_Display/n3929 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1032 (
    .a(\u2_Display/n6206 ),
    .b(\u2_Display/n5051 [0]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6241 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1033 (
    .a(\u2_Display/n6205 ),
    .b(\u2_Display/n5051 [1]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6240 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1034 (
    .a(\u2_Display/n6204 ),
    .b(\u2_Display/n5051 [2]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6239 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1035 (
    .a(\u2_Display/n6203 ),
    .b(\u2_Display/n5051 [3]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6238 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1036 (
    .a(\u2_Display/n6202 ),
    .b(\u2_Display/n5051 [4]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6237 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1037 (
    .a(\u2_Display/n6201 ),
    .b(\u2_Display/n5051 [5]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6236 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1038 (
    .a(\u2_Display/n6200 ),
    .b(\u2_Display/n5051 [6]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6235 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1039 (
    .a(\u2_Display/n6199 ),
    .b(\u2_Display/n5051 [7]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6234 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1040 (
    .a(\u2_Display/n6198 ),
    .b(\u2_Display/n5051 [8]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6233 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1041 (
    .a(\u2_Display/n6197 ),
    .b(\u2_Display/n5051 [9]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6232 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1042 (
    .a(\u2_Display/n6196 ),
    .b(\u2_Display/n5051 [10]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6231 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1043 (
    .a(\u2_Display/n6195 ),
    .b(\u2_Display/n5051 [11]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6230 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1044 (
    .a(\u2_Display/n6194 ),
    .b(\u2_Display/n5051 [12]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6229 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1045 (
    .a(\u2_Display/n6193 ),
    .b(\u2_Display/n5051 [13]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6228 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1046 (
    .a(\u2_Display/n6192 ),
    .b(\u2_Display/n5051 [14]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6227 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1047 (
    .a(\u2_Display/n6191 ),
    .b(\u2_Display/n5051 [15]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6226 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1048 (
    .a(\u2_Display/n6190 ),
    .b(\u2_Display/n5051 [16]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6225 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1049 (
    .a(\u2_Display/n6189 ),
    .b(\u2_Display/n5051 [17]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6224 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1050 (
    .a(\u2_Display/n6188 ),
    .b(\u2_Display/n5051 [18]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6223 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1051 (
    .a(\u2_Display/n6187 ),
    .b(\u2_Display/n5051 [19]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6222 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1052 (
    .a(\u2_Display/n6186 ),
    .b(\u2_Display/n5051 [20]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6221 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1053 (
    .a(\u2_Display/n6185 ),
    .b(\u2_Display/n5051 [21]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6220 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1054 (
    .a(\u2_Display/n6184 ),
    .b(\u2_Display/n5051 [22]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6219 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1055 (
    .a(\u2_Display/n6183 ),
    .b(\u2_Display/n5051 [23]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6218 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1056 (
    .a(\u2_Display/n6182 ),
    .b(\u2_Display/n5051 [24]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6217 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1057 (
    .a(\u2_Display/n6181 ),
    .b(\u2_Display/n5051 [25]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6216 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1058 (
    .a(\u2_Display/n6180 ),
    .b(\u2_Display/n5051 [26]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6215 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1059 (
    .a(\u2_Display/n6179 ),
    .b(\u2_Display/n5051 [27]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6214 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1060 (
    .a(\u2_Display/n6178 ),
    .b(\u2_Display/n5051 [28]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6213 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1061 (
    .a(\u2_Display/n6177 ),
    .b(\u2_Display/n5051 [29]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6212 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1062 (
    .a(\u2_Display/n6176 ),
    .b(\u2_Display/n5051 [30]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6211 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1063 (
    .a(\u2_Display/n6175 ),
    .b(\u2_Display/n5051 [31]),
    .c(\u2_Display/n5049 ),
    .o(\u2_Display/n6210 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1064 (
    .a(\u2_Display/n556 ),
    .b(\u2_Display/n559 [0]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n591 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1065 (
    .a(\u2_Display/n555 ),
    .b(\u2_Display/n559 [1]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n590 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1066 (
    .a(\u2_Display/n554 ),
    .b(\u2_Display/n559 [2]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n589 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1067 (
    .a(\u2_Display/n553 ),
    .b(\u2_Display/n559 [3]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n588 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1068 (
    .a(\u2_Display/n552 ),
    .b(\u2_Display/n559 [4]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n587 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1069 (
    .a(\u2_Display/n551 ),
    .b(\u2_Display/n559 [5]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n586 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1070 (
    .a(\u2_Display/n550 ),
    .b(\u2_Display/n559 [6]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n585 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1071 (
    .a(\u2_Display/n549 ),
    .b(\u2_Display/n559 [7]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n584 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1072 (
    .a(\u2_Display/n548 ),
    .b(\u2_Display/n559 [8]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n583 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1073 (
    .a(\u2_Display/n547 ),
    .b(\u2_Display/n559 [9]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n582 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1074 (
    .a(\u2_Display/n546 ),
    .b(\u2_Display/n559 [10]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n581 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1075 (
    .a(\u2_Display/n545 ),
    .b(\u2_Display/n559 [11]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n580 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1076 (
    .a(\u2_Display/n544 ),
    .b(\u2_Display/n559 [12]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n579 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1077 (
    .a(\u2_Display/n543 ),
    .b(\u2_Display/n559 [13]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n578 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1078 (
    .a(\u2_Display/n542 ),
    .b(\u2_Display/n559 [14]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n577 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1079 (
    .a(\u2_Display/n541 ),
    .b(\u2_Display/n559 [15]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n576 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1080 (
    .a(\u2_Display/n540 ),
    .b(\u2_Display/n559 [16]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n575 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1081 (
    .a(\u2_Display/n539 ),
    .b(\u2_Display/n559 [17]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n574 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1082 (
    .a(\u2_Display/n538 ),
    .b(\u2_Display/n559 [18]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n573 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1083 (
    .a(\u2_Display/n537 ),
    .b(\u2_Display/n559 [19]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n572 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1084 (
    .a(\u2_Display/n536 ),
    .b(\u2_Display/n559 [20]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n571 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1085 (
    .a(\u2_Display/n535 ),
    .b(\u2_Display/n559 [21]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n570 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1086 (
    .a(\u2_Display/n534 ),
    .b(\u2_Display/n559 [22]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n569 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1087 (
    .a(\u2_Display/n533 ),
    .b(\u2_Display/n559 [23]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n568 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1088 (
    .a(\u2_Display/n532 ),
    .b(\u2_Display/n559 [24]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n567 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1089 (
    .a(\u2_Display/n531 ),
    .b(\u2_Display/n559 [25]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n566 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1090 (
    .a(\u2_Display/n530 ),
    .b(\u2_Display/n559 [26]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n565 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1091 (
    .a(\u2_Display/n529 ),
    .b(\u2_Display/n559 [27]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n564 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1092 (
    .a(\u2_Display/n528 ),
    .b(\u2_Display/n559 [28]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n563 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1093 (
    .a(\u2_Display/n527 ),
    .b(\u2_Display/n559 [29]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n562 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1094 (
    .a(\u2_Display/n526 ),
    .b(\u2_Display/n559 [30]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n561 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1095 (
    .a(\u2_Display/n525 ),
    .b(\u2_Display/n559 [31]),
    .c(\u2_Display/n557 ),
    .o(\u2_Display/n560 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1096 (
    .a(\u2_Display/n1679 ),
    .b(\u2_Display/n1682 [0]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1714 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1097 (
    .a(\u2_Display/n1678 ),
    .b(\u2_Display/n1682 [1]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1713 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1098 (
    .a(\u2_Display/n1677 ),
    .b(\u2_Display/n1682 [2]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1712 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1099 (
    .a(\u2_Display/n1676 ),
    .b(\u2_Display/n1682 [3]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1711 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1100 (
    .a(\u2_Display/n1675 ),
    .b(\u2_Display/n1682 [4]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1710 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1101 (
    .a(\u2_Display/n1674 ),
    .b(\u2_Display/n1682 [5]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1709 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1102 (
    .a(\u2_Display/n1673 ),
    .b(\u2_Display/n1682 [6]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1708 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1103 (
    .a(\u2_Display/n1672 ),
    .b(\u2_Display/n1682 [7]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1707 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1104 (
    .a(\u2_Display/n1671 ),
    .b(\u2_Display/n1682 [8]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1706 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1105 (
    .a(\u2_Display/n1670 ),
    .b(\u2_Display/n1682 [9]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1705 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1106 (
    .a(\u2_Display/n1669 ),
    .b(\u2_Display/n1682 [10]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1704 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1107 (
    .a(\u2_Display/n1668 ),
    .b(\u2_Display/n1682 [11]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1703 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1108 (
    .a(\u2_Display/n1667 ),
    .b(\u2_Display/n1682 [12]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1702 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1109 (
    .a(\u2_Display/n1666 ),
    .b(\u2_Display/n1682 [13]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1701 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1110 (
    .a(\u2_Display/n1665 ),
    .b(\u2_Display/n1682 [14]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1700 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1111 (
    .a(\u2_Display/n1664 ),
    .b(\u2_Display/n1682 [15]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1699 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1112 (
    .a(\u2_Display/n1663 ),
    .b(\u2_Display/n1682 [16]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1698 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1113 (
    .a(\u2_Display/n1662 ),
    .b(\u2_Display/n1682 [17]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1697 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1114 (
    .a(\u2_Display/n1661 ),
    .b(\u2_Display/n1682 [18]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1696 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1115 (
    .a(\u2_Display/n1660 ),
    .b(\u2_Display/n1682 [19]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1695 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1116 (
    .a(\u2_Display/n1659 ),
    .b(\u2_Display/n1682 [20]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1694 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1117 (
    .a(\u2_Display/n1658 ),
    .b(\u2_Display/n1682 [21]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1693 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1118 (
    .a(\u2_Display/n1657 ),
    .b(\u2_Display/n1682 [22]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1692 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1119 (
    .a(\u2_Display/n1656 ),
    .b(\u2_Display/n1682 [23]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1691 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1120 (
    .a(\u2_Display/n1655 ),
    .b(\u2_Display/n1682 [24]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1690 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1121 (
    .a(\u2_Display/n1654 ),
    .b(\u2_Display/n1682 [25]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1689 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1122 (
    .a(\u2_Display/n1653 ),
    .b(\u2_Display/n1682 [26]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1688 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1123 (
    .a(\u2_Display/n1652 ),
    .b(\u2_Display/n1682 [27]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1687 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1124 (
    .a(\u2_Display/n1651 ),
    .b(\u2_Display/n1682 [28]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1686 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1125 (
    .a(\u2_Display/n1650 ),
    .b(\u2_Display/n1682 [29]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1685 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1126 (
    .a(\u2_Display/n1649 ),
    .b(\u2_Display/n1682 [30]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1684 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1127 (
    .a(\u2_Display/n1648 ),
    .b(\u2_Display/n1682 [31]),
    .c(\u2_Display/n1680 ),
    .o(\u2_Display/n1683 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1128 (
    .a(\u2_Display/n2802 ),
    .b(\u2_Display/n2805 [0]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2837 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1129 (
    .a(\u2_Display/n2801 ),
    .b(\u2_Display/n2805 [1]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2836 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1130 (
    .a(\u2_Display/n2800 ),
    .b(\u2_Display/n2805 [2]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2835 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1131 (
    .a(\u2_Display/n2799 ),
    .b(\u2_Display/n2805 [3]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2834 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1132 (
    .a(\u2_Display/n2798 ),
    .b(\u2_Display/n2805 [4]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2833 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1133 (
    .a(\u2_Display/n2797 ),
    .b(\u2_Display/n2805 [5]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2832 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1134 (
    .a(\u2_Display/n2796 ),
    .b(\u2_Display/n2805 [6]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2831 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1135 (
    .a(\u2_Display/n2795 ),
    .b(\u2_Display/n2805 [7]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2830 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1136 (
    .a(\u2_Display/n2794 ),
    .b(\u2_Display/n2805 [8]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2829 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1137 (
    .a(\u2_Display/n2793 ),
    .b(\u2_Display/n2805 [9]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2828 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1138 (
    .a(\u2_Display/n2792 ),
    .b(\u2_Display/n2805 [10]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2827 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1139 (
    .a(\u2_Display/n2791 ),
    .b(\u2_Display/n2805 [11]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2826 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1140 (
    .a(\u2_Display/n2790 ),
    .b(\u2_Display/n2805 [12]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2825 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1141 (
    .a(\u2_Display/n2789 ),
    .b(\u2_Display/n2805 [13]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2824 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1142 (
    .a(\u2_Display/n2788 ),
    .b(\u2_Display/n2805 [14]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2823 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1143 (
    .a(\u2_Display/n2787 ),
    .b(\u2_Display/n2805 [15]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2822 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1144 (
    .a(\u2_Display/n2786 ),
    .b(\u2_Display/n2805 [16]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2821 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1145 (
    .a(\u2_Display/n2785 ),
    .b(\u2_Display/n2805 [17]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2820 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1146 (
    .a(\u2_Display/n2784 ),
    .b(\u2_Display/n2805 [18]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2819 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1147 (
    .a(\u2_Display/n2783 ),
    .b(\u2_Display/n2805 [19]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2818 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1148 (
    .a(\u2_Display/n2782 ),
    .b(\u2_Display/n2805 [20]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2817 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1149 (
    .a(\u2_Display/n2781 ),
    .b(\u2_Display/n2805 [21]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2816 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1150 (
    .a(\u2_Display/n2780 ),
    .b(\u2_Display/n2805 [22]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2815 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1151 (
    .a(\u2_Display/n2779 ),
    .b(\u2_Display/n2805 [23]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2814 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1152 (
    .a(\u2_Display/n2778 ),
    .b(\u2_Display/n2805 [24]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2813 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1153 (
    .a(\u2_Display/n2777 ),
    .b(\u2_Display/n2805 [25]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2812 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1154 (
    .a(\u2_Display/n2776 ),
    .b(\u2_Display/n2805 [26]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2811 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1155 (
    .a(\u2_Display/n2775 ),
    .b(\u2_Display/n2805 [27]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2810 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1156 (
    .a(\u2_Display/n2774 ),
    .b(\u2_Display/n2805 [28]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2809 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1157 (
    .a(\u2_Display/n2773 ),
    .b(\u2_Display/n2805 [29]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2808 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1158 (
    .a(\u2_Display/n2772 ),
    .b(\u2_Display/n2805 [30]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2807 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1159 (
    .a(\u2_Display/n2771 ),
    .b(\u2_Display/n2805 [31]),
    .c(\u2_Display/n2803 ),
    .o(\u2_Display/n2806 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1160 (
    .a(on_off_pad[3]),
    .b(on_off_pad[2]),
    .o(\u2_Display/mux11_b0_sel_is_0_o ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1161 (
    .a(on_off_pad[4]),
    .b(on_off_pad[3]),
    .o(\u2_Display/mux5_b0_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1162 (
    .a(\u2_Display/n141 ),
    .b(\u2_Display/n144 ),
    .c(\u2_Display/n136 ),
    .d(\u2_Display/n138 ),
    .o(\u2_Display/n145 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1163 (
    .a(on_off_pad[1]),
    .b(on_off_pad[0]),
    .o(\u2_Display/mux19_b0_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1164 (
    .a(\u2_Display/n44 ),
    .b(\u2_Display/n45 ),
    .c(\u2_Display/n48 ),
    .d(\u2_Display/n50 ),
    .o(\u2_Display/n51 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1165 (
    .a(\u2_Display/n95 ),
    .b(\u2_Display/n97 ),
    .c(\u2_Display/n100 ),
    .d(\u2_Display/n103 ),
    .o(\u2_Display/n104 ));
  AL_MAP_LUT5 #(
    .EQN("((A*~(~D*C))*~(B)*~(E)+(A*~(~D*C))*B*~(E)+~((A*~(~D*C)))*B*E+(A*~(~D*C))*B*E)"),
    .INIT(32'hccccaa0a))
    _al_u1166 (
    .a(\u2_Display/n145 ),
    .b(\u2_Display/n104 ),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(on_off_pad[1]),
    .o(\u2_Display/n236 [0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u1167 (
    .a(\u2_Display/n236 [0]),
    .b(\u2_Display/n51 ),
    .c(on_off_pad[0]),
    .o(\u2_Display/n240 [0]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1168 (
    .a(\u2_Display/mux11_b0_sel_is_0_o ),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(on_off_pad[4]),
    .o(_al_u1168_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1169 (
    .a(_al_u1168_o),
    .b(rst_n_pad),
    .o(\u2_Display/mux21_b0_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1170 (
    .a(\u1_Driver/vcnt [6]),
    .b(\u1_Driver/vcnt [7]),
    .c(\u1_Driver/vcnt [8]),
    .d(\u1_Driver/vcnt [9]),
    .o(_al_u1170_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    _al_u1171 (
    .a(_al_u1170_o),
    .b(\u1_Driver/vcnt [0]),
    .c(\u1_Driver/vcnt [10]),
    .d(\u1_Driver/vcnt [2]),
    .e(\u1_Driver/vcnt [4]),
    .o(_al_u1171_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*A)"),
    .INIT(32'h02000000))
    _al_u1172 (
    .a(_al_u1171_o),
    .b(\u1_Driver/vcnt [1]),
    .c(\u1_Driver/vcnt [11]),
    .d(\u1_Driver/vcnt [3]),
    .e(\u1_Driver/vcnt [5]),
    .o(\u1_Driver/n6_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1173 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [9]),
    .o(\u1_Driver/n8 [9]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1174 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [8]),
    .o(\u1_Driver/n8 [8]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1175 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [7]),
    .o(\u1_Driver/n8 [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1176 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [6]),
    .o(\u1_Driver/n8 [6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1177 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [5]),
    .o(\u1_Driver/n8 [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1178 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [4]),
    .o(\u1_Driver/n8 [4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1179 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [3]),
    .o(\u1_Driver/n8 [3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1180 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [2]),
    .o(\u1_Driver/n8 [2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1181 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [11]),
    .o(\u1_Driver/n8 [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1182 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [10]),
    .o(\u1_Driver/n8 [10]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1183 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [1]),
    .o(\u1_Driver/n8 [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1184 (
    .a(\u1_Driver/n6_lutinv ),
    .b(\u1_Driver/n7 [0]),
    .o(\u1_Driver/n8 [0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1185 (
    .a(\u2_Display/n3960 ),
    .b(\u2_Display/n3963 [0]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3995 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1186 (
    .a(\u2_Display/n3959 ),
    .b(\u2_Display/n3963 [1]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3994 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1187 (
    .a(\u2_Display/n3958 ),
    .b(\u2_Display/n3963 [2]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3993 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1188 (
    .a(\u2_Display/n3957 ),
    .b(\u2_Display/n3963 [3]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3992 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1189 (
    .a(\u2_Display/n3956 ),
    .b(\u2_Display/n3963 [4]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3991 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1190 (
    .a(\u2_Display/n3955 ),
    .b(\u2_Display/n3963 [5]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3990 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1191 (
    .a(\u2_Display/n3954 ),
    .b(\u2_Display/n3963 [6]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3989 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1192 (
    .a(\u2_Display/n3953 ),
    .b(\u2_Display/n3963 [7]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3988 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1193 (
    .a(\u2_Display/n3952 ),
    .b(\u2_Display/n3963 [8]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3987 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1194 (
    .a(\u2_Display/n3951 ),
    .b(\u2_Display/n3963 [9]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3986 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1195 (
    .a(\u2_Display/n3950 ),
    .b(\u2_Display/n3963 [10]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3985 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1196 (
    .a(\u2_Display/n3949 ),
    .b(\u2_Display/n3963 [11]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3984 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1197 (
    .a(\u2_Display/n3948 ),
    .b(\u2_Display/n3963 [12]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3983 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1198 (
    .a(\u2_Display/n3947 ),
    .b(\u2_Display/n3963 [13]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3982 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1199 (
    .a(\u2_Display/n3946 ),
    .b(\u2_Display/n3963 [14]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3981 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1200 (
    .a(\u2_Display/n3945 ),
    .b(\u2_Display/n3963 [15]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3980 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1201 (
    .a(\u2_Display/n3944 ),
    .b(\u2_Display/n3963 [16]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3979 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1202 (
    .a(\u2_Display/n3943 ),
    .b(\u2_Display/n3963 [17]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3978 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1203 (
    .a(\u2_Display/n3942 ),
    .b(\u2_Display/n3963 [18]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3977 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1204 (
    .a(\u2_Display/n3941 ),
    .b(\u2_Display/n3963 [19]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3976 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1205 (
    .a(\u2_Display/n3940 ),
    .b(\u2_Display/n3963 [20]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3975 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1206 (
    .a(\u2_Display/n3939 ),
    .b(\u2_Display/n3963 [21]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3974 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1207 (
    .a(\u2_Display/n3938 ),
    .b(\u2_Display/n3963 [22]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3973 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1208 (
    .a(\u2_Display/n3937 ),
    .b(\u2_Display/n3963 [23]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3972 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1209 (
    .a(\u2_Display/n3936 ),
    .b(\u2_Display/n3963 [24]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3971 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1210 (
    .a(\u2_Display/n3935 ),
    .b(\u2_Display/n3963 [25]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3970 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1211 (
    .a(\u2_Display/n3934 ),
    .b(\u2_Display/n3963 [26]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3969 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1212 (
    .a(\u2_Display/n3933 ),
    .b(\u2_Display/n3963 [27]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3968 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1213 (
    .a(\u2_Display/n3932 ),
    .b(\u2_Display/n3963 [28]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3967 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1214 (
    .a(\u2_Display/n3931 ),
    .b(\u2_Display/n3963 [29]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3966 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1215 (
    .a(\u2_Display/n3930 ),
    .b(\u2_Display/n3963 [30]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3965 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1216 (
    .a(\u2_Display/n3929 ),
    .b(\u2_Display/n3963 [31]),
    .c(\u2_Display/n3961 ),
    .o(\u2_Display/n3964 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1217 (
    .a(\u2_Display/n6241 ),
    .b(\u2_Display/n5086 [0]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6276 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1218 (
    .a(\u2_Display/n6240 ),
    .b(\u2_Display/n5086 [1]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6275 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1219 (
    .a(\u2_Display/n6239 ),
    .b(\u2_Display/n5086 [2]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6274 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1220 (
    .a(\u2_Display/n6238 ),
    .b(\u2_Display/n5086 [3]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6273 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1221 (
    .a(\u2_Display/n6237 ),
    .b(\u2_Display/n5086 [4]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6272 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1222 (
    .a(\u2_Display/n6236 ),
    .b(\u2_Display/n5086 [5]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6271 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1223 (
    .a(\u2_Display/n6235 ),
    .b(\u2_Display/n5086 [6]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6270 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1224 (
    .a(\u2_Display/n6234 ),
    .b(\u2_Display/n5086 [7]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6269 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1225 (
    .a(\u2_Display/n6233 ),
    .b(\u2_Display/n5086 [8]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6268 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1226 (
    .a(\u2_Display/n6232 ),
    .b(\u2_Display/n5086 [9]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6267 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1227 (
    .a(\u2_Display/n6231 ),
    .b(\u2_Display/n5086 [10]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6266 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1228 (
    .a(\u2_Display/n6230 ),
    .b(\u2_Display/n5086 [11]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6265 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1229 (
    .a(\u2_Display/n6229 ),
    .b(\u2_Display/n5086 [12]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6264 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1230 (
    .a(\u2_Display/n6228 ),
    .b(\u2_Display/n5086 [13]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6263 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1231 (
    .a(\u2_Display/n6227 ),
    .b(\u2_Display/n5086 [14]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6262 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1232 (
    .a(\u2_Display/n6226 ),
    .b(\u2_Display/n5086 [15]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6261 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1233 (
    .a(\u2_Display/n6225 ),
    .b(\u2_Display/n5086 [16]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6260 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1234 (
    .a(\u2_Display/n6224 ),
    .b(\u2_Display/n5086 [17]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6259 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1235 (
    .a(\u2_Display/n6223 ),
    .b(\u2_Display/n5086 [18]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6258 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1236 (
    .a(\u2_Display/n6222 ),
    .b(\u2_Display/n5086 [19]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6257 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1237 (
    .a(\u2_Display/n6221 ),
    .b(\u2_Display/n5086 [20]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6256 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1238 (
    .a(\u2_Display/n6220 ),
    .b(\u2_Display/n5086 [21]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6255 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1239 (
    .a(\u2_Display/n6219 ),
    .b(\u2_Display/n5086 [22]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6254 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1240 (
    .a(\u2_Display/n6218 ),
    .b(\u2_Display/n5086 [23]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6253 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1241 (
    .a(\u2_Display/n6217 ),
    .b(\u2_Display/n5086 [24]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6252 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1242 (
    .a(\u2_Display/n6216 ),
    .b(\u2_Display/n5086 [25]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6251 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1243 (
    .a(\u2_Display/n6215 ),
    .b(\u2_Display/n5086 [26]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6250 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1244 (
    .a(\u2_Display/n6214 ),
    .b(\u2_Display/n5086 [27]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6249 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1245 (
    .a(\u2_Display/n6213 ),
    .b(\u2_Display/n5086 [28]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6248 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1246 (
    .a(\u2_Display/n6212 ),
    .b(\u2_Display/n5086 [29]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6247 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1247 (
    .a(\u2_Display/n6211 ),
    .b(\u2_Display/n5086 [30]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6246 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1248 (
    .a(\u2_Display/n6210 ),
    .b(\u2_Display/n5086 [31]),
    .c(\u2_Display/n5084 ),
    .o(\u2_Display/n6245 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1249 (
    .a(\u2_Display/n591 ),
    .b(\u2_Display/n594 [0]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n626 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1250 (
    .a(\u2_Display/n590 ),
    .b(\u2_Display/n594 [1]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n625 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1251 (
    .a(\u2_Display/n589 ),
    .b(\u2_Display/n594 [2]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n624 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1252 (
    .a(\u2_Display/n588 ),
    .b(\u2_Display/n594 [3]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n623 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1253 (
    .a(\u2_Display/n587 ),
    .b(\u2_Display/n594 [4]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n622 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1254 (
    .a(\u2_Display/n586 ),
    .b(\u2_Display/n594 [5]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n621 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1255 (
    .a(\u2_Display/n585 ),
    .b(\u2_Display/n594 [6]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n620 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1256 (
    .a(\u2_Display/n584 ),
    .b(\u2_Display/n594 [7]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n619 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1257 (
    .a(\u2_Display/n583 ),
    .b(\u2_Display/n594 [8]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n618 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1258 (
    .a(\u2_Display/n582 ),
    .b(\u2_Display/n594 [9]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n617 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1259 (
    .a(\u2_Display/n581 ),
    .b(\u2_Display/n594 [10]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n616 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1260 (
    .a(\u2_Display/n580 ),
    .b(\u2_Display/n594 [11]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n615 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1261 (
    .a(\u2_Display/n579 ),
    .b(\u2_Display/n594 [12]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n614 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1262 (
    .a(\u2_Display/n578 ),
    .b(\u2_Display/n594 [13]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n613 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1263 (
    .a(\u2_Display/n577 ),
    .b(\u2_Display/n594 [14]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n612 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1264 (
    .a(\u2_Display/n576 ),
    .b(\u2_Display/n594 [15]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n611 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1265 (
    .a(\u2_Display/n575 ),
    .b(\u2_Display/n594 [16]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n610 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1266 (
    .a(\u2_Display/n574 ),
    .b(\u2_Display/n594 [17]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n609 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1267 (
    .a(\u2_Display/n573 ),
    .b(\u2_Display/n594 [18]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n608 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1268 (
    .a(\u2_Display/n572 ),
    .b(\u2_Display/n594 [19]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n607 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1269 (
    .a(\u2_Display/n571 ),
    .b(\u2_Display/n594 [20]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n606 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1270 (
    .a(\u2_Display/n570 ),
    .b(\u2_Display/n594 [21]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n605 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1271 (
    .a(\u2_Display/n569 ),
    .b(\u2_Display/n594 [22]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n604 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1272 (
    .a(\u2_Display/n568 ),
    .b(\u2_Display/n594 [23]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n603 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1273 (
    .a(\u2_Display/n567 ),
    .b(\u2_Display/n594 [24]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n602 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1274 (
    .a(\u2_Display/n566 ),
    .b(\u2_Display/n594 [25]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n601 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1275 (
    .a(\u2_Display/n565 ),
    .b(\u2_Display/n594 [26]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n600 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1276 (
    .a(\u2_Display/n564 ),
    .b(\u2_Display/n594 [27]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n599 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1277 (
    .a(\u2_Display/n563 ),
    .b(\u2_Display/n594 [28]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n598 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1278 (
    .a(\u2_Display/n562 ),
    .b(\u2_Display/n594 [29]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n597 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1279 (
    .a(\u2_Display/n561 ),
    .b(\u2_Display/n594 [30]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n596 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1280 (
    .a(\u2_Display/n560 ),
    .b(\u2_Display/n594 [31]),
    .c(\u2_Display/n592 ),
    .o(\u2_Display/n595 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1281 (
    .a(\u2_Display/n1714 ),
    .b(\u2_Display/n1717 [0]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1749 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1282 (
    .a(\u2_Display/n1713 ),
    .b(\u2_Display/n1717 [1]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1748 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1283 (
    .a(\u2_Display/n1712 ),
    .b(\u2_Display/n1717 [2]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1747 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1284 (
    .a(\u2_Display/n1711 ),
    .b(\u2_Display/n1717 [3]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1746 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1285 (
    .a(\u2_Display/n1710 ),
    .b(\u2_Display/n1717 [4]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1745 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1286 (
    .a(\u2_Display/n1709 ),
    .b(\u2_Display/n1717 [5]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1744 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1287 (
    .a(\u2_Display/n1708 ),
    .b(\u2_Display/n1717 [6]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1743 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1288 (
    .a(\u2_Display/n1707 ),
    .b(\u2_Display/n1717 [7]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1742 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1289 (
    .a(\u2_Display/n1706 ),
    .b(\u2_Display/n1717 [8]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1741 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1290 (
    .a(\u2_Display/n1705 ),
    .b(\u2_Display/n1717 [9]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1740 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1291 (
    .a(\u2_Display/n1704 ),
    .b(\u2_Display/n1717 [10]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1739 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1292 (
    .a(\u2_Display/n1703 ),
    .b(\u2_Display/n1717 [11]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1738 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1293 (
    .a(\u2_Display/n1702 ),
    .b(\u2_Display/n1717 [12]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1737 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1294 (
    .a(\u2_Display/n1701 ),
    .b(\u2_Display/n1717 [13]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1736 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1295 (
    .a(\u2_Display/n1700 ),
    .b(\u2_Display/n1717 [14]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1735 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1296 (
    .a(\u2_Display/n1699 ),
    .b(\u2_Display/n1717 [15]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1734 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1297 (
    .a(\u2_Display/n1698 ),
    .b(\u2_Display/n1717 [16]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1733 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1298 (
    .a(\u2_Display/n1697 ),
    .b(\u2_Display/n1717 [17]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1732 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1299 (
    .a(\u2_Display/n1696 ),
    .b(\u2_Display/n1717 [18]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1731 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1300 (
    .a(\u2_Display/n1695 ),
    .b(\u2_Display/n1717 [19]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1730 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1301 (
    .a(\u2_Display/n1694 ),
    .b(\u2_Display/n1717 [20]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1729 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1302 (
    .a(\u2_Display/n1693 ),
    .b(\u2_Display/n1717 [21]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1728 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1303 (
    .a(\u2_Display/n1692 ),
    .b(\u2_Display/n1717 [22]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1727 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1304 (
    .a(\u2_Display/n1691 ),
    .b(\u2_Display/n1717 [23]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1726 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1305 (
    .a(\u2_Display/n1690 ),
    .b(\u2_Display/n1717 [24]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1725 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1306 (
    .a(\u2_Display/n1689 ),
    .b(\u2_Display/n1717 [25]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1724 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1307 (
    .a(\u2_Display/n1688 ),
    .b(\u2_Display/n1717 [26]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1723 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1308 (
    .a(\u2_Display/n1687 ),
    .b(\u2_Display/n1717 [27]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1722 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1309 (
    .a(\u2_Display/n1686 ),
    .b(\u2_Display/n1717 [28]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1721 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1310 (
    .a(\u2_Display/n1685 ),
    .b(\u2_Display/n1717 [29]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1720 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1311 (
    .a(\u2_Display/n1684 ),
    .b(\u2_Display/n1717 [30]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1719 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1312 (
    .a(\u2_Display/n1683 ),
    .b(\u2_Display/n1717 [31]),
    .c(\u2_Display/n1715 ),
    .o(\u2_Display/n1718 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1313 (
    .a(\u2_Display/n2837 ),
    .b(\u2_Display/n2840 [0]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2872 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1314 (
    .a(\u2_Display/n2836 ),
    .b(\u2_Display/n2840 [1]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2871 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1315 (
    .a(\u2_Display/n2835 ),
    .b(\u2_Display/n2840 [2]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2870 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1316 (
    .a(\u2_Display/n2834 ),
    .b(\u2_Display/n2840 [3]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2869 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1317 (
    .a(\u2_Display/n2833 ),
    .b(\u2_Display/n2840 [4]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2868 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1318 (
    .a(\u2_Display/n2832 ),
    .b(\u2_Display/n2840 [5]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2867 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1319 (
    .a(\u2_Display/n2831 ),
    .b(\u2_Display/n2840 [6]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2866 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1320 (
    .a(\u2_Display/n2830 ),
    .b(\u2_Display/n2840 [7]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2865 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1321 (
    .a(\u2_Display/n2829 ),
    .b(\u2_Display/n2840 [8]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2864 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1322 (
    .a(\u2_Display/n2828 ),
    .b(\u2_Display/n2840 [9]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2863 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1323 (
    .a(\u2_Display/n2827 ),
    .b(\u2_Display/n2840 [10]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2862 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1324 (
    .a(\u2_Display/n2826 ),
    .b(\u2_Display/n2840 [11]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2861 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1325 (
    .a(\u2_Display/n2825 ),
    .b(\u2_Display/n2840 [12]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2860 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1326 (
    .a(\u2_Display/n2824 ),
    .b(\u2_Display/n2840 [13]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2859 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1327 (
    .a(\u2_Display/n2823 ),
    .b(\u2_Display/n2840 [14]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2858 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1328 (
    .a(\u2_Display/n2822 ),
    .b(\u2_Display/n2840 [15]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2857 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1329 (
    .a(\u2_Display/n2821 ),
    .b(\u2_Display/n2840 [16]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2856 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1330 (
    .a(\u2_Display/n2820 ),
    .b(\u2_Display/n2840 [17]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2855 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1331 (
    .a(\u2_Display/n2819 ),
    .b(\u2_Display/n2840 [18]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2854 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1332 (
    .a(\u2_Display/n2818 ),
    .b(\u2_Display/n2840 [19]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2853 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1333 (
    .a(\u2_Display/n2817 ),
    .b(\u2_Display/n2840 [20]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2852 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1334 (
    .a(\u2_Display/n2816 ),
    .b(\u2_Display/n2840 [21]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2851 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1335 (
    .a(\u2_Display/n2815 ),
    .b(\u2_Display/n2840 [22]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2850 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1336 (
    .a(\u2_Display/n2814 ),
    .b(\u2_Display/n2840 [23]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2849 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1337 (
    .a(\u2_Display/n2813 ),
    .b(\u2_Display/n2840 [24]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2848 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1338 (
    .a(\u2_Display/n2812 ),
    .b(\u2_Display/n2840 [25]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2847 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1339 (
    .a(\u2_Display/n2811 ),
    .b(\u2_Display/n2840 [26]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2846 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1340 (
    .a(\u2_Display/n2810 ),
    .b(\u2_Display/n2840 [27]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2845 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1341 (
    .a(\u2_Display/n2809 ),
    .b(\u2_Display/n2840 [28]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2844 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1342 (
    .a(\u2_Display/n2808 ),
    .b(\u2_Display/n2840 [29]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2843 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1343 (
    .a(\u2_Display/n2807 ),
    .b(\u2_Display/n2840 [30]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2842 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1344 (
    .a(\u2_Display/n2806 ),
    .b(\u2_Display/n2840 [31]),
    .c(\u2_Display/n2838 ),
    .o(\u2_Display/n2841 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1345 (
    .a(\u2_Display/n [27]),
    .b(\u2_Display/n [28]),
    .c(\u2_Display/n [29]),
    .d(\u2_Display/n [3]),
    .o(_al_u1345_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1346 (
    .a(\u2_Display/n [23]),
    .b(\u2_Display/n [24]),
    .c(\u2_Display/n [25]),
    .d(\u2_Display/n [26]),
    .o(_al_u1346_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u1347 (
    .a(\u2_Display/n [30]),
    .b(\u2_Display/n [4]),
    .c(\u2_Display/n [5]),
    .d(\u2_Display/n [6]),
    .o(_al_u1347_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u1348 (
    .a(_al_u1347_o),
    .b(\u2_Display/n [7]),
    .c(\u2_Display/n [8]),
    .d(\u2_Display/n [9]),
    .o(_al_u1348_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u1349 (
    .a(\u2_Display/n [12]),
    .b(\u2_Display/n [13]),
    .c(\u2_Display/n [14]),
    .d(\u2_Display/n [15]),
    .o(_al_u1349_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'h0010))
    _al_u1350 (
    .a(\u2_Display/n [0]),
    .b(\u2_Display/n [1]),
    .c(\u2_Display/n [10]),
    .d(\u2_Display/n [11]),
    .o(_al_u1350_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1351 (
    .a(\u2_Display/n [2]),
    .b(\u2_Display/n [20]),
    .c(\u2_Display/n [21]),
    .d(\u2_Display/n [22]),
    .o(_al_u1351_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1352 (
    .a(\u2_Display/n [16]),
    .b(\u2_Display/n [17]),
    .c(\u2_Display/n [18]),
    .d(\u2_Display/n [19]),
    .o(_al_u1352_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1353 (
    .a(_al_u1349_o),
    .b(_al_u1350_o),
    .c(_al_u1351_o),
    .d(_al_u1352_o),
    .o(_al_u1353_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1354 (
    .a(_al_u1353_o),
    .b(_al_u1348_o),
    .c(_al_u1345_o),
    .d(_al_u1346_o),
    .o(\u2_Display/n35 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1355 (
    .a(\u2_Display/n3995 ),
    .b(\u2_Display/n3998 [0]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4030 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1356 (
    .a(\u2_Display/n3994 ),
    .b(\u2_Display/n3998 [1]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4029 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1357 (
    .a(\u2_Display/n3993 ),
    .b(\u2_Display/n3998 [2]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4028 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1358 (
    .a(\u2_Display/n3992 ),
    .b(\u2_Display/n3998 [3]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4027 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1359 (
    .a(\u2_Display/n3991 ),
    .b(\u2_Display/n3998 [4]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4026 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1360 (
    .a(\u2_Display/n3990 ),
    .b(\u2_Display/n3998 [5]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4025 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1361 (
    .a(\u2_Display/n3989 ),
    .b(\u2_Display/n3998 [6]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4024 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1362 (
    .a(\u2_Display/n3988 ),
    .b(\u2_Display/n3998 [7]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4023 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1363 (
    .a(\u2_Display/n3987 ),
    .b(\u2_Display/n3998 [8]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4022 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1364 (
    .a(\u2_Display/n3986 ),
    .b(\u2_Display/n3998 [9]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4021 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1365 (
    .a(\u2_Display/n3985 ),
    .b(\u2_Display/n3998 [10]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4020 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1366 (
    .a(\u2_Display/n3984 ),
    .b(\u2_Display/n3998 [11]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4019 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1367 (
    .a(\u2_Display/n3983 ),
    .b(\u2_Display/n3998 [12]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4018 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1368 (
    .a(\u2_Display/n3982 ),
    .b(\u2_Display/n3998 [13]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4017 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1369 (
    .a(\u2_Display/n3981 ),
    .b(\u2_Display/n3998 [14]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4016 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1370 (
    .a(\u2_Display/n3980 ),
    .b(\u2_Display/n3998 [15]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4015 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1371 (
    .a(\u2_Display/n3979 ),
    .b(\u2_Display/n3998 [16]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4014 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1372 (
    .a(\u2_Display/n3978 ),
    .b(\u2_Display/n3998 [17]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4013 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1373 (
    .a(\u2_Display/n3977 ),
    .b(\u2_Display/n3998 [18]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4012 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1374 (
    .a(\u2_Display/n3976 ),
    .b(\u2_Display/n3998 [19]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4011 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1375 (
    .a(\u2_Display/n3975 ),
    .b(\u2_Display/n3998 [20]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4010 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1376 (
    .a(\u2_Display/n3974 ),
    .b(\u2_Display/n3998 [21]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4009 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1377 (
    .a(\u2_Display/n3973 ),
    .b(\u2_Display/n3998 [22]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4008 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1378 (
    .a(\u2_Display/n3972 ),
    .b(\u2_Display/n3998 [23]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4007 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1379 (
    .a(\u2_Display/n3971 ),
    .b(\u2_Display/n3998 [24]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4006 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1380 (
    .a(\u2_Display/n3970 ),
    .b(\u2_Display/n3998 [25]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4005 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1381 (
    .a(\u2_Display/n3969 ),
    .b(\u2_Display/n3998 [26]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4004 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1382 (
    .a(\u2_Display/n3968 ),
    .b(\u2_Display/n3998 [27]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4003 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1383 (
    .a(\u2_Display/n3967 ),
    .b(\u2_Display/n3998 [28]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4002 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1384 (
    .a(\u2_Display/n3966 ),
    .b(\u2_Display/n3998 [29]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4001 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1385 (
    .a(\u2_Display/n3965 ),
    .b(\u2_Display/n3998 [30]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n4000 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1386 (
    .a(\u2_Display/n3964 ),
    .b(\u2_Display/n3998 [31]),
    .c(\u2_Display/n3996 ),
    .o(\u2_Display/n3999 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1387 (
    .a(\u2_Display/n6276 ),
    .b(\u2_Display/n5121 [0]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6311 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1388 (
    .a(\u2_Display/n6275 ),
    .b(\u2_Display/n5121 [1]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6310 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1389 (
    .a(\u2_Display/n6274 ),
    .b(\u2_Display/n5121 [2]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6309 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1390 (
    .a(\u2_Display/n6273 ),
    .b(\u2_Display/n5121 [3]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6308 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1391 (
    .a(\u2_Display/n6272 ),
    .b(\u2_Display/n5121 [4]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6307 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1392 (
    .a(\u2_Display/n6271 ),
    .b(\u2_Display/n5121 [5]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6306 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1393 (
    .a(\u2_Display/n6270 ),
    .b(\u2_Display/n5121 [6]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6305 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1394 (
    .a(\u2_Display/n6269 ),
    .b(\u2_Display/n5121 [7]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6304 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1395 (
    .a(\u2_Display/n6268 ),
    .b(\u2_Display/n5121 [8]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6303 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1396 (
    .a(\u2_Display/n6267 ),
    .b(\u2_Display/n5121 [9]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6302 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1397 (
    .a(\u2_Display/n6266 ),
    .b(\u2_Display/n5121 [10]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6301 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1398 (
    .a(\u2_Display/n6265 ),
    .b(\u2_Display/n5121 [11]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6300 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1399 (
    .a(\u2_Display/n6264 ),
    .b(\u2_Display/n5121 [12]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6299 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1400 (
    .a(\u2_Display/n6263 ),
    .b(\u2_Display/n5121 [13]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6298 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1401 (
    .a(\u2_Display/n6262 ),
    .b(\u2_Display/n5121 [14]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6297 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1402 (
    .a(\u2_Display/n6261 ),
    .b(\u2_Display/n5121 [15]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6296 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1403 (
    .a(\u2_Display/n6260 ),
    .b(\u2_Display/n5121 [16]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6295 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1404 (
    .a(\u2_Display/n6259 ),
    .b(\u2_Display/n5121 [17]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6294 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1405 (
    .a(\u2_Display/n6258 ),
    .b(\u2_Display/n5121 [18]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6293 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1406 (
    .a(\u2_Display/n6257 ),
    .b(\u2_Display/n5121 [19]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6292 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1407 (
    .a(\u2_Display/n6256 ),
    .b(\u2_Display/n5121 [20]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6291 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1408 (
    .a(\u2_Display/n6255 ),
    .b(\u2_Display/n5121 [21]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6290 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1409 (
    .a(\u2_Display/n6254 ),
    .b(\u2_Display/n5121 [22]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6289 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1410 (
    .a(\u2_Display/n6253 ),
    .b(\u2_Display/n5121 [23]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6288 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1411 (
    .a(\u2_Display/n6252 ),
    .b(\u2_Display/n5121 [24]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6287 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1412 (
    .a(\u2_Display/n6251 ),
    .b(\u2_Display/n5121 [25]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6286 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1413 (
    .a(\u2_Display/n6250 ),
    .b(\u2_Display/n5121 [26]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6285 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1414 (
    .a(\u2_Display/n6249 ),
    .b(\u2_Display/n5121 [27]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6284 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1415 (
    .a(\u2_Display/n6248 ),
    .b(\u2_Display/n5121 [28]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6283 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1416 (
    .a(\u2_Display/n6247 ),
    .b(\u2_Display/n5121 [29]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6282 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1417 (
    .a(\u2_Display/n6246 ),
    .b(\u2_Display/n5121 [30]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6281 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1418 (
    .a(\u2_Display/n6245 ),
    .b(\u2_Display/n5121 [31]),
    .c(\u2_Display/n5119 ),
    .o(\u2_Display/n6280 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1419 (
    .a(\u2_Display/n626 ),
    .b(\u2_Display/n629 [0]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n661 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1420 (
    .a(\u2_Display/n625 ),
    .b(\u2_Display/n629 [1]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n660 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1421 (
    .a(\u2_Display/n624 ),
    .b(\u2_Display/n629 [2]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n659 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1422 (
    .a(\u2_Display/n623 ),
    .b(\u2_Display/n629 [3]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n658 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1423 (
    .a(\u2_Display/n622 ),
    .b(\u2_Display/n629 [4]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n657 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1424 (
    .a(\u2_Display/n621 ),
    .b(\u2_Display/n629 [5]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n656 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1425 (
    .a(\u2_Display/n620 ),
    .b(\u2_Display/n629 [6]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n655 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1426 (
    .a(\u2_Display/n619 ),
    .b(\u2_Display/n629 [7]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n654 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1427 (
    .a(\u2_Display/n618 ),
    .b(\u2_Display/n629 [8]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n653 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1428 (
    .a(\u2_Display/n617 ),
    .b(\u2_Display/n629 [9]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n652 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1429 (
    .a(\u2_Display/n616 ),
    .b(\u2_Display/n629 [10]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n651 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1430 (
    .a(\u2_Display/n615 ),
    .b(\u2_Display/n629 [11]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n650 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1431 (
    .a(\u2_Display/n614 ),
    .b(\u2_Display/n629 [12]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n649 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1432 (
    .a(\u2_Display/n613 ),
    .b(\u2_Display/n629 [13]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n648 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1433 (
    .a(\u2_Display/n612 ),
    .b(\u2_Display/n629 [14]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n647 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1434 (
    .a(\u2_Display/n611 ),
    .b(\u2_Display/n629 [15]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n646 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1435 (
    .a(\u2_Display/n610 ),
    .b(\u2_Display/n629 [16]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n645 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1436 (
    .a(\u2_Display/n609 ),
    .b(\u2_Display/n629 [17]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n644 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1437 (
    .a(\u2_Display/n608 ),
    .b(\u2_Display/n629 [18]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n643 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1438 (
    .a(\u2_Display/n607 ),
    .b(\u2_Display/n629 [19]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n642 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1439 (
    .a(\u2_Display/n606 ),
    .b(\u2_Display/n629 [20]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n641 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1440 (
    .a(\u2_Display/n605 ),
    .b(\u2_Display/n629 [21]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n640 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1441 (
    .a(\u2_Display/n604 ),
    .b(\u2_Display/n629 [22]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n639 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1442 (
    .a(\u2_Display/n603 ),
    .b(\u2_Display/n629 [23]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n638 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1443 (
    .a(\u2_Display/n602 ),
    .b(\u2_Display/n629 [24]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n637 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1444 (
    .a(\u2_Display/n601 ),
    .b(\u2_Display/n629 [25]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n636 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1445 (
    .a(\u2_Display/n600 ),
    .b(\u2_Display/n629 [26]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n635 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1446 (
    .a(\u2_Display/n599 ),
    .b(\u2_Display/n629 [27]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n634 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1447 (
    .a(\u2_Display/n598 ),
    .b(\u2_Display/n629 [28]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n633 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1448 (
    .a(\u2_Display/n597 ),
    .b(\u2_Display/n629 [29]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n632 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1449 (
    .a(\u2_Display/n596 ),
    .b(\u2_Display/n629 [30]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n631 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1450 (
    .a(\u2_Display/n595 ),
    .b(\u2_Display/n629 [31]),
    .c(\u2_Display/n627 ),
    .o(\u2_Display/n630 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1451 (
    .a(\u2_Display/n1749 ),
    .b(\u2_Display/n1752 [0]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1784 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1452 (
    .a(\u2_Display/n1748 ),
    .b(\u2_Display/n1752 [1]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1783 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1453 (
    .a(\u2_Display/n1747 ),
    .b(\u2_Display/n1752 [2]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1782 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1454 (
    .a(\u2_Display/n1746 ),
    .b(\u2_Display/n1752 [3]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1781 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1455 (
    .a(\u2_Display/n1745 ),
    .b(\u2_Display/n1752 [4]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1780 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1456 (
    .a(\u2_Display/n1744 ),
    .b(\u2_Display/n1752 [5]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1779 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1457 (
    .a(\u2_Display/n1743 ),
    .b(\u2_Display/n1752 [6]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1778 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1458 (
    .a(\u2_Display/n1742 ),
    .b(\u2_Display/n1752 [7]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1777 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1459 (
    .a(\u2_Display/n1741 ),
    .b(\u2_Display/n1752 [8]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1776 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1460 (
    .a(\u2_Display/n1740 ),
    .b(\u2_Display/n1752 [9]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1775 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1461 (
    .a(\u2_Display/n1739 ),
    .b(\u2_Display/n1752 [10]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1774 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1462 (
    .a(\u2_Display/n1738 ),
    .b(\u2_Display/n1752 [11]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1773 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1463 (
    .a(\u2_Display/n1737 ),
    .b(\u2_Display/n1752 [12]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1772 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1464 (
    .a(\u2_Display/n1736 ),
    .b(\u2_Display/n1752 [13]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1771 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1465 (
    .a(\u2_Display/n1735 ),
    .b(\u2_Display/n1752 [14]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1770 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1466 (
    .a(\u2_Display/n1734 ),
    .b(\u2_Display/n1752 [15]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1769 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1467 (
    .a(\u2_Display/n1733 ),
    .b(\u2_Display/n1752 [16]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1768 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1468 (
    .a(\u2_Display/n1732 ),
    .b(\u2_Display/n1752 [17]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1767 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1469 (
    .a(\u2_Display/n1731 ),
    .b(\u2_Display/n1752 [18]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1766 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1470 (
    .a(\u2_Display/n1730 ),
    .b(\u2_Display/n1752 [19]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1765 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1471 (
    .a(\u2_Display/n1729 ),
    .b(\u2_Display/n1752 [20]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1764 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1472 (
    .a(\u2_Display/n1728 ),
    .b(\u2_Display/n1752 [21]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1763 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1473 (
    .a(\u2_Display/n1727 ),
    .b(\u2_Display/n1752 [22]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1762 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1474 (
    .a(\u2_Display/n1726 ),
    .b(\u2_Display/n1752 [23]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1761 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1475 (
    .a(\u2_Display/n1725 ),
    .b(\u2_Display/n1752 [24]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1760 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1476 (
    .a(\u2_Display/n1724 ),
    .b(\u2_Display/n1752 [25]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1759 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1477 (
    .a(\u2_Display/n1723 ),
    .b(\u2_Display/n1752 [26]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1758 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1478 (
    .a(\u2_Display/n1722 ),
    .b(\u2_Display/n1752 [27]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1757 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1479 (
    .a(\u2_Display/n1721 ),
    .b(\u2_Display/n1752 [28]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1756 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1480 (
    .a(\u2_Display/n1720 ),
    .b(\u2_Display/n1752 [29]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1755 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1481 (
    .a(\u2_Display/n1719 ),
    .b(\u2_Display/n1752 [30]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1754 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1482 (
    .a(\u2_Display/n1718 ),
    .b(\u2_Display/n1752 [31]),
    .c(\u2_Display/n1750 ),
    .o(\u2_Display/n1753 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1483 (
    .a(\u2_Display/n2872 ),
    .b(\u2_Display/n2875 [0]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2907 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1484 (
    .a(\u2_Display/n2871 ),
    .b(\u2_Display/n2875 [1]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2906 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1485 (
    .a(\u2_Display/n2870 ),
    .b(\u2_Display/n2875 [2]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2905 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1486 (
    .a(\u2_Display/n2869 ),
    .b(\u2_Display/n2875 [3]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2904 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1487 (
    .a(\u2_Display/n2868 ),
    .b(\u2_Display/n2875 [4]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2903 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1488 (
    .a(\u2_Display/n2867 ),
    .b(\u2_Display/n2875 [5]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2902 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1489 (
    .a(\u2_Display/n2866 ),
    .b(\u2_Display/n2875 [6]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2901 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1490 (
    .a(\u2_Display/n2865 ),
    .b(\u2_Display/n2875 [7]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2900 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1491 (
    .a(\u2_Display/n2864 ),
    .b(\u2_Display/n2875 [8]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2899 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1492 (
    .a(\u2_Display/n2863 ),
    .b(\u2_Display/n2875 [9]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2898 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1493 (
    .a(\u2_Display/n2862 ),
    .b(\u2_Display/n2875 [10]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2897 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1494 (
    .a(\u2_Display/n2861 ),
    .b(\u2_Display/n2875 [11]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2896 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1495 (
    .a(\u2_Display/n2860 ),
    .b(\u2_Display/n2875 [12]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2895 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1496 (
    .a(\u2_Display/n2859 ),
    .b(\u2_Display/n2875 [13]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2894 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1497 (
    .a(\u2_Display/n2858 ),
    .b(\u2_Display/n2875 [14]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2893 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1498 (
    .a(\u2_Display/n2857 ),
    .b(\u2_Display/n2875 [15]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2892 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1499 (
    .a(\u2_Display/n2856 ),
    .b(\u2_Display/n2875 [16]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2891 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1500 (
    .a(\u2_Display/n2855 ),
    .b(\u2_Display/n2875 [17]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2890 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1501 (
    .a(\u2_Display/n2854 ),
    .b(\u2_Display/n2875 [18]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2889 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1502 (
    .a(\u2_Display/n2853 ),
    .b(\u2_Display/n2875 [19]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2888 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1503 (
    .a(\u2_Display/n2852 ),
    .b(\u2_Display/n2875 [20]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2887 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1504 (
    .a(\u2_Display/n2851 ),
    .b(\u2_Display/n2875 [21]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2886 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1505 (
    .a(\u2_Display/n2850 ),
    .b(\u2_Display/n2875 [22]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2885 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1506 (
    .a(\u2_Display/n2849 ),
    .b(\u2_Display/n2875 [23]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2884 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1507 (
    .a(\u2_Display/n2848 ),
    .b(\u2_Display/n2875 [24]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2883 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1508 (
    .a(\u2_Display/n2847 ),
    .b(\u2_Display/n2875 [25]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2882 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1509 (
    .a(\u2_Display/n2846 ),
    .b(\u2_Display/n2875 [26]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2881 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1510 (
    .a(\u2_Display/n2845 ),
    .b(\u2_Display/n2875 [27]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2880 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1511 (
    .a(\u2_Display/n2844 ),
    .b(\u2_Display/n2875 [28]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2879 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1512 (
    .a(\u2_Display/n2843 ),
    .b(\u2_Display/n2875 [29]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2878 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1513 (
    .a(\u2_Display/n2842 ),
    .b(\u2_Display/n2875 [30]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2877 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1514 (
    .a(\u2_Display/n2841 ),
    .b(\u2_Display/n2875 [31]),
    .c(\u2_Display/n2873 ),
    .o(\u2_Display/n2876 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1515 (
    .a(\u2_Display/n4030 ),
    .b(\u2_Display/n4033 [0]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4065 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1516 (
    .a(\u2_Display/n4029 ),
    .b(\u2_Display/n4033 [1]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4064 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1517 (
    .a(\u2_Display/n4028 ),
    .b(\u2_Display/n4033 [2]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4063 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1518 (
    .a(\u2_Display/n4027 ),
    .b(\u2_Display/n4033 [3]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4062 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1519 (
    .a(\u2_Display/n4026 ),
    .b(\u2_Display/n4033 [4]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4061 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1520 (
    .a(\u2_Display/n4025 ),
    .b(\u2_Display/n4033 [5]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4060 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1521 (
    .a(\u2_Display/n4024 ),
    .b(\u2_Display/n4033 [6]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4059 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1522 (
    .a(\u2_Display/n4023 ),
    .b(\u2_Display/n4033 [7]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4058 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1523 (
    .a(\u2_Display/n4022 ),
    .b(\u2_Display/n4033 [8]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4057 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1524 (
    .a(\u2_Display/n4021 ),
    .b(\u2_Display/n4033 [9]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4056 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1525 (
    .a(\u2_Display/n4020 ),
    .b(\u2_Display/n4033 [10]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4055 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1526 (
    .a(\u2_Display/n4019 ),
    .b(\u2_Display/n4033 [11]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4054 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1527 (
    .a(\u2_Display/n4018 ),
    .b(\u2_Display/n4033 [12]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4053 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1528 (
    .a(\u2_Display/n4017 ),
    .b(\u2_Display/n4033 [13]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4052 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1529 (
    .a(\u2_Display/n4016 ),
    .b(\u2_Display/n4033 [14]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4051 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1530 (
    .a(\u2_Display/n4015 ),
    .b(\u2_Display/n4033 [15]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4050 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1531 (
    .a(\u2_Display/n4014 ),
    .b(\u2_Display/n4033 [16]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4049 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1532 (
    .a(\u2_Display/n4013 ),
    .b(\u2_Display/n4033 [17]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4048 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1533 (
    .a(\u2_Display/n4012 ),
    .b(\u2_Display/n4033 [18]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4047 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1534 (
    .a(\u2_Display/n4011 ),
    .b(\u2_Display/n4033 [19]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4046 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1535 (
    .a(\u2_Display/n4010 ),
    .b(\u2_Display/n4033 [20]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4045 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1536 (
    .a(\u2_Display/n4009 ),
    .b(\u2_Display/n4033 [21]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4044 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1537 (
    .a(\u2_Display/n4008 ),
    .b(\u2_Display/n4033 [22]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4043 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1538 (
    .a(\u2_Display/n4007 ),
    .b(\u2_Display/n4033 [23]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4042 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1539 (
    .a(\u2_Display/n4006 ),
    .b(\u2_Display/n4033 [24]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4041 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1540 (
    .a(\u2_Display/n4005 ),
    .b(\u2_Display/n4033 [25]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4040 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1541 (
    .a(\u2_Display/n4004 ),
    .b(\u2_Display/n4033 [26]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4039 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1542 (
    .a(\u2_Display/n4003 ),
    .b(\u2_Display/n4033 [27]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4038 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1543 (
    .a(\u2_Display/n4002 ),
    .b(\u2_Display/n4033 [28]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4037 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1544 (
    .a(\u2_Display/n4001 ),
    .b(\u2_Display/n4033 [29]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4036 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1545 (
    .a(\u2_Display/n4000 ),
    .b(\u2_Display/n4033 [30]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4035 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1546 (
    .a(\u2_Display/n3999 ),
    .b(\u2_Display/n4033 [31]),
    .c(\u2_Display/n4031 ),
    .o(\u2_Display/n4034 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1547 (
    .a(\u2_Display/n6311 ),
    .b(\u2_Display/n5156 [0]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6346 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1548 (
    .a(\u2_Display/n6310 ),
    .b(\u2_Display/n5156 [1]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6345 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1549 (
    .a(\u2_Display/n6309 ),
    .b(\u2_Display/n5156 [2]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6344 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1550 (
    .a(\u2_Display/n6308 ),
    .b(\u2_Display/n5156 [3]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6343 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1551 (
    .a(\u2_Display/n6307 ),
    .b(\u2_Display/n5156 [4]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6342 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1552 (
    .a(\u2_Display/n6306 ),
    .b(\u2_Display/n5156 [5]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6341 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1553 (
    .a(\u2_Display/n6305 ),
    .b(\u2_Display/n5156 [6]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6340 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1554 (
    .a(\u2_Display/n6304 ),
    .b(\u2_Display/n5156 [7]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6339 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1555 (
    .a(\u2_Display/n6303 ),
    .b(\u2_Display/n5156 [8]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6338 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1556 (
    .a(\u2_Display/n6302 ),
    .b(\u2_Display/n5156 [9]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6337 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1557 (
    .a(\u2_Display/n6301 ),
    .b(\u2_Display/n5156 [10]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6336 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1558 (
    .a(\u2_Display/n6300 ),
    .b(\u2_Display/n5156 [11]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6335 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1559 (
    .a(\u2_Display/n6299 ),
    .b(\u2_Display/n5156 [12]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6334 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1560 (
    .a(\u2_Display/n6298 ),
    .b(\u2_Display/n5156 [13]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6333 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1561 (
    .a(\u2_Display/n6297 ),
    .b(\u2_Display/n5156 [14]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6332 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1562 (
    .a(\u2_Display/n6296 ),
    .b(\u2_Display/n5156 [15]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6331 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1563 (
    .a(\u2_Display/n6295 ),
    .b(\u2_Display/n5156 [16]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6330 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1564 (
    .a(\u2_Display/n6294 ),
    .b(\u2_Display/n5156 [17]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6329 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1565 (
    .a(\u2_Display/n6293 ),
    .b(\u2_Display/n5156 [18]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6328 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1566 (
    .a(\u2_Display/n6292 ),
    .b(\u2_Display/n5156 [19]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6327 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1567 (
    .a(\u2_Display/n6291 ),
    .b(\u2_Display/n5156 [20]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6326 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1568 (
    .a(\u2_Display/n6290 ),
    .b(\u2_Display/n5156 [21]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6325 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1569 (
    .a(\u2_Display/n6289 ),
    .b(\u2_Display/n5156 [22]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6324 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1570 (
    .a(\u2_Display/n6288 ),
    .b(\u2_Display/n5156 [23]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6323 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1571 (
    .a(\u2_Display/n6287 ),
    .b(\u2_Display/n5156 [24]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6322 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1572 (
    .a(\u2_Display/n6286 ),
    .b(\u2_Display/n5156 [25]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6321 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1573 (
    .a(\u2_Display/n6285 ),
    .b(\u2_Display/n5156 [26]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6320 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1574 (
    .a(\u2_Display/n6284 ),
    .b(\u2_Display/n5156 [27]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6319 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1575 (
    .a(\u2_Display/n6283 ),
    .b(\u2_Display/n5156 [28]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6318 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1576 (
    .a(\u2_Display/n6282 ),
    .b(\u2_Display/n5156 [29]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6317 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1577 (
    .a(\u2_Display/n6281 ),
    .b(\u2_Display/n5156 [30]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6316 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1578 (
    .a(\u2_Display/n6280 ),
    .b(\u2_Display/n5156 [31]),
    .c(\u2_Display/n5154 ),
    .o(\u2_Display/n6315 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1579 (
    .a(\u2_Display/n661 ),
    .b(\u2_Display/n664 [0]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n696 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1580 (
    .a(\u2_Display/n660 ),
    .b(\u2_Display/n664 [1]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n695 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1581 (
    .a(\u2_Display/n659 ),
    .b(\u2_Display/n664 [2]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n694 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1582 (
    .a(\u2_Display/n658 ),
    .b(\u2_Display/n664 [3]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n693 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1583 (
    .a(\u2_Display/n657 ),
    .b(\u2_Display/n664 [4]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n692 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1584 (
    .a(\u2_Display/n656 ),
    .b(\u2_Display/n664 [5]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n691 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1585 (
    .a(\u2_Display/n655 ),
    .b(\u2_Display/n664 [6]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n690 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1586 (
    .a(\u2_Display/n654 ),
    .b(\u2_Display/n664 [7]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n689 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1587 (
    .a(\u2_Display/n653 ),
    .b(\u2_Display/n664 [8]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n688 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1588 (
    .a(\u2_Display/n652 ),
    .b(\u2_Display/n664 [9]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n687 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1589 (
    .a(\u2_Display/n651 ),
    .b(\u2_Display/n664 [10]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n686 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1590 (
    .a(\u2_Display/n650 ),
    .b(\u2_Display/n664 [11]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n685 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1591 (
    .a(\u2_Display/n649 ),
    .b(\u2_Display/n664 [12]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n684 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1592 (
    .a(\u2_Display/n648 ),
    .b(\u2_Display/n664 [13]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n683 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1593 (
    .a(\u2_Display/n647 ),
    .b(\u2_Display/n664 [14]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n682 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1594 (
    .a(\u2_Display/n646 ),
    .b(\u2_Display/n664 [15]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n681 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1595 (
    .a(\u2_Display/n645 ),
    .b(\u2_Display/n664 [16]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n680 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1596 (
    .a(\u2_Display/n644 ),
    .b(\u2_Display/n664 [17]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n679 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1597 (
    .a(\u2_Display/n643 ),
    .b(\u2_Display/n664 [18]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n678 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1598 (
    .a(\u2_Display/n642 ),
    .b(\u2_Display/n664 [19]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n677 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1599 (
    .a(\u2_Display/n641 ),
    .b(\u2_Display/n664 [20]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n676 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1600 (
    .a(\u2_Display/n640 ),
    .b(\u2_Display/n664 [21]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n675 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1601 (
    .a(\u2_Display/n639 ),
    .b(\u2_Display/n664 [22]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n674 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1602 (
    .a(\u2_Display/n638 ),
    .b(\u2_Display/n664 [23]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n673 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1603 (
    .a(\u2_Display/n637 ),
    .b(\u2_Display/n664 [24]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n672 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1604 (
    .a(\u2_Display/n636 ),
    .b(\u2_Display/n664 [25]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n671 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1605 (
    .a(\u2_Display/n635 ),
    .b(\u2_Display/n664 [26]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n670 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1606 (
    .a(\u2_Display/n634 ),
    .b(\u2_Display/n664 [27]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n669 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1607 (
    .a(\u2_Display/n633 ),
    .b(\u2_Display/n664 [28]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n668 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1608 (
    .a(\u2_Display/n632 ),
    .b(\u2_Display/n664 [29]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n667 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1609 (
    .a(\u2_Display/n631 ),
    .b(\u2_Display/n664 [30]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n666 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1610 (
    .a(\u2_Display/n630 ),
    .b(\u2_Display/n664 [31]),
    .c(\u2_Display/n662 ),
    .o(\u2_Display/n665 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1611 (
    .a(\u2_Display/n1784 ),
    .b(\u2_Display/n1787 [0]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1819 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1612 (
    .a(\u2_Display/n1783 ),
    .b(\u2_Display/n1787 [1]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1818 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1613 (
    .a(\u2_Display/n1782 ),
    .b(\u2_Display/n1787 [2]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1817 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1614 (
    .a(\u2_Display/n1781 ),
    .b(\u2_Display/n1787 [3]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1816 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1615 (
    .a(\u2_Display/n1780 ),
    .b(\u2_Display/n1787 [4]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1815 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1616 (
    .a(\u2_Display/n1779 ),
    .b(\u2_Display/n1787 [5]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1814 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1617 (
    .a(\u2_Display/n1778 ),
    .b(\u2_Display/n1787 [6]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1813 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1618 (
    .a(\u2_Display/n1777 ),
    .b(\u2_Display/n1787 [7]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1812 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1619 (
    .a(\u2_Display/n1776 ),
    .b(\u2_Display/n1787 [8]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1811 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1620 (
    .a(\u2_Display/n1775 ),
    .b(\u2_Display/n1787 [9]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1810 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1621 (
    .a(\u2_Display/n1774 ),
    .b(\u2_Display/n1787 [10]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1809 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1622 (
    .a(\u2_Display/n1773 ),
    .b(\u2_Display/n1787 [11]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1808 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1623 (
    .a(\u2_Display/n1772 ),
    .b(\u2_Display/n1787 [12]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1807 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1624 (
    .a(\u2_Display/n1771 ),
    .b(\u2_Display/n1787 [13]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1806 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1625 (
    .a(\u2_Display/n1770 ),
    .b(\u2_Display/n1787 [14]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1805 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1626 (
    .a(\u2_Display/n1769 ),
    .b(\u2_Display/n1787 [15]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1804 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1627 (
    .a(\u2_Display/n1768 ),
    .b(\u2_Display/n1787 [16]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1803 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1628 (
    .a(\u2_Display/n1767 ),
    .b(\u2_Display/n1787 [17]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1802 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1629 (
    .a(\u2_Display/n1766 ),
    .b(\u2_Display/n1787 [18]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1801 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1630 (
    .a(\u2_Display/n1765 ),
    .b(\u2_Display/n1787 [19]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1800 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1631 (
    .a(\u2_Display/n1764 ),
    .b(\u2_Display/n1787 [20]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1799 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1632 (
    .a(\u2_Display/n1763 ),
    .b(\u2_Display/n1787 [21]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1798 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1633 (
    .a(\u2_Display/n1762 ),
    .b(\u2_Display/n1787 [22]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1797 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1634 (
    .a(\u2_Display/n1761 ),
    .b(\u2_Display/n1787 [23]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1796 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1635 (
    .a(\u2_Display/n1760 ),
    .b(\u2_Display/n1787 [24]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1795 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1636 (
    .a(\u2_Display/n1759 ),
    .b(\u2_Display/n1787 [25]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1794 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1637 (
    .a(\u2_Display/n1758 ),
    .b(\u2_Display/n1787 [26]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1793 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1638 (
    .a(\u2_Display/n1757 ),
    .b(\u2_Display/n1787 [27]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1792 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1639 (
    .a(\u2_Display/n1756 ),
    .b(\u2_Display/n1787 [28]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1791 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1640 (
    .a(\u2_Display/n1755 ),
    .b(\u2_Display/n1787 [29]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1790 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1641 (
    .a(\u2_Display/n1754 ),
    .b(\u2_Display/n1787 [30]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1789 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1642 (
    .a(\u2_Display/n1753 ),
    .b(\u2_Display/n1787 [31]),
    .c(\u2_Display/n1785 ),
    .o(\u2_Display/n1788 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1643 (
    .a(\u2_Display/n2907 ),
    .b(\u2_Display/n2910 [0]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2942 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1644 (
    .a(\u2_Display/n2906 ),
    .b(\u2_Display/n2910 [1]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2941 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1645 (
    .a(\u2_Display/n2905 ),
    .b(\u2_Display/n2910 [2]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2940 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1646 (
    .a(\u2_Display/n2904 ),
    .b(\u2_Display/n2910 [3]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2939 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1647 (
    .a(\u2_Display/n2903 ),
    .b(\u2_Display/n2910 [4]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2938 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1648 (
    .a(\u2_Display/n2902 ),
    .b(\u2_Display/n2910 [5]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2937 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1649 (
    .a(\u2_Display/n2901 ),
    .b(\u2_Display/n2910 [6]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2936 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1650 (
    .a(\u2_Display/n2900 ),
    .b(\u2_Display/n2910 [7]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2935 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1651 (
    .a(\u2_Display/n2899 ),
    .b(\u2_Display/n2910 [8]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2934 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1652 (
    .a(\u2_Display/n2898 ),
    .b(\u2_Display/n2910 [9]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2933 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1653 (
    .a(\u2_Display/n2897 ),
    .b(\u2_Display/n2910 [10]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2932 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1654 (
    .a(\u2_Display/n2896 ),
    .b(\u2_Display/n2910 [11]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2931 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1655 (
    .a(\u2_Display/n2895 ),
    .b(\u2_Display/n2910 [12]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2930 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1656 (
    .a(\u2_Display/n2894 ),
    .b(\u2_Display/n2910 [13]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2929 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1657 (
    .a(\u2_Display/n2893 ),
    .b(\u2_Display/n2910 [14]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2928 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1658 (
    .a(\u2_Display/n2892 ),
    .b(\u2_Display/n2910 [15]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2927 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1659 (
    .a(\u2_Display/n2891 ),
    .b(\u2_Display/n2910 [16]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2926 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1660 (
    .a(\u2_Display/n2890 ),
    .b(\u2_Display/n2910 [17]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2925 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1661 (
    .a(\u2_Display/n2889 ),
    .b(\u2_Display/n2910 [18]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2924 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1662 (
    .a(\u2_Display/n2888 ),
    .b(\u2_Display/n2910 [19]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2923 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1663 (
    .a(\u2_Display/n2887 ),
    .b(\u2_Display/n2910 [20]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2922 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1664 (
    .a(\u2_Display/n2886 ),
    .b(\u2_Display/n2910 [21]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2921 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1665 (
    .a(\u2_Display/n2885 ),
    .b(\u2_Display/n2910 [22]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2920 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1666 (
    .a(\u2_Display/n2884 ),
    .b(\u2_Display/n2910 [23]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2919 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1667 (
    .a(\u2_Display/n2883 ),
    .b(\u2_Display/n2910 [24]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2918 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1668 (
    .a(\u2_Display/n2882 ),
    .b(\u2_Display/n2910 [25]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2917 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1669 (
    .a(\u2_Display/n2881 ),
    .b(\u2_Display/n2910 [26]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2916 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1670 (
    .a(\u2_Display/n2880 ),
    .b(\u2_Display/n2910 [27]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2915 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1671 (
    .a(\u2_Display/n2879 ),
    .b(\u2_Display/n2910 [28]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2914 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1672 (
    .a(\u2_Display/n2878 ),
    .b(\u2_Display/n2910 [29]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2913 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1673 (
    .a(\u2_Display/n2877 ),
    .b(\u2_Display/n2910 [30]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2912 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1674 (
    .a(\u2_Display/n2876 ),
    .b(\u2_Display/n2910 [31]),
    .c(\u2_Display/n2908 ),
    .o(\u2_Display/n2911 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1675 (
    .a(\u2_Display/n4065 ),
    .b(\u2_Display/n4068 [0]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4100 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1676 (
    .a(\u2_Display/n4064 ),
    .b(\u2_Display/n4068 [1]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4099 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1677 (
    .a(\u2_Display/n4063 ),
    .b(\u2_Display/n4068 [2]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4098 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1678 (
    .a(\u2_Display/n4062 ),
    .b(\u2_Display/n4068 [3]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4097 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1679 (
    .a(\u2_Display/n4061 ),
    .b(\u2_Display/n4068 [4]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4096 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1680 (
    .a(\u2_Display/n4060 ),
    .b(\u2_Display/n4068 [5]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4095 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1681 (
    .a(\u2_Display/n4059 ),
    .b(\u2_Display/n4068 [6]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4094 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1682 (
    .a(\u2_Display/n4058 ),
    .b(\u2_Display/n4068 [7]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4093 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1683 (
    .a(\u2_Display/n4057 ),
    .b(\u2_Display/n4068 [8]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4092 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1684 (
    .a(\u2_Display/n4056 ),
    .b(\u2_Display/n4068 [9]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4091 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1685 (
    .a(\u2_Display/n4055 ),
    .b(\u2_Display/n4068 [10]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4090 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1686 (
    .a(\u2_Display/n4054 ),
    .b(\u2_Display/n4068 [11]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4089 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1687 (
    .a(\u2_Display/n4053 ),
    .b(\u2_Display/n4068 [12]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4088 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1688 (
    .a(\u2_Display/n4052 ),
    .b(\u2_Display/n4068 [13]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4087 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1689 (
    .a(\u2_Display/n4051 ),
    .b(\u2_Display/n4068 [14]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4086 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1690 (
    .a(\u2_Display/n4050 ),
    .b(\u2_Display/n4068 [15]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4085 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1691 (
    .a(\u2_Display/n4049 ),
    .b(\u2_Display/n4068 [16]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4084 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1692 (
    .a(\u2_Display/n4048 ),
    .b(\u2_Display/n4068 [17]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4083 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1693 (
    .a(\u2_Display/n4047 ),
    .b(\u2_Display/n4068 [18]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4082 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1694 (
    .a(\u2_Display/n4046 ),
    .b(\u2_Display/n4068 [19]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4081 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1695 (
    .a(\u2_Display/n4045 ),
    .b(\u2_Display/n4068 [20]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4080 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1696 (
    .a(\u2_Display/n4044 ),
    .b(\u2_Display/n4068 [21]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4079 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1697 (
    .a(\u2_Display/n4043 ),
    .b(\u2_Display/n4068 [22]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4078 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1698 (
    .a(\u2_Display/n4042 ),
    .b(\u2_Display/n4068 [23]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4077 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1699 (
    .a(\u2_Display/n4041 ),
    .b(\u2_Display/n4068 [24]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4076 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1700 (
    .a(\u2_Display/n4040 ),
    .b(\u2_Display/n4068 [25]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4075 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1701 (
    .a(\u2_Display/n4039 ),
    .b(\u2_Display/n4068 [26]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4074 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1702 (
    .a(\u2_Display/n4038 ),
    .b(\u2_Display/n4068 [27]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4073 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1703 (
    .a(\u2_Display/n4037 ),
    .b(\u2_Display/n4068 [28]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4072 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1704 (
    .a(\u2_Display/n4036 ),
    .b(\u2_Display/n4068 [29]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4071 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1705 (
    .a(\u2_Display/n4035 ),
    .b(\u2_Display/n4068 [30]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4070 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1706 (
    .a(\u2_Display/n4034 ),
    .b(\u2_Display/n4068 [31]),
    .c(\u2_Display/n4066 ),
    .o(\u2_Display/n4069 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1707 (
    .a(\u2_Display/n6346 ),
    .b(\u2_Display/n5191 [0]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5223 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1708 (
    .a(\u2_Display/n6345 ),
    .b(\u2_Display/n5191 [1]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5222 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1709 (
    .a(\u2_Display/n6344 ),
    .b(\u2_Display/n5191 [2]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5221 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1710 (
    .a(\u2_Display/n6343 ),
    .b(\u2_Display/n5191 [3]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5220 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1711 (
    .a(\u2_Display/n6342 ),
    .b(\u2_Display/n5191 [4]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5219 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1712 (
    .a(\u2_Display/n6341 ),
    .b(\u2_Display/n5191 [5]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5218 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1713 (
    .a(\u2_Display/n6340 ),
    .b(\u2_Display/n5191 [6]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5217 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1714 (
    .a(\u2_Display/n6339 ),
    .b(\u2_Display/n5191 [7]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5216 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1715 (
    .a(\u2_Display/n6338 ),
    .b(\u2_Display/n5191 [8]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5215 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1716 (
    .a(\u2_Display/n6337 ),
    .b(\u2_Display/n5191 [9]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5214 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1717 (
    .a(\u2_Display/n6336 ),
    .b(\u2_Display/n5191 [10]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5213 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1718 (
    .a(\u2_Display/n6335 ),
    .b(\u2_Display/n5191 [11]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5212 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1719 (
    .a(\u2_Display/n6334 ),
    .b(\u2_Display/n5191 [12]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5211 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1720 (
    .a(\u2_Display/n6333 ),
    .b(\u2_Display/n5191 [13]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5210 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1721 (
    .a(\u2_Display/n6332 ),
    .b(\u2_Display/n5191 [14]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5209 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1722 (
    .a(\u2_Display/n6331 ),
    .b(\u2_Display/n5191 [15]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5208 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1723 (
    .a(\u2_Display/n6330 ),
    .b(\u2_Display/n5191 [16]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5207 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1724 (
    .a(\u2_Display/n6329 ),
    .b(\u2_Display/n5191 [17]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5206 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1725 (
    .a(\u2_Display/n6328 ),
    .b(\u2_Display/n5191 [18]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5205 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1726 (
    .a(\u2_Display/n6327 ),
    .b(\u2_Display/n5191 [19]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5204 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1727 (
    .a(\u2_Display/n6326 ),
    .b(\u2_Display/n5191 [20]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5203 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1728 (
    .a(\u2_Display/n6325 ),
    .b(\u2_Display/n5191 [21]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5202 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1729 (
    .a(\u2_Display/n6324 ),
    .b(\u2_Display/n5191 [22]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5201 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1730 (
    .a(\u2_Display/n6323 ),
    .b(\u2_Display/n5191 [23]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5200 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1731 (
    .a(\u2_Display/n6322 ),
    .b(\u2_Display/n5191 [24]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5199 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1732 (
    .a(\u2_Display/n6321 ),
    .b(\u2_Display/n5191 [25]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5198 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1733 (
    .a(\u2_Display/n6320 ),
    .b(\u2_Display/n5191 [26]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5197 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1734 (
    .a(\u2_Display/n6319 ),
    .b(\u2_Display/n5191 [27]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n5196 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1735 (
    .a(\u2_Display/n6318 ),
    .b(\u2_Display/n5191 [28]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n6353 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1736 (
    .a(\u2_Display/n6317 ),
    .b(\u2_Display/n5191 [29]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n6352 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1737 (
    .a(\u2_Display/n6316 ),
    .b(\u2_Display/n5191 [30]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n6351 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1738 (
    .a(\u2_Display/n6315 ),
    .b(\u2_Display/n5191 [31]),
    .c(\u2_Display/n5189 ),
    .o(\u2_Display/n6350 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1739 (
    .a(\u2_Display/n696 ),
    .b(\u2_Display/n699 [0]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n731 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1740 (
    .a(\u2_Display/n695 ),
    .b(\u2_Display/n699 [1]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n730 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1741 (
    .a(\u2_Display/n694 ),
    .b(\u2_Display/n699 [2]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n729 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1742 (
    .a(\u2_Display/n693 ),
    .b(\u2_Display/n699 [3]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n728 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1743 (
    .a(\u2_Display/n692 ),
    .b(\u2_Display/n699 [4]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n727 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1744 (
    .a(\u2_Display/n691 ),
    .b(\u2_Display/n699 [5]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n726 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1745 (
    .a(\u2_Display/n690 ),
    .b(\u2_Display/n699 [6]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n725 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1746 (
    .a(\u2_Display/n689 ),
    .b(\u2_Display/n699 [7]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n724 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1747 (
    .a(\u2_Display/n688 ),
    .b(\u2_Display/n699 [8]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n723 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1748 (
    .a(\u2_Display/n687 ),
    .b(\u2_Display/n699 [9]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n722 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1749 (
    .a(\u2_Display/n686 ),
    .b(\u2_Display/n699 [10]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n721 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1750 (
    .a(\u2_Display/n685 ),
    .b(\u2_Display/n699 [11]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n720 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1751 (
    .a(\u2_Display/n684 ),
    .b(\u2_Display/n699 [12]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n719 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1752 (
    .a(\u2_Display/n683 ),
    .b(\u2_Display/n699 [13]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n718 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1753 (
    .a(\u2_Display/n682 ),
    .b(\u2_Display/n699 [14]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n717 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1754 (
    .a(\u2_Display/n681 ),
    .b(\u2_Display/n699 [15]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n716 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1755 (
    .a(\u2_Display/n680 ),
    .b(\u2_Display/n699 [16]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n715 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1756 (
    .a(\u2_Display/n679 ),
    .b(\u2_Display/n699 [17]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n714 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1757 (
    .a(\u2_Display/n678 ),
    .b(\u2_Display/n699 [18]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n713 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1758 (
    .a(\u2_Display/n677 ),
    .b(\u2_Display/n699 [19]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n712 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1759 (
    .a(\u2_Display/n676 ),
    .b(\u2_Display/n699 [20]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n711 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1760 (
    .a(\u2_Display/n675 ),
    .b(\u2_Display/n699 [21]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n710 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1761 (
    .a(\u2_Display/n674 ),
    .b(\u2_Display/n699 [22]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n709 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1762 (
    .a(\u2_Display/n673 ),
    .b(\u2_Display/n699 [23]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n708 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1763 (
    .a(\u2_Display/n672 ),
    .b(\u2_Display/n699 [24]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n707 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1764 (
    .a(\u2_Display/n671 ),
    .b(\u2_Display/n699 [25]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n706 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1765 (
    .a(\u2_Display/n670 ),
    .b(\u2_Display/n699 [26]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n705 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1766 (
    .a(\u2_Display/n669 ),
    .b(\u2_Display/n699 [27]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n704 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1767 (
    .a(\u2_Display/n668 ),
    .b(\u2_Display/n699 [28]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n703 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1768 (
    .a(\u2_Display/n667 ),
    .b(\u2_Display/n699 [29]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n702 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1769 (
    .a(\u2_Display/n666 ),
    .b(\u2_Display/n699 [30]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n701 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1770 (
    .a(\u2_Display/n665 ),
    .b(\u2_Display/n699 [31]),
    .c(\u2_Display/n697 ),
    .o(\u2_Display/n700 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1771 (
    .a(\u2_Display/n1819 ),
    .b(\u2_Display/n1822 [0]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1854 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1772 (
    .a(\u2_Display/n1818 ),
    .b(\u2_Display/n1822 [1]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1853 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1773 (
    .a(\u2_Display/n1817 ),
    .b(\u2_Display/n1822 [2]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1852 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1774 (
    .a(\u2_Display/n1816 ),
    .b(\u2_Display/n1822 [3]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1851 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1775 (
    .a(\u2_Display/n1815 ),
    .b(\u2_Display/n1822 [4]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1850 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1776 (
    .a(\u2_Display/n1814 ),
    .b(\u2_Display/n1822 [5]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1849 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1777 (
    .a(\u2_Display/n1813 ),
    .b(\u2_Display/n1822 [6]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1848 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1778 (
    .a(\u2_Display/n1812 ),
    .b(\u2_Display/n1822 [7]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1847 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1779 (
    .a(\u2_Display/n1811 ),
    .b(\u2_Display/n1822 [8]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1846 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1780 (
    .a(\u2_Display/n1810 ),
    .b(\u2_Display/n1822 [9]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1845 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1781 (
    .a(\u2_Display/n1809 ),
    .b(\u2_Display/n1822 [10]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1844 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1782 (
    .a(\u2_Display/n1808 ),
    .b(\u2_Display/n1822 [11]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1843 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1783 (
    .a(\u2_Display/n1807 ),
    .b(\u2_Display/n1822 [12]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1842 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1784 (
    .a(\u2_Display/n1806 ),
    .b(\u2_Display/n1822 [13]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1841 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1785 (
    .a(\u2_Display/n1805 ),
    .b(\u2_Display/n1822 [14]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1840 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1786 (
    .a(\u2_Display/n1804 ),
    .b(\u2_Display/n1822 [15]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1839 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1787 (
    .a(\u2_Display/n1803 ),
    .b(\u2_Display/n1822 [16]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1838 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1788 (
    .a(\u2_Display/n1802 ),
    .b(\u2_Display/n1822 [17]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1837 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1789 (
    .a(\u2_Display/n1801 ),
    .b(\u2_Display/n1822 [18]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1836 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1790 (
    .a(\u2_Display/n1800 ),
    .b(\u2_Display/n1822 [19]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1835 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1791 (
    .a(\u2_Display/n1799 ),
    .b(\u2_Display/n1822 [20]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1834 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1792 (
    .a(\u2_Display/n1798 ),
    .b(\u2_Display/n1822 [21]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1833 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1793 (
    .a(\u2_Display/n1797 ),
    .b(\u2_Display/n1822 [22]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1832 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1794 (
    .a(\u2_Display/n1796 ),
    .b(\u2_Display/n1822 [23]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1831 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1795 (
    .a(\u2_Display/n1795 ),
    .b(\u2_Display/n1822 [24]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1830 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1796 (
    .a(\u2_Display/n1794 ),
    .b(\u2_Display/n1822 [25]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1829 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1797 (
    .a(\u2_Display/n1793 ),
    .b(\u2_Display/n1822 [26]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1828 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1798 (
    .a(\u2_Display/n1792 ),
    .b(\u2_Display/n1822 [27]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1827 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1799 (
    .a(\u2_Display/n1791 ),
    .b(\u2_Display/n1822 [28]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1826 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1800 (
    .a(\u2_Display/n1790 ),
    .b(\u2_Display/n1822 [29]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1825 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1801 (
    .a(\u2_Display/n1789 ),
    .b(\u2_Display/n1822 [30]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1824 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1802 (
    .a(\u2_Display/n1788 ),
    .b(\u2_Display/n1822 [31]),
    .c(\u2_Display/n1820 ),
    .o(\u2_Display/n1823 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1803 (
    .a(\u2_Display/n2942 ),
    .b(\u2_Display/n2945 [0]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2977 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1804 (
    .a(\u2_Display/n2941 ),
    .b(\u2_Display/n2945 [1]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2976 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1805 (
    .a(\u2_Display/n2940 ),
    .b(\u2_Display/n2945 [2]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2975 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1806 (
    .a(\u2_Display/n2939 ),
    .b(\u2_Display/n2945 [3]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2974 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1807 (
    .a(\u2_Display/n2938 ),
    .b(\u2_Display/n2945 [4]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2973 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1808 (
    .a(\u2_Display/n2937 ),
    .b(\u2_Display/n2945 [5]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2972 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1809 (
    .a(\u2_Display/n2936 ),
    .b(\u2_Display/n2945 [6]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2971 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1810 (
    .a(\u2_Display/n2935 ),
    .b(\u2_Display/n2945 [7]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2970 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1811 (
    .a(\u2_Display/n2934 ),
    .b(\u2_Display/n2945 [8]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2969 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1812 (
    .a(\u2_Display/n2933 ),
    .b(\u2_Display/n2945 [9]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2968 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1813 (
    .a(\u2_Display/n2932 ),
    .b(\u2_Display/n2945 [10]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2967 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1814 (
    .a(\u2_Display/n2931 ),
    .b(\u2_Display/n2945 [11]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2966 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1815 (
    .a(\u2_Display/n2930 ),
    .b(\u2_Display/n2945 [12]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2965 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1816 (
    .a(\u2_Display/n2929 ),
    .b(\u2_Display/n2945 [13]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2964 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1817 (
    .a(\u2_Display/n2928 ),
    .b(\u2_Display/n2945 [14]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2963 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1818 (
    .a(\u2_Display/n2927 ),
    .b(\u2_Display/n2945 [15]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2962 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1819 (
    .a(\u2_Display/n2926 ),
    .b(\u2_Display/n2945 [16]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2961 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1820 (
    .a(\u2_Display/n2925 ),
    .b(\u2_Display/n2945 [17]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2960 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1821 (
    .a(\u2_Display/n2924 ),
    .b(\u2_Display/n2945 [18]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2959 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1822 (
    .a(\u2_Display/n2923 ),
    .b(\u2_Display/n2945 [19]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2958 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1823 (
    .a(\u2_Display/n2922 ),
    .b(\u2_Display/n2945 [20]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2957 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1824 (
    .a(\u2_Display/n2921 ),
    .b(\u2_Display/n2945 [21]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2956 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1825 (
    .a(\u2_Display/n2920 ),
    .b(\u2_Display/n2945 [22]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2955 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1826 (
    .a(\u2_Display/n2919 ),
    .b(\u2_Display/n2945 [23]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2954 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1827 (
    .a(\u2_Display/n2918 ),
    .b(\u2_Display/n2945 [24]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2953 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1828 (
    .a(\u2_Display/n2917 ),
    .b(\u2_Display/n2945 [25]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2952 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1829 (
    .a(\u2_Display/n2916 ),
    .b(\u2_Display/n2945 [26]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2951 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1830 (
    .a(\u2_Display/n2915 ),
    .b(\u2_Display/n2945 [27]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2950 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1831 (
    .a(\u2_Display/n2914 ),
    .b(\u2_Display/n2945 [28]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2949 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1832 (
    .a(\u2_Display/n2913 ),
    .b(\u2_Display/n2945 [29]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2948 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1833 (
    .a(\u2_Display/n2912 ),
    .b(\u2_Display/n2945 [30]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2947 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1834 (
    .a(\u2_Display/n2911 ),
    .b(\u2_Display/n2945 [31]),
    .c(\u2_Display/n2943 ),
    .o(\u2_Display/n2946 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1835 (
    .a(\u2_Display/n4100 ),
    .b(\u2_Display/n4103 [0]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4135 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1836 (
    .a(\u2_Display/n4099 ),
    .b(\u2_Display/n4103 [1]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4134 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1837 (
    .a(\u2_Display/n4098 ),
    .b(\u2_Display/n4103 [2]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4133 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1838 (
    .a(\u2_Display/n4097 ),
    .b(\u2_Display/n4103 [3]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4132 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1839 (
    .a(\u2_Display/n4096 ),
    .b(\u2_Display/n4103 [4]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4131 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1840 (
    .a(\u2_Display/n4095 ),
    .b(\u2_Display/n4103 [5]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4130 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1841 (
    .a(\u2_Display/n4094 ),
    .b(\u2_Display/n4103 [6]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4129 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1842 (
    .a(\u2_Display/n4093 ),
    .b(\u2_Display/n4103 [7]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4128 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1843 (
    .a(\u2_Display/n4092 ),
    .b(\u2_Display/n4103 [8]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4127 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1844 (
    .a(\u2_Display/n4091 ),
    .b(\u2_Display/n4103 [9]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4126 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1845 (
    .a(\u2_Display/n4090 ),
    .b(\u2_Display/n4103 [10]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4125 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1846 (
    .a(\u2_Display/n4089 ),
    .b(\u2_Display/n4103 [11]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4124 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1847 (
    .a(\u2_Display/n4088 ),
    .b(\u2_Display/n4103 [12]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4123 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1848 (
    .a(\u2_Display/n4087 ),
    .b(\u2_Display/n4103 [13]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4122 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1849 (
    .a(\u2_Display/n4086 ),
    .b(\u2_Display/n4103 [14]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4121 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1850 (
    .a(\u2_Display/n4085 ),
    .b(\u2_Display/n4103 [15]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4120 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1851 (
    .a(\u2_Display/n4084 ),
    .b(\u2_Display/n4103 [16]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4119 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1852 (
    .a(\u2_Display/n4083 ),
    .b(\u2_Display/n4103 [17]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4118 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1853 (
    .a(\u2_Display/n4082 ),
    .b(\u2_Display/n4103 [18]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4117 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1854 (
    .a(\u2_Display/n4081 ),
    .b(\u2_Display/n4103 [19]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4116 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1855 (
    .a(\u2_Display/n4080 ),
    .b(\u2_Display/n4103 [20]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4115 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1856 (
    .a(\u2_Display/n4079 ),
    .b(\u2_Display/n4103 [21]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4114 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1857 (
    .a(\u2_Display/n4078 ),
    .b(\u2_Display/n4103 [22]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4113 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1858 (
    .a(\u2_Display/n4077 ),
    .b(\u2_Display/n4103 [23]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4112 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1859 (
    .a(\u2_Display/n4076 ),
    .b(\u2_Display/n4103 [24]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4111 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1860 (
    .a(\u2_Display/n4075 ),
    .b(\u2_Display/n4103 [25]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4110 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1861 (
    .a(\u2_Display/n4074 ),
    .b(\u2_Display/n4103 [26]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4109 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1862 (
    .a(\u2_Display/n4073 ),
    .b(\u2_Display/n4103 [27]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4108 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1863 (
    .a(\u2_Display/n4072 ),
    .b(\u2_Display/n4103 [28]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4107 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1864 (
    .a(\u2_Display/n4071 ),
    .b(\u2_Display/n4103 [29]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4106 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1865 (
    .a(\u2_Display/n4070 ),
    .b(\u2_Display/n4103 [30]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4105 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1866 (
    .a(\u2_Display/n4069 ),
    .b(\u2_Display/n4103 [31]),
    .c(\u2_Display/n4101 ),
    .o(\u2_Display/n4104 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1867 (
    .a(\u2_Display/n5223 ),
    .b(\u2_Display/n5226 [0]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5258 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1868 (
    .a(\u2_Display/n5222 ),
    .b(\u2_Display/n5226 [1]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5257 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1869 (
    .a(\u2_Display/n5221 ),
    .b(\u2_Display/n5226 [2]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5256 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1870 (
    .a(\u2_Display/n5220 ),
    .b(\u2_Display/n5226 [3]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5255 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1871 (
    .a(\u2_Display/n5219 ),
    .b(\u2_Display/n5226 [4]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5254 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1872 (
    .a(\u2_Display/n5218 ),
    .b(\u2_Display/n5226 [5]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5253 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1873 (
    .a(\u2_Display/n5217 ),
    .b(\u2_Display/n5226 [6]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5252 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1874 (
    .a(\u2_Display/n5216 ),
    .b(\u2_Display/n5226 [7]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5251 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1875 (
    .a(\u2_Display/n5215 ),
    .b(\u2_Display/n5226 [8]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5250 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1876 (
    .a(\u2_Display/n5214 ),
    .b(\u2_Display/n5226 [9]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5249 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1877 (
    .a(\u2_Display/n5213 ),
    .b(\u2_Display/n5226 [10]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5248 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1878 (
    .a(\u2_Display/n5212 ),
    .b(\u2_Display/n5226 [11]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5247 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1879 (
    .a(\u2_Display/n5211 ),
    .b(\u2_Display/n5226 [12]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5246 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1880 (
    .a(\u2_Display/n5210 ),
    .b(\u2_Display/n5226 [13]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5245 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1881 (
    .a(\u2_Display/n5209 ),
    .b(\u2_Display/n5226 [14]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5244 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1882 (
    .a(\u2_Display/n5208 ),
    .b(\u2_Display/n5226 [15]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5243 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1883 (
    .a(\u2_Display/n5207 ),
    .b(\u2_Display/n5226 [16]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5242 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1884 (
    .a(\u2_Display/n5206 ),
    .b(\u2_Display/n5226 [17]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5241 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1885 (
    .a(\u2_Display/n5205 ),
    .b(\u2_Display/n5226 [18]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5240 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1886 (
    .a(\u2_Display/n5204 ),
    .b(\u2_Display/n5226 [19]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5239 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1887 (
    .a(\u2_Display/n5203 ),
    .b(\u2_Display/n5226 [20]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5238 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1888 (
    .a(\u2_Display/n5202 ),
    .b(\u2_Display/n5226 [21]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5237 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1889 (
    .a(\u2_Display/n5201 ),
    .b(\u2_Display/n5226 [22]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5236 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1890 (
    .a(\u2_Display/n5200 ),
    .b(\u2_Display/n5226 [23]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5235 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1891 (
    .a(\u2_Display/n5199 ),
    .b(\u2_Display/n5226 [24]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5234 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1892 (
    .a(\u2_Display/n5198 ),
    .b(\u2_Display/n5226 [25]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5233 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1893 (
    .a(\u2_Display/n5197 ),
    .b(\u2_Display/n5226 [26]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5232 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1894 (
    .a(\u2_Display/n5196 ),
    .b(\u2_Display/n5226 [27]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5231 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1895 (
    .a(\u2_Display/n6353 ),
    .b(\u2_Display/n5226 [28]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5230 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1896 (
    .a(\u2_Display/n6352 ),
    .b(\u2_Display/n5226 [29]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5229 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1897 (
    .a(\u2_Display/n6351 ),
    .b(\u2_Display/n5226 [30]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5228 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1898 (
    .a(\u2_Display/n6350 ),
    .b(\u2_Display/n5226 [31]),
    .c(\u2_Display/n5224 ),
    .o(\u2_Display/n5227 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1899 (
    .a(\u2_Display/n731 ),
    .b(\u2_Display/n734 [0]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n766 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1900 (
    .a(\u2_Display/n730 ),
    .b(\u2_Display/n734 [1]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n765 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1901 (
    .a(\u2_Display/n729 ),
    .b(\u2_Display/n734 [2]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n764 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1902 (
    .a(\u2_Display/n728 ),
    .b(\u2_Display/n734 [3]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n763 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1903 (
    .a(\u2_Display/n727 ),
    .b(\u2_Display/n734 [4]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n762 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1904 (
    .a(\u2_Display/n726 ),
    .b(\u2_Display/n734 [5]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n761 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1905 (
    .a(\u2_Display/n725 ),
    .b(\u2_Display/n734 [6]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n760 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1906 (
    .a(\u2_Display/n724 ),
    .b(\u2_Display/n734 [7]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n759 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1907 (
    .a(\u2_Display/n723 ),
    .b(\u2_Display/n734 [8]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n758 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1908 (
    .a(\u2_Display/n722 ),
    .b(\u2_Display/n734 [9]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n757 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1909 (
    .a(\u2_Display/n721 ),
    .b(\u2_Display/n734 [10]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n756 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1910 (
    .a(\u2_Display/n720 ),
    .b(\u2_Display/n734 [11]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n755 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1911 (
    .a(\u2_Display/n719 ),
    .b(\u2_Display/n734 [12]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n754 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1912 (
    .a(\u2_Display/n718 ),
    .b(\u2_Display/n734 [13]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n753 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1913 (
    .a(\u2_Display/n717 ),
    .b(\u2_Display/n734 [14]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n752 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1914 (
    .a(\u2_Display/n716 ),
    .b(\u2_Display/n734 [15]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n751 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1915 (
    .a(\u2_Display/n715 ),
    .b(\u2_Display/n734 [16]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n750 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1916 (
    .a(\u2_Display/n714 ),
    .b(\u2_Display/n734 [17]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n749 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1917 (
    .a(\u2_Display/n713 ),
    .b(\u2_Display/n734 [18]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n748 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1918 (
    .a(\u2_Display/n712 ),
    .b(\u2_Display/n734 [19]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n747 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1919 (
    .a(\u2_Display/n711 ),
    .b(\u2_Display/n734 [20]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n746 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1920 (
    .a(\u2_Display/n710 ),
    .b(\u2_Display/n734 [21]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n745 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1921 (
    .a(\u2_Display/n709 ),
    .b(\u2_Display/n734 [22]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n744 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1922 (
    .a(\u2_Display/n708 ),
    .b(\u2_Display/n734 [23]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n743 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1923 (
    .a(\u2_Display/n707 ),
    .b(\u2_Display/n734 [24]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n742 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1924 (
    .a(\u2_Display/n706 ),
    .b(\u2_Display/n734 [25]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n741 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1925 (
    .a(\u2_Display/n705 ),
    .b(\u2_Display/n734 [26]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n740 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1926 (
    .a(\u2_Display/n704 ),
    .b(\u2_Display/n734 [27]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n739 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1927 (
    .a(\u2_Display/n703 ),
    .b(\u2_Display/n734 [28]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n738 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1928 (
    .a(\u2_Display/n702 ),
    .b(\u2_Display/n734 [29]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n737 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1929 (
    .a(\u2_Display/n701 ),
    .b(\u2_Display/n734 [30]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n736 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1930 (
    .a(\u2_Display/n700 ),
    .b(\u2_Display/n734 [31]),
    .c(\u2_Display/n732 ),
    .o(\u2_Display/n735 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1931 (
    .a(\u2_Display/n1854 ),
    .b(\u2_Display/n1857 [0]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1889 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1932 (
    .a(\u2_Display/n1853 ),
    .b(\u2_Display/n1857 [1]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1888 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1933 (
    .a(\u2_Display/n1852 ),
    .b(\u2_Display/n1857 [2]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1887 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1934 (
    .a(\u2_Display/n1851 ),
    .b(\u2_Display/n1857 [3]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1886 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1935 (
    .a(\u2_Display/n1850 ),
    .b(\u2_Display/n1857 [4]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1885 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1936 (
    .a(\u2_Display/n1849 ),
    .b(\u2_Display/n1857 [5]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1884 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1937 (
    .a(\u2_Display/n1848 ),
    .b(\u2_Display/n1857 [6]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1883 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1938 (
    .a(\u2_Display/n1847 ),
    .b(\u2_Display/n1857 [7]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1882 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1939 (
    .a(\u2_Display/n1846 ),
    .b(\u2_Display/n1857 [8]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1881 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1940 (
    .a(\u2_Display/n1845 ),
    .b(\u2_Display/n1857 [9]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1880 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1941 (
    .a(\u2_Display/n1844 ),
    .b(\u2_Display/n1857 [10]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1879 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1942 (
    .a(\u2_Display/n1843 ),
    .b(\u2_Display/n1857 [11]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1878 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1943 (
    .a(\u2_Display/n1842 ),
    .b(\u2_Display/n1857 [12]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1877 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1944 (
    .a(\u2_Display/n1841 ),
    .b(\u2_Display/n1857 [13]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1876 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1945 (
    .a(\u2_Display/n1840 ),
    .b(\u2_Display/n1857 [14]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1875 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1946 (
    .a(\u2_Display/n1839 ),
    .b(\u2_Display/n1857 [15]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1874 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1947 (
    .a(\u2_Display/n1838 ),
    .b(\u2_Display/n1857 [16]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1873 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1948 (
    .a(\u2_Display/n1837 ),
    .b(\u2_Display/n1857 [17]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1872 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1949 (
    .a(\u2_Display/n1836 ),
    .b(\u2_Display/n1857 [18]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1871 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1950 (
    .a(\u2_Display/n1835 ),
    .b(\u2_Display/n1857 [19]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1870 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1951 (
    .a(\u2_Display/n1834 ),
    .b(\u2_Display/n1857 [20]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1869 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1952 (
    .a(\u2_Display/n1833 ),
    .b(\u2_Display/n1857 [21]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1868 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1953 (
    .a(\u2_Display/n1832 ),
    .b(\u2_Display/n1857 [22]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1867 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1954 (
    .a(\u2_Display/n1831 ),
    .b(\u2_Display/n1857 [23]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1866 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1955 (
    .a(\u2_Display/n1830 ),
    .b(\u2_Display/n1857 [24]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1865 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1956 (
    .a(\u2_Display/n1829 ),
    .b(\u2_Display/n1857 [25]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1864 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1957 (
    .a(\u2_Display/n1828 ),
    .b(\u2_Display/n1857 [26]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1863 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1958 (
    .a(\u2_Display/n1827 ),
    .b(\u2_Display/n1857 [27]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1862 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1959 (
    .a(\u2_Display/n1826 ),
    .b(\u2_Display/n1857 [28]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1861 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1960 (
    .a(\u2_Display/n1825 ),
    .b(\u2_Display/n1857 [29]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1860 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1961 (
    .a(\u2_Display/n1824 ),
    .b(\u2_Display/n1857 [30]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1859 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1962 (
    .a(\u2_Display/n1823 ),
    .b(\u2_Display/n1857 [31]),
    .c(\u2_Display/n1855 ),
    .o(\u2_Display/n1858 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1963 (
    .a(\u2_Display/n2977 ),
    .b(\u2_Display/n2980 [0]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3012 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1964 (
    .a(\u2_Display/n2976 ),
    .b(\u2_Display/n2980 [1]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3011 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1965 (
    .a(\u2_Display/n2975 ),
    .b(\u2_Display/n2980 [2]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3010 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1966 (
    .a(\u2_Display/n2974 ),
    .b(\u2_Display/n2980 [3]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3009 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1967 (
    .a(\u2_Display/n2973 ),
    .b(\u2_Display/n2980 [4]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3008 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1968 (
    .a(\u2_Display/n2972 ),
    .b(\u2_Display/n2980 [5]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3007 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1969 (
    .a(\u2_Display/n2971 ),
    .b(\u2_Display/n2980 [6]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3006 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1970 (
    .a(\u2_Display/n2970 ),
    .b(\u2_Display/n2980 [7]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3005 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1971 (
    .a(\u2_Display/n2969 ),
    .b(\u2_Display/n2980 [8]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3004 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1972 (
    .a(\u2_Display/n2968 ),
    .b(\u2_Display/n2980 [9]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3003 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1973 (
    .a(\u2_Display/n2967 ),
    .b(\u2_Display/n2980 [10]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3002 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1974 (
    .a(\u2_Display/n2966 ),
    .b(\u2_Display/n2980 [11]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3001 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1975 (
    .a(\u2_Display/n2965 ),
    .b(\u2_Display/n2980 [12]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n3000 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1976 (
    .a(\u2_Display/n2964 ),
    .b(\u2_Display/n2980 [13]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2999 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1977 (
    .a(\u2_Display/n2963 ),
    .b(\u2_Display/n2980 [14]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2998 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1978 (
    .a(\u2_Display/n2962 ),
    .b(\u2_Display/n2980 [15]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2997 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1979 (
    .a(\u2_Display/n2961 ),
    .b(\u2_Display/n2980 [16]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2996 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1980 (
    .a(\u2_Display/n2960 ),
    .b(\u2_Display/n2980 [17]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2995 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1981 (
    .a(\u2_Display/n2959 ),
    .b(\u2_Display/n2980 [18]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2994 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1982 (
    .a(\u2_Display/n2958 ),
    .b(\u2_Display/n2980 [19]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2993 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1983 (
    .a(\u2_Display/n2957 ),
    .b(\u2_Display/n2980 [20]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2992 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1984 (
    .a(\u2_Display/n2956 ),
    .b(\u2_Display/n2980 [21]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2991 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1985 (
    .a(\u2_Display/n2955 ),
    .b(\u2_Display/n2980 [22]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2990 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1986 (
    .a(\u2_Display/n2954 ),
    .b(\u2_Display/n2980 [23]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2989 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1987 (
    .a(\u2_Display/n2953 ),
    .b(\u2_Display/n2980 [24]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2988 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1988 (
    .a(\u2_Display/n2952 ),
    .b(\u2_Display/n2980 [25]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2987 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1989 (
    .a(\u2_Display/n2951 ),
    .b(\u2_Display/n2980 [26]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2986 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1990 (
    .a(\u2_Display/n2950 ),
    .b(\u2_Display/n2980 [27]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2985 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1991 (
    .a(\u2_Display/n2949 ),
    .b(\u2_Display/n2980 [28]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2984 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1992 (
    .a(\u2_Display/n2948 ),
    .b(\u2_Display/n2980 [29]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2983 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1993 (
    .a(\u2_Display/n2947 ),
    .b(\u2_Display/n2980 [30]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2982 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1994 (
    .a(\u2_Display/n2946 ),
    .b(\u2_Display/n2980 [31]),
    .c(\u2_Display/n2978 ),
    .o(\u2_Display/n2981 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1995 (
    .a(\u2_Display/n4135 ),
    .b(\u2_Display/n4138 [0]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4170 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1996 (
    .a(\u2_Display/n4134 ),
    .b(\u2_Display/n4138 [1]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4169 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1997 (
    .a(\u2_Display/n4133 ),
    .b(\u2_Display/n4138 [2]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4168 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1998 (
    .a(\u2_Display/n4132 ),
    .b(\u2_Display/n4138 [3]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4167 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1999 (
    .a(\u2_Display/n4131 ),
    .b(\u2_Display/n4138 [4]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4166 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2000 (
    .a(\u2_Display/n4130 ),
    .b(\u2_Display/n4138 [5]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4165 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2001 (
    .a(\u2_Display/n4129 ),
    .b(\u2_Display/n4138 [6]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4164 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2002 (
    .a(\u2_Display/n4128 ),
    .b(\u2_Display/n4138 [7]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4163 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2003 (
    .a(\u2_Display/n4127 ),
    .b(\u2_Display/n4138 [8]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4162 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2004 (
    .a(\u2_Display/n4126 ),
    .b(\u2_Display/n4138 [9]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4161 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2005 (
    .a(\u2_Display/n4125 ),
    .b(\u2_Display/n4138 [10]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4160 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2006 (
    .a(\u2_Display/n4124 ),
    .b(\u2_Display/n4138 [11]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4159 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2007 (
    .a(\u2_Display/n4123 ),
    .b(\u2_Display/n4138 [12]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4158 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2008 (
    .a(\u2_Display/n4122 ),
    .b(\u2_Display/n4138 [13]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4157 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2009 (
    .a(\u2_Display/n4121 ),
    .b(\u2_Display/n4138 [14]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4156 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2010 (
    .a(\u2_Display/n4120 ),
    .b(\u2_Display/n4138 [15]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4155 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2011 (
    .a(\u2_Display/n4119 ),
    .b(\u2_Display/n4138 [16]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4154 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2012 (
    .a(\u2_Display/n4118 ),
    .b(\u2_Display/n4138 [17]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4153 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2013 (
    .a(\u2_Display/n4117 ),
    .b(\u2_Display/n4138 [18]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4152 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2014 (
    .a(\u2_Display/n4116 ),
    .b(\u2_Display/n4138 [19]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4151 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2015 (
    .a(\u2_Display/n4115 ),
    .b(\u2_Display/n4138 [20]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4150 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2016 (
    .a(\u2_Display/n4114 ),
    .b(\u2_Display/n4138 [21]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4149 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2017 (
    .a(\u2_Display/n4113 ),
    .b(\u2_Display/n4138 [22]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4148 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2018 (
    .a(\u2_Display/n4112 ),
    .b(\u2_Display/n4138 [23]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4147 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2019 (
    .a(\u2_Display/n4111 ),
    .b(\u2_Display/n4138 [24]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4146 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2020 (
    .a(\u2_Display/n4110 ),
    .b(\u2_Display/n4138 [25]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4145 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2021 (
    .a(\u2_Display/n4109 ),
    .b(\u2_Display/n4138 [26]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4144 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2022 (
    .a(\u2_Display/n4108 ),
    .b(\u2_Display/n4138 [27]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4143 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2023 (
    .a(\u2_Display/n4107 ),
    .b(\u2_Display/n4138 [28]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4142 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2024 (
    .a(\u2_Display/n4106 ),
    .b(\u2_Display/n4138 [29]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4141 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2025 (
    .a(\u2_Display/n4105 ),
    .b(\u2_Display/n4138 [30]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4140 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2026 (
    .a(\u2_Display/n4104 ),
    .b(\u2_Display/n4138 [31]),
    .c(\u2_Display/n4136 ),
    .o(\u2_Display/n4139 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2027 (
    .a(\u2_Display/n5258 ),
    .b(\u2_Display/n5261 [0]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5293 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2028 (
    .a(\u2_Display/n5257 ),
    .b(\u2_Display/n5261 [1]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5292 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2029 (
    .a(\u2_Display/n5256 ),
    .b(\u2_Display/n5261 [2]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5291 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2030 (
    .a(\u2_Display/n5255 ),
    .b(\u2_Display/n5261 [3]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5290 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2031 (
    .a(\u2_Display/n5254 ),
    .b(\u2_Display/n5261 [4]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5289 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2032 (
    .a(\u2_Display/n5253 ),
    .b(\u2_Display/n5261 [5]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5288 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2033 (
    .a(\u2_Display/n5252 ),
    .b(\u2_Display/n5261 [6]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5287 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2034 (
    .a(\u2_Display/n5251 ),
    .b(\u2_Display/n5261 [7]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5286 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2035 (
    .a(\u2_Display/n5250 ),
    .b(\u2_Display/n5261 [8]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5285 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2036 (
    .a(\u2_Display/n5249 ),
    .b(\u2_Display/n5261 [9]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5284 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2037 (
    .a(\u2_Display/n5248 ),
    .b(\u2_Display/n5261 [10]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5283 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2038 (
    .a(\u2_Display/n5247 ),
    .b(\u2_Display/n5261 [11]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5282 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2039 (
    .a(\u2_Display/n5246 ),
    .b(\u2_Display/n5261 [12]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5281 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2040 (
    .a(\u2_Display/n5245 ),
    .b(\u2_Display/n5261 [13]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5280 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2041 (
    .a(\u2_Display/n5244 ),
    .b(\u2_Display/n5261 [14]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5279 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2042 (
    .a(\u2_Display/n5243 ),
    .b(\u2_Display/n5261 [15]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5278 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2043 (
    .a(\u2_Display/n5242 ),
    .b(\u2_Display/n5261 [16]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5277 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2044 (
    .a(\u2_Display/n5241 ),
    .b(\u2_Display/n5261 [17]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5276 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2045 (
    .a(\u2_Display/n5240 ),
    .b(\u2_Display/n5261 [18]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5275 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2046 (
    .a(\u2_Display/n5239 ),
    .b(\u2_Display/n5261 [19]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5274 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2047 (
    .a(\u2_Display/n5238 ),
    .b(\u2_Display/n5261 [20]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5273 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2048 (
    .a(\u2_Display/n5237 ),
    .b(\u2_Display/n5261 [21]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5272 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2049 (
    .a(\u2_Display/n5236 ),
    .b(\u2_Display/n5261 [22]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5271 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2050 (
    .a(\u2_Display/n5235 ),
    .b(\u2_Display/n5261 [23]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5270 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2051 (
    .a(\u2_Display/n5234 ),
    .b(\u2_Display/n5261 [24]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5269 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2052 (
    .a(\u2_Display/n5233 ),
    .b(\u2_Display/n5261 [25]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5268 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2053 (
    .a(\u2_Display/n5232 ),
    .b(\u2_Display/n5261 [26]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5267 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2054 (
    .a(\u2_Display/n5231 ),
    .b(\u2_Display/n5261 [27]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5266 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2055 (
    .a(\u2_Display/n5230 ),
    .b(\u2_Display/n5261 [28]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5265 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2056 (
    .a(\u2_Display/n5229 ),
    .b(\u2_Display/n5261 [29]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5264 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2057 (
    .a(\u2_Display/n5228 ),
    .b(\u2_Display/n5261 [30]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5263 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2058 (
    .a(\u2_Display/n5227 ),
    .b(\u2_Display/n5261 [31]),
    .c(\u2_Display/n5259 ),
    .o(\u2_Display/n5262 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2059 (
    .a(\u2_Display/n766 ),
    .b(\u2_Display/n769 [0]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n801 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2060 (
    .a(\u2_Display/n765 ),
    .b(\u2_Display/n769 [1]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n800 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2061 (
    .a(\u2_Display/n764 ),
    .b(\u2_Display/n769 [2]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n799 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2062 (
    .a(\u2_Display/n763 ),
    .b(\u2_Display/n769 [3]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n798 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2063 (
    .a(\u2_Display/n762 ),
    .b(\u2_Display/n769 [4]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n797 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2064 (
    .a(\u2_Display/n761 ),
    .b(\u2_Display/n769 [5]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n796 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2065 (
    .a(\u2_Display/n760 ),
    .b(\u2_Display/n769 [6]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n795 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2066 (
    .a(\u2_Display/n759 ),
    .b(\u2_Display/n769 [7]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n794 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2067 (
    .a(\u2_Display/n758 ),
    .b(\u2_Display/n769 [8]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n793 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2068 (
    .a(\u2_Display/n757 ),
    .b(\u2_Display/n769 [9]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n792 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2069 (
    .a(\u2_Display/n756 ),
    .b(\u2_Display/n769 [10]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n791 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2070 (
    .a(\u2_Display/n755 ),
    .b(\u2_Display/n769 [11]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n790 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2071 (
    .a(\u2_Display/n754 ),
    .b(\u2_Display/n769 [12]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n789 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2072 (
    .a(\u2_Display/n753 ),
    .b(\u2_Display/n769 [13]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n788 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2073 (
    .a(\u2_Display/n752 ),
    .b(\u2_Display/n769 [14]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n787 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2074 (
    .a(\u2_Display/n751 ),
    .b(\u2_Display/n769 [15]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n786 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2075 (
    .a(\u2_Display/n750 ),
    .b(\u2_Display/n769 [16]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n785 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2076 (
    .a(\u2_Display/n749 ),
    .b(\u2_Display/n769 [17]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n784 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2077 (
    .a(\u2_Display/n748 ),
    .b(\u2_Display/n769 [18]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n783 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2078 (
    .a(\u2_Display/n747 ),
    .b(\u2_Display/n769 [19]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n782 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2079 (
    .a(\u2_Display/n746 ),
    .b(\u2_Display/n769 [20]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n781 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2080 (
    .a(\u2_Display/n745 ),
    .b(\u2_Display/n769 [21]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n780 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2081 (
    .a(\u2_Display/n744 ),
    .b(\u2_Display/n769 [22]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n779 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2082 (
    .a(\u2_Display/n743 ),
    .b(\u2_Display/n769 [23]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n778 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2083 (
    .a(\u2_Display/n742 ),
    .b(\u2_Display/n769 [24]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n777 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2084 (
    .a(\u2_Display/n741 ),
    .b(\u2_Display/n769 [25]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n776 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2085 (
    .a(\u2_Display/n740 ),
    .b(\u2_Display/n769 [26]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n775 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2086 (
    .a(\u2_Display/n739 ),
    .b(\u2_Display/n769 [27]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n774 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2087 (
    .a(\u2_Display/n738 ),
    .b(\u2_Display/n769 [28]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n773 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2088 (
    .a(\u2_Display/n737 ),
    .b(\u2_Display/n769 [29]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n772 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2089 (
    .a(\u2_Display/n736 ),
    .b(\u2_Display/n769 [30]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n771 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2090 (
    .a(\u2_Display/n735 ),
    .b(\u2_Display/n769 [31]),
    .c(\u2_Display/n767 ),
    .o(\u2_Display/n770 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2091 (
    .a(\u2_Display/n1889 ),
    .b(\u2_Display/n1892 [0]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1924 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2092 (
    .a(\u2_Display/n1888 ),
    .b(\u2_Display/n1892 [1]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1923 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2093 (
    .a(\u2_Display/n1887 ),
    .b(\u2_Display/n1892 [2]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1922 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2094 (
    .a(\u2_Display/n1886 ),
    .b(\u2_Display/n1892 [3]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1921 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2095 (
    .a(\u2_Display/n1885 ),
    .b(\u2_Display/n1892 [4]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1920 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2096 (
    .a(\u2_Display/n1884 ),
    .b(\u2_Display/n1892 [5]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1919 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2097 (
    .a(\u2_Display/n1883 ),
    .b(\u2_Display/n1892 [6]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1918 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2098 (
    .a(\u2_Display/n1882 ),
    .b(\u2_Display/n1892 [7]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1917 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2099 (
    .a(\u2_Display/n1881 ),
    .b(\u2_Display/n1892 [8]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1916 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2100 (
    .a(\u2_Display/n1880 ),
    .b(\u2_Display/n1892 [9]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1915 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2101 (
    .a(\u2_Display/n1879 ),
    .b(\u2_Display/n1892 [10]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1914 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2102 (
    .a(\u2_Display/n1878 ),
    .b(\u2_Display/n1892 [11]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1913 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2103 (
    .a(\u2_Display/n1877 ),
    .b(\u2_Display/n1892 [12]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1912 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2104 (
    .a(\u2_Display/n1876 ),
    .b(\u2_Display/n1892 [13]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1911 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2105 (
    .a(\u2_Display/n1875 ),
    .b(\u2_Display/n1892 [14]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1910 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2106 (
    .a(\u2_Display/n1874 ),
    .b(\u2_Display/n1892 [15]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1909 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2107 (
    .a(\u2_Display/n1873 ),
    .b(\u2_Display/n1892 [16]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1908 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2108 (
    .a(\u2_Display/n1872 ),
    .b(\u2_Display/n1892 [17]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1907 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2109 (
    .a(\u2_Display/n1871 ),
    .b(\u2_Display/n1892 [18]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1906 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2110 (
    .a(\u2_Display/n1870 ),
    .b(\u2_Display/n1892 [19]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1905 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2111 (
    .a(\u2_Display/n1869 ),
    .b(\u2_Display/n1892 [20]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1904 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2112 (
    .a(\u2_Display/n1868 ),
    .b(\u2_Display/n1892 [21]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1903 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2113 (
    .a(\u2_Display/n1867 ),
    .b(\u2_Display/n1892 [22]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1902 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2114 (
    .a(\u2_Display/n1866 ),
    .b(\u2_Display/n1892 [23]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1901 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2115 (
    .a(\u2_Display/n1865 ),
    .b(\u2_Display/n1892 [24]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1900 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2116 (
    .a(\u2_Display/n1864 ),
    .b(\u2_Display/n1892 [25]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1899 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2117 (
    .a(\u2_Display/n1863 ),
    .b(\u2_Display/n1892 [26]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1898 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2118 (
    .a(\u2_Display/n1862 ),
    .b(\u2_Display/n1892 [27]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1897 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2119 (
    .a(\u2_Display/n1861 ),
    .b(\u2_Display/n1892 [28]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1896 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2120 (
    .a(\u2_Display/n1860 ),
    .b(\u2_Display/n1892 [29]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1895 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2121 (
    .a(\u2_Display/n1859 ),
    .b(\u2_Display/n1892 [30]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1894 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2122 (
    .a(\u2_Display/n1858 ),
    .b(\u2_Display/n1892 [31]),
    .c(\u2_Display/n1890 ),
    .o(\u2_Display/n1893 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2123 (
    .a(\u2_Display/n3012 ),
    .b(\u2_Display/n3015 [0]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3047 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2124 (
    .a(\u2_Display/n3011 ),
    .b(\u2_Display/n3015 [1]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3046 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2125 (
    .a(\u2_Display/n3010 ),
    .b(\u2_Display/n3015 [2]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3045 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2126 (
    .a(\u2_Display/n3009 ),
    .b(\u2_Display/n3015 [3]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3044 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2127 (
    .a(\u2_Display/n3008 ),
    .b(\u2_Display/n3015 [4]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3043 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2128 (
    .a(\u2_Display/n3007 ),
    .b(\u2_Display/n3015 [5]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3042 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2129 (
    .a(\u2_Display/n3006 ),
    .b(\u2_Display/n3015 [6]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3041 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2130 (
    .a(\u2_Display/n3005 ),
    .b(\u2_Display/n3015 [7]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3040 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2131 (
    .a(\u2_Display/n3004 ),
    .b(\u2_Display/n3015 [8]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3039 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2132 (
    .a(\u2_Display/n3003 ),
    .b(\u2_Display/n3015 [9]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3038 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2133 (
    .a(\u2_Display/n3002 ),
    .b(\u2_Display/n3015 [10]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3037 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2134 (
    .a(\u2_Display/n3001 ),
    .b(\u2_Display/n3015 [11]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3036 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2135 (
    .a(\u2_Display/n3000 ),
    .b(\u2_Display/n3015 [12]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3035 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2136 (
    .a(\u2_Display/n2999 ),
    .b(\u2_Display/n3015 [13]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3034 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2137 (
    .a(\u2_Display/n2998 ),
    .b(\u2_Display/n3015 [14]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3033 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2138 (
    .a(\u2_Display/n2997 ),
    .b(\u2_Display/n3015 [15]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3032 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2139 (
    .a(\u2_Display/n2996 ),
    .b(\u2_Display/n3015 [16]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3031 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2140 (
    .a(\u2_Display/n2995 ),
    .b(\u2_Display/n3015 [17]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3030 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2141 (
    .a(\u2_Display/n2994 ),
    .b(\u2_Display/n3015 [18]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3029 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2142 (
    .a(\u2_Display/n2993 ),
    .b(\u2_Display/n3015 [19]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3028 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2143 (
    .a(\u2_Display/n2992 ),
    .b(\u2_Display/n3015 [20]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3027 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2144 (
    .a(\u2_Display/n2991 ),
    .b(\u2_Display/n3015 [21]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3026 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2145 (
    .a(\u2_Display/n2990 ),
    .b(\u2_Display/n3015 [22]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3025 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2146 (
    .a(\u2_Display/n2989 ),
    .b(\u2_Display/n3015 [23]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3024 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2147 (
    .a(\u2_Display/n2988 ),
    .b(\u2_Display/n3015 [24]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3023 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2148 (
    .a(\u2_Display/n2987 ),
    .b(\u2_Display/n3015 [25]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3022 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2149 (
    .a(\u2_Display/n2986 ),
    .b(\u2_Display/n3015 [26]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3021 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2150 (
    .a(\u2_Display/n2985 ),
    .b(\u2_Display/n3015 [27]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3020 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2151 (
    .a(\u2_Display/n2984 ),
    .b(\u2_Display/n3015 [28]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3019 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2152 (
    .a(\u2_Display/n2983 ),
    .b(\u2_Display/n3015 [29]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3018 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2153 (
    .a(\u2_Display/n2982 ),
    .b(\u2_Display/n3015 [30]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3017 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2154 (
    .a(\u2_Display/n2981 ),
    .b(\u2_Display/n3015 [31]),
    .c(\u2_Display/n3013 ),
    .o(\u2_Display/n3016 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2155 (
    .a(\u2_Display/n4170 ),
    .b(\u2_Display/n4173 [0]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4205 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2156 (
    .a(\u2_Display/n4169 ),
    .b(\u2_Display/n4173 [1]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4204 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2157 (
    .a(\u2_Display/n4168 ),
    .b(\u2_Display/n4173 [2]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4203 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2158 (
    .a(\u2_Display/n4167 ),
    .b(\u2_Display/n4173 [3]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4202 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2159 (
    .a(\u2_Display/n4166 ),
    .b(\u2_Display/n4173 [4]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4201 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2160 (
    .a(\u2_Display/n4165 ),
    .b(\u2_Display/n4173 [5]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4200 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2161 (
    .a(\u2_Display/n4164 ),
    .b(\u2_Display/n4173 [6]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4199 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2162 (
    .a(\u2_Display/n4163 ),
    .b(\u2_Display/n4173 [7]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4198 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2163 (
    .a(\u2_Display/n4162 ),
    .b(\u2_Display/n4173 [8]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4197 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2164 (
    .a(\u2_Display/n4161 ),
    .b(\u2_Display/n4173 [9]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4196 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2165 (
    .a(\u2_Display/n4160 ),
    .b(\u2_Display/n4173 [10]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4195 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2166 (
    .a(\u2_Display/n4159 ),
    .b(\u2_Display/n4173 [11]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4194 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2167 (
    .a(\u2_Display/n4158 ),
    .b(\u2_Display/n4173 [12]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4193 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2168 (
    .a(\u2_Display/n4157 ),
    .b(\u2_Display/n4173 [13]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4192 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2169 (
    .a(\u2_Display/n4156 ),
    .b(\u2_Display/n4173 [14]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4191 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2170 (
    .a(\u2_Display/n4155 ),
    .b(\u2_Display/n4173 [15]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4190 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2171 (
    .a(\u2_Display/n4154 ),
    .b(\u2_Display/n4173 [16]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4189 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2172 (
    .a(\u2_Display/n4153 ),
    .b(\u2_Display/n4173 [17]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4188 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2173 (
    .a(\u2_Display/n4152 ),
    .b(\u2_Display/n4173 [18]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4187 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2174 (
    .a(\u2_Display/n4151 ),
    .b(\u2_Display/n4173 [19]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4186 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2175 (
    .a(\u2_Display/n4150 ),
    .b(\u2_Display/n4173 [20]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4185 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2176 (
    .a(\u2_Display/n4149 ),
    .b(\u2_Display/n4173 [21]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4184 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2177 (
    .a(\u2_Display/n4148 ),
    .b(\u2_Display/n4173 [22]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4183 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2178 (
    .a(\u2_Display/n4147 ),
    .b(\u2_Display/n4173 [23]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4182 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2179 (
    .a(\u2_Display/n4146 ),
    .b(\u2_Display/n4173 [24]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4181 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2180 (
    .a(\u2_Display/n4145 ),
    .b(\u2_Display/n4173 [25]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4180 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2181 (
    .a(\u2_Display/n4144 ),
    .b(\u2_Display/n4173 [26]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4179 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2182 (
    .a(\u2_Display/n4143 ),
    .b(\u2_Display/n4173 [27]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4178 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2183 (
    .a(\u2_Display/n4142 ),
    .b(\u2_Display/n4173 [28]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4177 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2184 (
    .a(\u2_Display/n4141 ),
    .b(\u2_Display/n4173 [29]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4176 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2185 (
    .a(\u2_Display/n4140 ),
    .b(\u2_Display/n4173 [30]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4175 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2186 (
    .a(\u2_Display/n4139 ),
    .b(\u2_Display/n4173 [31]),
    .c(\u2_Display/n4171 ),
    .o(\u2_Display/n4174 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2187 (
    .a(\u2_Display/n5293 ),
    .b(\u2_Display/n5296 [0]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5328 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2188 (
    .a(\u2_Display/n5292 ),
    .b(\u2_Display/n5296 [1]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5327 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2189 (
    .a(\u2_Display/n5291 ),
    .b(\u2_Display/n5296 [2]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5326 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2190 (
    .a(\u2_Display/n5290 ),
    .b(\u2_Display/n5296 [3]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5325 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2191 (
    .a(\u2_Display/n5289 ),
    .b(\u2_Display/n5296 [4]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5324 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2192 (
    .a(\u2_Display/n5288 ),
    .b(\u2_Display/n5296 [5]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5323 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2193 (
    .a(\u2_Display/n5287 ),
    .b(\u2_Display/n5296 [6]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5322 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2194 (
    .a(\u2_Display/n5286 ),
    .b(\u2_Display/n5296 [7]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5321 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2195 (
    .a(\u2_Display/n5285 ),
    .b(\u2_Display/n5296 [8]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5320 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2196 (
    .a(\u2_Display/n5284 ),
    .b(\u2_Display/n5296 [9]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5319 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2197 (
    .a(\u2_Display/n5283 ),
    .b(\u2_Display/n5296 [10]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5318 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2198 (
    .a(\u2_Display/n5282 ),
    .b(\u2_Display/n5296 [11]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5317 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2199 (
    .a(\u2_Display/n5281 ),
    .b(\u2_Display/n5296 [12]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5316 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2200 (
    .a(\u2_Display/n5280 ),
    .b(\u2_Display/n5296 [13]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5315 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2201 (
    .a(\u2_Display/n5279 ),
    .b(\u2_Display/n5296 [14]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5314 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2202 (
    .a(\u2_Display/n5278 ),
    .b(\u2_Display/n5296 [15]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5313 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2203 (
    .a(\u2_Display/n5277 ),
    .b(\u2_Display/n5296 [16]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5312 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2204 (
    .a(\u2_Display/n5276 ),
    .b(\u2_Display/n5296 [17]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5311 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2205 (
    .a(\u2_Display/n5275 ),
    .b(\u2_Display/n5296 [18]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5310 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2206 (
    .a(\u2_Display/n5274 ),
    .b(\u2_Display/n5296 [19]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5309 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2207 (
    .a(\u2_Display/n5273 ),
    .b(\u2_Display/n5296 [20]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5308 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2208 (
    .a(\u2_Display/n5272 ),
    .b(\u2_Display/n5296 [21]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5307 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2209 (
    .a(\u2_Display/n5271 ),
    .b(\u2_Display/n5296 [22]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5306 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2210 (
    .a(\u2_Display/n5270 ),
    .b(\u2_Display/n5296 [23]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5305 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2211 (
    .a(\u2_Display/n5269 ),
    .b(\u2_Display/n5296 [24]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5304 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2212 (
    .a(\u2_Display/n5268 ),
    .b(\u2_Display/n5296 [25]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5303 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2213 (
    .a(\u2_Display/n5267 ),
    .b(\u2_Display/n5296 [26]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5302 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2214 (
    .a(\u2_Display/n5266 ),
    .b(\u2_Display/n5296 [27]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5301 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2215 (
    .a(\u2_Display/n5265 ),
    .b(\u2_Display/n5296 [28]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5300 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2216 (
    .a(\u2_Display/n5264 ),
    .b(\u2_Display/n5296 [29]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5299 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2217 (
    .a(\u2_Display/n5263 ),
    .b(\u2_Display/n5296 [30]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5298 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2218 (
    .a(\u2_Display/n5262 ),
    .b(\u2_Display/n5296 [31]),
    .c(\u2_Display/n5294 ),
    .o(\u2_Display/n5297 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2219 (
    .a(\u2_Display/n801 ),
    .b(\u2_Display/n804 [0]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n836 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2220 (
    .a(\u2_Display/n800 ),
    .b(\u2_Display/n804 [1]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n835 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2221 (
    .a(\u2_Display/n799 ),
    .b(\u2_Display/n804 [2]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n834 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2222 (
    .a(\u2_Display/n798 ),
    .b(\u2_Display/n804 [3]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n833 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2223 (
    .a(\u2_Display/n797 ),
    .b(\u2_Display/n804 [4]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n832 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2224 (
    .a(\u2_Display/n796 ),
    .b(\u2_Display/n804 [5]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n831 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2225 (
    .a(\u2_Display/n795 ),
    .b(\u2_Display/n804 [6]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n830 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2226 (
    .a(\u2_Display/n794 ),
    .b(\u2_Display/n804 [7]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n829 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2227 (
    .a(\u2_Display/n793 ),
    .b(\u2_Display/n804 [8]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n828 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2228 (
    .a(\u2_Display/n792 ),
    .b(\u2_Display/n804 [9]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n827 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2229 (
    .a(\u2_Display/n791 ),
    .b(\u2_Display/n804 [10]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n826 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2230 (
    .a(\u2_Display/n790 ),
    .b(\u2_Display/n804 [11]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n825 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2231 (
    .a(\u2_Display/n789 ),
    .b(\u2_Display/n804 [12]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n824 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2232 (
    .a(\u2_Display/n788 ),
    .b(\u2_Display/n804 [13]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n823 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2233 (
    .a(\u2_Display/n787 ),
    .b(\u2_Display/n804 [14]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n822 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2234 (
    .a(\u2_Display/n786 ),
    .b(\u2_Display/n804 [15]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n821 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2235 (
    .a(\u2_Display/n785 ),
    .b(\u2_Display/n804 [16]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n820 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2236 (
    .a(\u2_Display/n784 ),
    .b(\u2_Display/n804 [17]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n819 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2237 (
    .a(\u2_Display/n783 ),
    .b(\u2_Display/n804 [18]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n818 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2238 (
    .a(\u2_Display/n782 ),
    .b(\u2_Display/n804 [19]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n817 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2239 (
    .a(\u2_Display/n781 ),
    .b(\u2_Display/n804 [20]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n816 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2240 (
    .a(\u2_Display/n780 ),
    .b(\u2_Display/n804 [21]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n815 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2241 (
    .a(\u2_Display/n779 ),
    .b(\u2_Display/n804 [22]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n814 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2242 (
    .a(\u2_Display/n778 ),
    .b(\u2_Display/n804 [23]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n813 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2243 (
    .a(\u2_Display/n777 ),
    .b(\u2_Display/n804 [24]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n812 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2244 (
    .a(\u2_Display/n776 ),
    .b(\u2_Display/n804 [25]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n811 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2245 (
    .a(\u2_Display/n775 ),
    .b(\u2_Display/n804 [26]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n810 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2246 (
    .a(\u2_Display/n774 ),
    .b(\u2_Display/n804 [27]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n809 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2247 (
    .a(\u2_Display/n773 ),
    .b(\u2_Display/n804 [28]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n808 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2248 (
    .a(\u2_Display/n772 ),
    .b(\u2_Display/n804 [29]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n807 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2249 (
    .a(\u2_Display/n771 ),
    .b(\u2_Display/n804 [30]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n806 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2250 (
    .a(\u2_Display/n770 ),
    .b(\u2_Display/n804 [31]),
    .c(\u2_Display/n802 ),
    .o(\u2_Display/n805 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2251 (
    .a(\u2_Display/n1924 ),
    .b(\u2_Display/n1927 [0]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1959 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2252 (
    .a(\u2_Display/n1923 ),
    .b(\u2_Display/n1927 [1]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1958 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2253 (
    .a(\u2_Display/n1922 ),
    .b(\u2_Display/n1927 [2]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1957 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2254 (
    .a(\u2_Display/n1921 ),
    .b(\u2_Display/n1927 [3]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1956 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2255 (
    .a(\u2_Display/n1920 ),
    .b(\u2_Display/n1927 [4]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1955 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2256 (
    .a(\u2_Display/n1919 ),
    .b(\u2_Display/n1927 [5]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1954 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2257 (
    .a(\u2_Display/n1918 ),
    .b(\u2_Display/n1927 [6]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1953 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2258 (
    .a(\u2_Display/n1917 ),
    .b(\u2_Display/n1927 [7]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1952 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2259 (
    .a(\u2_Display/n1916 ),
    .b(\u2_Display/n1927 [8]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1951 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2260 (
    .a(\u2_Display/n1915 ),
    .b(\u2_Display/n1927 [9]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1950 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2261 (
    .a(\u2_Display/n1914 ),
    .b(\u2_Display/n1927 [10]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1949 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2262 (
    .a(\u2_Display/n1913 ),
    .b(\u2_Display/n1927 [11]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1948 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2263 (
    .a(\u2_Display/n1912 ),
    .b(\u2_Display/n1927 [12]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1947 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2264 (
    .a(\u2_Display/n1911 ),
    .b(\u2_Display/n1927 [13]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1946 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2265 (
    .a(\u2_Display/n1910 ),
    .b(\u2_Display/n1927 [14]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1945 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2266 (
    .a(\u2_Display/n1909 ),
    .b(\u2_Display/n1927 [15]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1944 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2267 (
    .a(\u2_Display/n1908 ),
    .b(\u2_Display/n1927 [16]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1943 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2268 (
    .a(\u2_Display/n1907 ),
    .b(\u2_Display/n1927 [17]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1942 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2269 (
    .a(\u2_Display/n1906 ),
    .b(\u2_Display/n1927 [18]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1941 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2270 (
    .a(\u2_Display/n1905 ),
    .b(\u2_Display/n1927 [19]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1940 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2271 (
    .a(\u2_Display/n1904 ),
    .b(\u2_Display/n1927 [20]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1939 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2272 (
    .a(\u2_Display/n1903 ),
    .b(\u2_Display/n1927 [21]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1938 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2273 (
    .a(\u2_Display/n1902 ),
    .b(\u2_Display/n1927 [22]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1937 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2274 (
    .a(\u2_Display/n1901 ),
    .b(\u2_Display/n1927 [23]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1936 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2275 (
    .a(\u2_Display/n1900 ),
    .b(\u2_Display/n1927 [24]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1935 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2276 (
    .a(\u2_Display/n1899 ),
    .b(\u2_Display/n1927 [25]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1934 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2277 (
    .a(\u2_Display/n1898 ),
    .b(\u2_Display/n1927 [26]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1933 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2278 (
    .a(\u2_Display/n1897 ),
    .b(\u2_Display/n1927 [27]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1932 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2279 (
    .a(\u2_Display/n1896 ),
    .b(\u2_Display/n1927 [28]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1931 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2280 (
    .a(\u2_Display/n1895 ),
    .b(\u2_Display/n1927 [29]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1930 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2281 (
    .a(\u2_Display/n1894 ),
    .b(\u2_Display/n1927 [30]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1929 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2282 (
    .a(\u2_Display/n1893 ),
    .b(\u2_Display/n1927 [31]),
    .c(\u2_Display/n1925 ),
    .o(\u2_Display/n1928 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2283 (
    .a(\u2_Display/n3047 ),
    .b(\u2_Display/n3050 [0]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3082 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2284 (
    .a(\u2_Display/n3046 ),
    .b(\u2_Display/n3050 [1]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3081 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2285 (
    .a(\u2_Display/n3045 ),
    .b(\u2_Display/n3050 [2]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3080 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2286 (
    .a(\u2_Display/n3044 ),
    .b(\u2_Display/n3050 [3]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3079 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2287 (
    .a(\u2_Display/n3043 ),
    .b(\u2_Display/n3050 [4]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3078 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2288 (
    .a(\u2_Display/n3042 ),
    .b(\u2_Display/n3050 [5]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3077 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2289 (
    .a(\u2_Display/n3041 ),
    .b(\u2_Display/n3050 [6]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3076 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2290 (
    .a(\u2_Display/n3040 ),
    .b(\u2_Display/n3050 [7]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3075 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2291 (
    .a(\u2_Display/n3039 ),
    .b(\u2_Display/n3050 [8]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3074 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2292 (
    .a(\u2_Display/n3038 ),
    .b(\u2_Display/n3050 [9]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3073 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2293 (
    .a(\u2_Display/n3037 ),
    .b(\u2_Display/n3050 [10]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3072 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2294 (
    .a(\u2_Display/n3036 ),
    .b(\u2_Display/n3050 [11]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3071 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2295 (
    .a(\u2_Display/n3035 ),
    .b(\u2_Display/n3050 [12]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3070 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2296 (
    .a(\u2_Display/n3034 ),
    .b(\u2_Display/n3050 [13]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3069 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2297 (
    .a(\u2_Display/n3033 ),
    .b(\u2_Display/n3050 [14]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3068 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2298 (
    .a(\u2_Display/n3032 ),
    .b(\u2_Display/n3050 [15]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3067 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2299 (
    .a(\u2_Display/n3031 ),
    .b(\u2_Display/n3050 [16]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3066 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2300 (
    .a(\u2_Display/n3030 ),
    .b(\u2_Display/n3050 [17]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3065 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2301 (
    .a(\u2_Display/n3029 ),
    .b(\u2_Display/n3050 [18]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3064 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2302 (
    .a(\u2_Display/n3028 ),
    .b(\u2_Display/n3050 [19]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3063 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2303 (
    .a(\u2_Display/n3027 ),
    .b(\u2_Display/n3050 [20]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3062 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2304 (
    .a(\u2_Display/n3026 ),
    .b(\u2_Display/n3050 [21]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3061 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2305 (
    .a(\u2_Display/n3025 ),
    .b(\u2_Display/n3050 [22]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3060 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2306 (
    .a(\u2_Display/n3024 ),
    .b(\u2_Display/n3050 [23]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3059 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2307 (
    .a(\u2_Display/n3023 ),
    .b(\u2_Display/n3050 [24]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3058 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2308 (
    .a(\u2_Display/n3022 ),
    .b(\u2_Display/n3050 [25]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3057 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2309 (
    .a(\u2_Display/n3021 ),
    .b(\u2_Display/n3050 [26]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3056 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2310 (
    .a(\u2_Display/n3020 ),
    .b(\u2_Display/n3050 [27]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3055 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2311 (
    .a(\u2_Display/n3019 ),
    .b(\u2_Display/n3050 [28]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3054 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2312 (
    .a(\u2_Display/n3018 ),
    .b(\u2_Display/n3050 [29]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3053 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2313 (
    .a(\u2_Display/n3017 ),
    .b(\u2_Display/n3050 [30]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3052 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2314 (
    .a(\u2_Display/n3016 ),
    .b(\u2_Display/n3050 [31]),
    .c(\u2_Display/n3048 ),
    .o(\u2_Display/n3051 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2315 (
    .a(\u2_Display/n4205 ),
    .b(\u2_Display/n4208 [0]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4240 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2316 (
    .a(\u2_Display/n4204 ),
    .b(\u2_Display/n4208 [1]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4239 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2317 (
    .a(\u2_Display/n4203 ),
    .b(\u2_Display/n4208 [2]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4238 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2318 (
    .a(\u2_Display/n4202 ),
    .b(\u2_Display/n4208 [3]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4237 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2319 (
    .a(\u2_Display/n4201 ),
    .b(\u2_Display/n4208 [4]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4236 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2320 (
    .a(\u2_Display/n4200 ),
    .b(\u2_Display/n4208 [5]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4235 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2321 (
    .a(\u2_Display/n4199 ),
    .b(\u2_Display/n4208 [6]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4234 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2322 (
    .a(\u2_Display/n4198 ),
    .b(\u2_Display/n4208 [7]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4233 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2323 (
    .a(\u2_Display/n4197 ),
    .b(\u2_Display/n4208 [8]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4232 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2324 (
    .a(\u2_Display/n4196 ),
    .b(\u2_Display/n4208 [9]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4231 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2325 (
    .a(\u2_Display/n4195 ),
    .b(\u2_Display/n4208 [10]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4230 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2326 (
    .a(\u2_Display/n4194 ),
    .b(\u2_Display/n4208 [11]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4229 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2327 (
    .a(\u2_Display/n4193 ),
    .b(\u2_Display/n4208 [12]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4228 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2328 (
    .a(\u2_Display/n4192 ),
    .b(\u2_Display/n4208 [13]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4227 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2329 (
    .a(\u2_Display/n4191 ),
    .b(\u2_Display/n4208 [14]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4226 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2330 (
    .a(\u2_Display/n4190 ),
    .b(\u2_Display/n4208 [15]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4225 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2331 (
    .a(\u2_Display/n4189 ),
    .b(\u2_Display/n4208 [16]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4224 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2332 (
    .a(\u2_Display/n4188 ),
    .b(\u2_Display/n4208 [17]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4223 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2333 (
    .a(\u2_Display/n4187 ),
    .b(\u2_Display/n4208 [18]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4222 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2334 (
    .a(\u2_Display/n4186 ),
    .b(\u2_Display/n4208 [19]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4221 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2335 (
    .a(\u2_Display/n4185 ),
    .b(\u2_Display/n4208 [20]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4220 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2336 (
    .a(\u2_Display/n4184 ),
    .b(\u2_Display/n4208 [21]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4219 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2337 (
    .a(\u2_Display/n4183 ),
    .b(\u2_Display/n4208 [22]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4218 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2338 (
    .a(\u2_Display/n4182 ),
    .b(\u2_Display/n4208 [23]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4217 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2339 (
    .a(\u2_Display/n4181 ),
    .b(\u2_Display/n4208 [24]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4216 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2340 (
    .a(\u2_Display/n4180 ),
    .b(\u2_Display/n4208 [25]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4215 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2341 (
    .a(\u2_Display/n4179 ),
    .b(\u2_Display/n4208 [26]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4214 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2342 (
    .a(\u2_Display/n4178 ),
    .b(\u2_Display/n4208 [27]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4213 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2343 (
    .a(\u2_Display/n4177 ),
    .b(\u2_Display/n4208 [28]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4212 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2344 (
    .a(\u2_Display/n4176 ),
    .b(\u2_Display/n4208 [29]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4211 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2345 (
    .a(\u2_Display/n4175 ),
    .b(\u2_Display/n4208 [30]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4210 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2346 (
    .a(\u2_Display/n4174 ),
    .b(\u2_Display/n4208 [31]),
    .c(\u2_Display/n4206 ),
    .o(\u2_Display/n4209 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2347 (
    .a(\u2_Display/n5328 ),
    .b(\u2_Display/n5331 [0]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5363 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2348 (
    .a(\u2_Display/n5327 ),
    .b(\u2_Display/n5331 [1]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5362 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2349 (
    .a(\u2_Display/n5326 ),
    .b(\u2_Display/n5331 [2]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5361 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2350 (
    .a(\u2_Display/n5325 ),
    .b(\u2_Display/n5331 [3]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5360 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2351 (
    .a(\u2_Display/n5324 ),
    .b(\u2_Display/n5331 [4]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5359 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2352 (
    .a(\u2_Display/n5323 ),
    .b(\u2_Display/n5331 [5]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5358 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2353 (
    .a(\u2_Display/n5322 ),
    .b(\u2_Display/n5331 [6]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5357 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2354 (
    .a(\u2_Display/n5321 ),
    .b(\u2_Display/n5331 [7]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5356 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2355 (
    .a(\u2_Display/n5320 ),
    .b(\u2_Display/n5331 [8]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5355 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2356 (
    .a(\u2_Display/n5319 ),
    .b(\u2_Display/n5331 [9]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5354 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2357 (
    .a(\u2_Display/n5318 ),
    .b(\u2_Display/n5331 [10]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5353 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2358 (
    .a(\u2_Display/n5317 ),
    .b(\u2_Display/n5331 [11]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5352 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2359 (
    .a(\u2_Display/n5316 ),
    .b(\u2_Display/n5331 [12]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5351 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2360 (
    .a(\u2_Display/n5315 ),
    .b(\u2_Display/n5331 [13]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5350 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2361 (
    .a(\u2_Display/n5314 ),
    .b(\u2_Display/n5331 [14]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5349 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2362 (
    .a(\u2_Display/n5313 ),
    .b(\u2_Display/n5331 [15]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5348 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2363 (
    .a(\u2_Display/n5312 ),
    .b(\u2_Display/n5331 [16]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5347 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2364 (
    .a(\u2_Display/n5311 ),
    .b(\u2_Display/n5331 [17]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5346 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2365 (
    .a(\u2_Display/n5310 ),
    .b(\u2_Display/n5331 [18]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5345 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2366 (
    .a(\u2_Display/n5309 ),
    .b(\u2_Display/n5331 [19]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5344 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2367 (
    .a(\u2_Display/n5308 ),
    .b(\u2_Display/n5331 [20]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5343 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2368 (
    .a(\u2_Display/n5307 ),
    .b(\u2_Display/n5331 [21]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5342 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2369 (
    .a(\u2_Display/n5306 ),
    .b(\u2_Display/n5331 [22]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5341 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2370 (
    .a(\u2_Display/n5305 ),
    .b(\u2_Display/n5331 [23]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5340 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2371 (
    .a(\u2_Display/n5304 ),
    .b(\u2_Display/n5331 [24]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5339 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2372 (
    .a(\u2_Display/n5303 ),
    .b(\u2_Display/n5331 [25]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5338 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2373 (
    .a(\u2_Display/n5302 ),
    .b(\u2_Display/n5331 [26]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5337 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2374 (
    .a(\u2_Display/n5301 ),
    .b(\u2_Display/n5331 [27]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5336 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2375 (
    .a(\u2_Display/n5300 ),
    .b(\u2_Display/n5331 [28]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5335 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2376 (
    .a(\u2_Display/n5299 ),
    .b(\u2_Display/n5331 [29]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5334 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2377 (
    .a(\u2_Display/n5298 ),
    .b(\u2_Display/n5331 [30]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5333 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2378 (
    .a(\u2_Display/n5297 ),
    .b(\u2_Display/n5331 [31]),
    .c(\u2_Display/n5329 ),
    .o(\u2_Display/n5332 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2379 (
    .a(\u2_Display/n836 ),
    .b(\u2_Display/n839 [0]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n871 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2380 (
    .a(\u2_Display/n835 ),
    .b(\u2_Display/n839 [1]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n870 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2381 (
    .a(\u2_Display/n834 ),
    .b(\u2_Display/n839 [2]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n869 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2382 (
    .a(\u2_Display/n833 ),
    .b(\u2_Display/n839 [3]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n868 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2383 (
    .a(\u2_Display/n832 ),
    .b(\u2_Display/n839 [4]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n867 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2384 (
    .a(\u2_Display/n831 ),
    .b(\u2_Display/n839 [5]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n866 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2385 (
    .a(\u2_Display/n830 ),
    .b(\u2_Display/n839 [6]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n865 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2386 (
    .a(\u2_Display/n829 ),
    .b(\u2_Display/n839 [7]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n864 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2387 (
    .a(\u2_Display/n828 ),
    .b(\u2_Display/n839 [8]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n863 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2388 (
    .a(\u2_Display/n827 ),
    .b(\u2_Display/n839 [9]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n862 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2389 (
    .a(\u2_Display/n826 ),
    .b(\u2_Display/n839 [10]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n861 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2390 (
    .a(\u2_Display/n825 ),
    .b(\u2_Display/n839 [11]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n860 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2391 (
    .a(\u2_Display/n824 ),
    .b(\u2_Display/n839 [12]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n859 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2392 (
    .a(\u2_Display/n823 ),
    .b(\u2_Display/n839 [13]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n858 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2393 (
    .a(\u2_Display/n822 ),
    .b(\u2_Display/n839 [14]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n857 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2394 (
    .a(\u2_Display/n821 ),
    .b(\u2_Display/n839 [15]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n856 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2395 (
    .a(\u2_Display/n820 ),
    .b(\u2_Display/n839 [16]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n855 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2396 (
    .a(\u2_Display/n819 ),
    .b(\u2_Display/n839 [17]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n854 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2397 (
    .a(\u2_Display/n818 ),
    .b(\u2_Display/n839 [18]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n853 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2398 (
    .a(\u2_Display/n817 ),
    .b(\u2_Display/n839 [19]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n852 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2399 (
    .a(\u2_Display/n816 ),
    .b(\u2_Display/n839 [20]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n851 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2400 (
    .a(\u2_Display/n815 ),
    .b(\u2_Display/n839 [21]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n850 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2401 (
    .a(\u2_Display/n814 ),
    .b(\u2_Display/n839 [22]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n849 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2402 (
    .a(\u2_Display/n813 ),
    .b(\u2_Display/n839 [23]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n848 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2403 (
    .a(\u2_Display/n812 ),
    .b(\u2_Display/n839 [24]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n847 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2404 (
    .a(\u2_Display/n811 ),
    .b(\u2_Display/n839 [25]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n846 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2405 (
    .a(\u2_Display/n810 ),
    .b(\u2_Display/n839 [26]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n845 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2406 (
    .a(\u2_Display/n809 ),
    .b(\u2_Display/n839 [27]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n844 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2407 (
    .a(\u2_Display/n808 ),
    .b(\u2_Display/n839 [28]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n843 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2408 (
    .a(\u2_Display/n807 ),
    .b(\u2_Display/n839 [29]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n842 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2409 (
    .a(\u2_Display/n806 ),
    .b(\u2_Display/n839 [30]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n841 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2410 (
    .a(\u2_Display/n805 ),
    .b(\u2_Display/n839 [31]),
    .c(\u2_Display/n837 ),
    .o(\u2_Display/n840 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2411 (
    .a(\u2_Display/n1959 ),
    .b(\u2_Display/n1962 [0]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1994 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2412 (
    .a(\u2_Display/n1958 ),
    .b(\u2_Display/n1962 [1]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1993 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2413 (
    .a(\u2_Display/n1957 ),
    .b(\u2_Display/n1962 [2]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1992 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2414 (
    .a(\u2_Display/n1956 ),
    .b(\u2_Display/n1962 [3]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1991 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2415 (
    .a(\u2_Display/n1955 ),
    .b(\u2_Display/n1962 [4]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1990 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2416 (
    .a(\u2_Display/n1954 ),
    .b(\u2_Display/n1962 [5]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1989 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2417 (
    .a(\u2_Display/n1953 ),
    .b(\u2_Display/n1962 [6]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1988 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2418 (
    .a(\u2_Display/n1952 ),
    .b(\u2_Display/n1962 [7]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1987 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2419 (
    .a(\u2_Display/n1951 ),
    .b(\u2_Display/n1962 [8]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1986 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2420 (
    .a(\u2_Display/n1950 ),
    .b(\u2_Display/n1962 [9]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1985 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2421 (
    .a(\u2_Display/n1949 ),
    .b(\u2_Display/n1962 [10]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1984 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2422 (
    .a(\u2_Display/n1948 ),
    .b(\u2_Display/n1962 [11]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1983 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2423 (
    .a(\u2_Display/n1947 ),
    .b(\u2_Display/n1962 [12]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1982 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2424 (
    .a(\u2_Display/n1946 ),
    .b(\u2_Display/n1962 [13]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1981 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2425 (
    .a(\u2_Display/n1945 ),
    .b(\u2_Display/n1962 [14]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1980 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2426 (
    .a(\u2_Display/n1944 ),
    .b(\u2_Display/n1962 [15]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1979 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2427 (
    .a(\u2_Display/n1943 ),
    .b(\u2_Display/n1962 [16]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1978 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2428 (
    .a(\u2_Display/n1942 ),
    .b(\u2_Display/n1962 [17]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1977 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2429 (
    .a(\u2_Display/n1941 ),
    .b(\u2_Display/n1962 [18]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1976 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2430 (
    .a(\u2_Display/n1940 ),
    .b(\u2_Display/n1962 [19]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1975 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2431 (
    .a(\u2_Display/n1939 ),
    .b(\u2_Display/n1962 [20]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1974 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2432 (
    .a(\u2_Display/n1938 ),
    .b(\u2_Display/n1962 [21]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1973 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2433 (
    .a(\u2_Display/n1937 ),
    .b(\u2_Display/n1962 [22]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1972 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2434 (
    .a(\u2_Display/n1936 ),
    .b(\u2_Display/n1962 [23]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1971 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2435 (
    .a(\u2_Display/n1935 ),
    .b(\u2_Display/n1962 [24]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1970 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2436 (
    .a(\u2_Display/n1934 ),
    .b(\u2_Display/n1962 [25]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1969 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2437 (
    .a(\u2_Display/n1933 ),
    .b(\u2_Display/n1962 [26]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1968 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2438 (
    .a(\u2_Display/n1932 ),
    .b(\u2_Display/n1962 [27]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1967 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2439 (
    .a(\u2_Display/n1931 ),
    .b(\u2_Display/n1962 [28]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1966 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2440 (
    .a(\u2_Display/n1930 ),
    .b(\u2_Display/n1962 [29]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1965 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2441 (
    .a(\u2_Display/n1929 ),
    .b(\u2_Display/n1962 [30]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1964 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2442 (
    .a(\u2_Display/n1928 ),
    .b(\u2_Display/n1962 [31]),
    .c(\u2_Display/n1960 ),
    .o(\u2_Display/n1963 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2443 (
    .a(\u2_Display/n3082 ),
    .b(\u2_Display/n3085 [0]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3117 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2444 (
    .a(\u2_Display/n3081 ),
    .b(\u2_Display/n3085 [1]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3116 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2445 (
    .a(\u2_Display/n3080 ),
    .b(\u2_Display/n3085 [2]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3115 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2446 (
    .a(\u2_Display/n3079 ),
    .b(\u2_Display/n3085 [3]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3114 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2447 (
    .a(\u2_Display/n3078 ),
    .b(\u2_Display/n3085 [4]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3113 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2448 (
    .a(\u2_Display/n3077 ),
    .b(\u2_Display/n3085 [5]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3112 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2449 (
    .a(\u2_Display/n3076 ),
    .b(\u2_Display/n3085 [6]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3111 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2450 (
    .a(\u2_Display/n3075 ),
    .b(\u2_Display/n3085 [7]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3110 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2451 (
    .a(\u2_Display/n3074 ),
    .b(\u2_Display/n3085 [8]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3109 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2452 (
    .a(\u2_Display/n3073 ),
    .b(\u2_Display/n3085 [9]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3108 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2453 (
    .a(\u2_Display/n3072 ),
    .b(\u2_Display/n3085 [10]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3107 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2454 (
    .a(\u2_Display/n3071 ),
    .b(\u2_Display/n3085 [11]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3106 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2455 (
    .a(\u2_Display/n3070 ),
    .b(\u2_Display/n3085 [12]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3105 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2456 (
    .a(\u2_Display/n3069 ),
    .b(\u2_Display/n3085 [13]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3104 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2457 (
    .a(\u2_Display/n3068 ),
    .b(\u2_Display/n3085 [14]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3103 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2458 (
    .a(\u2_Display/n3067 ),
    .b(\u2_Display/n3085 [15]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3102 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2459 (
    .a(\u2_Display/n3066 ),
    .b(\u2_Display/n3085 [16]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3101 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2460 (
    .a(\u2_Display/n3065 ),
    .b(\u2_Display/n3085 [17]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3100 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2461 (
    .a(\u2_Display/n3064 ),
    .b(\u2_Display/n3085 [18]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3099 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2462 (
    .a(\u2_Display/n3063 ),
    .b(\u2_Display/n3085 [19]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3098 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2463 (
    .a(\u2_Display/n3062 ),
    .b(\u2_Display/n3085 [20]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3097 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2464 (
    .a(\u2_Display/n3061 ),
    .b(\u2_Display/n3085 [21]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3096 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2465 (
    .a(\u2_Display/n3060 ),
    .b(\u2_Display/n3085 [22]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3095 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2466 (
    .a(\u2_Display/n3059 ),
    .b(\u2_Display/n3085 [23]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3094 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2467 (
    .a(\u2_Display/n3058 ),
    .b(\u2_Display/n3085 [24]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3093 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2468 (
    .a(\u2_Display/n3057 ),
    .b(\u2_Display/n3085 [25]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3092 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2469 (
    .a(\u2_Display/n3056 ),
    .b(\u2_Display/n3085 [26]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3091 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2470 (
    .a(\u2_Display/n3055 ),
    .b(\u2_Display/n3085 [27]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3090 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2471 (
    .a(\u2_Display/n3054 ),
    .b(\u2_Display/n3085 [28]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3089 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2472 (
    .a(\u2_Display/n3053 ),
    .b(\u2_Display/n3085 [29]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3088 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2473 (
    .a(\u2_Display/n3052 ),
    .b(\u2_Display/n3085 [30]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3087 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2474 (
    .a(\u2_Display/n3051 ),
    .b(\u2_Display/n3085 [31]),
    .c(\u2_Display/n3083 ),
    .o(\u2_Display/n3086 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2475 (
    .a(\u2_Display/n4240 ),
    .b(\u2_Display/n4243 [0]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4275 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2476 (
    .a(\u2_Display/n4239 ),
    .b(\u2_Display/n4243 [1]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4274 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2477 (
    .a(\u2_Display/n4238 ),
    .b(\u2_Display/n4243 [2]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4273 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2478 (
    .a(\u2_Display/n4237 ),
    .b(\u2_Display/n4243 [3]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4272 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2479 (
    .a(\u2_Display/n4236 ),
    .b(\u2_Display/n4243 [4]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4271 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2480 (
    .a(\u2_Display/n4235 ),
    .b(\u2_Display/n4243 [5]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4270 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2481 (
    .a(\u2_Display/n4234 ),
    .b(\u2_Display/n4243 [6]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4269 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2482 (
    .a(\u2_Display/n4233 ),
    .b(\u2_Display/n4243 [7]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4268 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2483 (
    .a(\u2_Display/n4232 ),
    .b(\u2_Display/n4243 [8]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4267 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2484 (
    .a(\u2_Display/n4231 ),
    .b(\u2_Display/n4243 [9]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4266 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2485 (
    .a(\u2_Display/n4230 ),
    .b(\u2_Display/n4243 [10]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4265 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2486 (
    .a(\u2_Display/n4229 ),
    .b(\u2_Display/n4243 [11]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4264 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2487 (
    .a(\u2_Display/n4228 ),
    .b(\u2_Display/n4243 [12]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4263 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2488 (
    .a(\u2_Display/n4227 ),
    .b(\u2_Display/n4243 [13]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4262 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2489 (
    .a(\u2_Display/n4226 ),
    .b(\u2_Display/n4243 [14]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4261 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2490 (
    .a(\u2_Display/n4225 ),
    .b(\u2_Display/n4243 [15]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4260 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2491 (
    .a(\u2_Display/n4224 ),
    .b(\u2_Display/n4243 [16]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4259 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2492 (
    .a(\u2_Display/n4223 ),
    .b(\u2_Display/n4243 [17]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4258 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2493 (
    .a(\u2_Display/n4222 ),
    .b(\u2_Display/n4243 [18]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4257 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2494 (
    .a(\u2_Display/n4221 ),
    .b(\u2_Display/n4243 [19]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4256 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2495 (
    .a(\u2_Display/n4220 ),
    .b(\u2_Display/n4243 [20]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4255 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2496 (
    .a(\u2_Display/n4219 ),
    .b(\u2_Display/n4243 [21]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4254 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2497 (
    .a(\u2_Display/n4218 ),
    .b(\u2_Display/n4243 [22]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4253 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2498 (
    .a(\u2_Display/n4217 ),
    .b(\u2_Display/n4243 [23]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4252 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2499 (
    .a(\u2_Display/n4216 ),
    .b(\u2_Display/n4243 [24]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4251 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2500 (
    .a(\u2_Display/n4215 ),
    .b(\u2_Display/n4243 [25]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4250 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2501 (
    .a(\u2_Display/n4214 ),
    .b(\u2_Display/n4243 [26]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4249 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2502 (
    .a(\u2_Display/n4213 ),
    .b(\u2_Display/n4243 [27]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4248 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2503 (
    .a(\u2_Display/n4212 ),
    .b(\u2_Display/n4243 [28]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4247 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2504 (
    .a(\u2_Display/n4211 ),
    .b(\u2_Display/n4243 [29]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4246 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2505 (
    .a(\u2_Display/n4210 ),
    .b(\u2_Display/n4243 [30]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4245 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2506 (
    .a(\u2_Display/n4209 ),
    .b(\u2_Display/n4243 [31]),
    .c(\u2_Display/n4241 ),
    .o(\u2_Display/n4244 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2507 (
    .a(\u2_Display/n5363 ),
    .b(\u2_Display/n5366 [0]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5398 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2508 (
    .a(\u2_Display/n5362 ),
    .b(\u2_Display/n5366 [1]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5397 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2509 (
    .a(\u2_Display/n5361 ),
    .b(\u2_Display/n5366 [2]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5396 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2510 (
    .a(\u2_Display/n5360 ),
    .b(\u2_Display/n5366 [3]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5395 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2511 (
    .a(\u2_Display/n5359 ),
    .b(\u2_Display/n5366 [4]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5394 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2512 (
    .a(\u2_Display/n5358 ),
    .b(\u2_Display/n5366 [5]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5393 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2513 (
    .a(\u2_Display/n5357 ),
    .b(\u2_Display/n5366 [6]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5392 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2514 (
    .a(\u2_Display/n5356 ),
    .b(\u2_Display/n5366 [7]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5391 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2515 (
    .a(\u2_Display/n5355 ),
    .b(\u2_Display/n5366 [8]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5390 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2516 (
    .a(\u2_Display/n5354 ),
    .b(\u2_Display/n5366 [9]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5389 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2517 (
    .a(\u2_Display/n5353 ),
    .b(\u2_Display/n5366 [10]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5388 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2518 (
    .a(\u2_Display/n5352 ),
    .b(\u2_Display/n5366 [11]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5387 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2519 (
    .a(\u2_Display/n5351 ),
    .b(\u2_Display/n5366 [12]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5386 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2520 (
    .a(\u2_Display/n5350 ),
    .b(\u2_Display/n5366 [13]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5385 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2521 (
    .a(\u2_Display/n5349 ),
    .b(\u2_Display/n5366 [14]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5384 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2522 (
    .a(\u2_Display/n5348 ),
    .b(\u2_Display/n5366 [15]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5383 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2523 (
    .a(\u2_Display/n5347 ),
    .b(\u2_Display/n5366 [16]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5382 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2524 (
    .a(\u2_Display/n5346 ),
    .b(\u2_Display/n5366 [17]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5381 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2525 (
    .a(\u2_Display/n5345 ),
    .b(\u2_Display/n5366 [18]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5380 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2526 (
    .a(\u2_Display/n5344 ),
    .b(\u2_Display/n5366 [19]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5379 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2527 (
    .a(\u2_Display/n5343 ),
    .b(\u2_Display/n5366 [20]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5378 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2528 (
    .a(\u2_Display/n5342 ),
    .b(\u2_Display/n5366 [21]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5377 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2529 (
    .a(\u2_Display/n5341 ),
    .b(\u2_Display/n5366 [22]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5376 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2530 (
    .a(\u2_Display/n5340 ),
    .b(\u2_Display/n5366 [23]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5375 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2531 (
    .a(\u2_Display/n5339 ),
    .b(\u2_Display/n5366 [24]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5374 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2532 (
    .a(\u2_Display/n5338 ),
    .b(\u2_Display/n5366 [25]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5373 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2533 (
    .a(\u2_Display/n5337 ),
    .b(\u2_Display/n5366 [26]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5372 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2534 (
    .a(\u2_Display/n5336 ),
    .b(\u2_Display/n5366 [27]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5371 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2535 (
    .a(\u2_Display/n5335 ),
    .b(\u2_Display/n5366 [28]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5370 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2536 (
    .a(\u2_Display/n5334 ),
    .b(\u2_Display/n5366 [29]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5369 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2537 (
    .a(\u2_Display/n5333 ),
    .b(\u2_Display/n5366 [30]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5368 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2538 (
    .a(\u2_Display/n5332 ),
    .b(\u2_Display/n5366 [31]),
    .c(\u2_Display/n5364 ),
    .o(\u2_Display/n5367 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2539 (
    .a(\u2_Display/n871 ),
    .b(\u2_Display/n874 [0]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n906 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2540 (
    .a(\u2_Display/n870 ),
    .b(\u2_Display/n874 [1]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n905 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2541 (
    .a(\u2_Display/n869 ),
    .b(\u2_Display/n874 [2]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n904 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2542 (
    .a(\u2_Display/n868 ),
    .b(\u2_Display/n874 [3]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n903 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2543 (
    .a(\u2_Display/n867 ),
    .b(\u2_Display/n874 [4]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n902 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2544 (
    .a(\u2_Display/n866 ),
    .b(\u2_Display/n874 [5]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n901 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2545 (
    .a(\u2_Display/n865 ),
    .b(\u2_Display/n874 [6]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n900 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2546 (
    .a(\u2_Display/n864 ),
    .b(\u2_Display/n874 [7]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n899 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2547 (
    .a(\u2_Display/n863 ),
    .b(\u2_Display/n874 [8]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n898 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2548 (
    .a(\u2_Display/n862 ),
    .b(\u2_Display/n874 [9]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n897 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2549 (
    .a(\u2_Display/n861 ),
    .b(\u2_Display/n874 [10]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n896 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2550 (
    .a(\u2_Display/n860 ),
    .b(\u2_Display/n874 [11]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n895 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2551 (
    .a(\u2_Display/n859 ),
    .b(\u2_Display/n874 [12]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n894 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2552 (
    .a(\u2_Display/n858 ),
    .b(\u2_Display/n874 [13]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n893 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2553 (
    .a(\u2_Display/n857 ),
    .b(\u2_Display/n874 [14]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n892 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2554 (
    .a(\u2_Display/n856 ),
    .b(\u2_Display/n874 [15]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n891 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2555 (
    .a(\u2_Display/n855 ),
    .b(\u2_Display/n874 [16]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n890 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2556 (
    .a(\u2_Display/n854 ),
    .b(\u2_Display/n874 [17]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n889 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2557 (
    .a(\u2_Display/n853 ),
    .b(\u2_Display/n874 [18]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n888 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2558 (
    .a(\u2_Display/n852 ),
    .b(\u2_Display/n874 [19]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n887 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2559 (
    .a(\u2_Display/n851 ),
    .b(\u2_Display/n874 [20]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n886 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2560 (
    .a(\u2_Display/n850 ),
    .b(\u2_Display/n874 [21]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n885 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2561 (
    .a(\u2_Display/n849 ),
    .b(\u2_Display/n874 [22]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n884 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2562 (
    .a(\u2_Display/n848 ),
    .b(\u2_Display/n874 [23]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n883 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2563 (
    .a(\u2_Display/n847 ),
    .b(\u2_Display/n874 [24]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n882 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2564 (
    .a(\u2_Display/n846 ),
    .b(\u2_Display/n874 [25]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n881 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2565 (
    .a(\u2_Display/n845 ),
    .b(\u2_Display/n874 [26]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n880 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2566 (
    .a(\u2_Display/n844 ),
    .b(\u2_Display/n874 [27]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n879 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2567 (
    .a(\u2_Display/n843 ),
    .b(\u2_Display/n874 [28]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n878 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2568 (
    .a(\u2_Display/n842 ),
    .b(\u2_Display/n874 [29]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n877 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2569 (
    .a(\u2_Display/n841 ),
    .b(\u2_Display/n874 [30]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n876 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2570 (
    .a(\u2_Display/n840 ),
    .b(\u2_Display/n874 [31]),
    .c(\u2_Display/n872 ),
    .o(\u2_Display/n875 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2571 (
    .a(\u2_Display/n1994 ),
    .b(\u2_Display/n1997 [0]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2029 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2572 (
    .a(\u2_Display/n1993 ),
    .b(\u2_Display/n1997 [1]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2028 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2573 (
    .a(\u2_Display/n1992 ),
    .b(\u2_Display/n1997 [2]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2027 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2574 (
    .a(\u2_Display/n1991 ),
    .b(\u2_Display/n1997 [3]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2026 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2575 (
    .a(\u2_Display/n1990 ),
    .b(\u2_Display/n1997 [4]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2025 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2576 (
    .a(\u2_Display/n1989 ),
    .b(\u2_Display/n1997 [5]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2024 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2577 (
    .a(\u2_Display/n1988 ),
    .b(\u2_Display/n1997 [6]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2023 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2578 (
    .a(\u2_Display/n1987 ),
    .b(\u2_Display/n1997 [7]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2022 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2579 (
    .a(\u2_Display/n1986 ),
    .b(\u2_Display/n1997 [8]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2021 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2580 (
    .a(\u2_Display/n1985 ),
    .b(\u2_Display/n1997 [9]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2020 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2581 (
    .a(\u2_Display/n1984 ),
    .b(\u2_Display/n1997 [10]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2019 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2582 (
    .a(\u2_Display/n1983 ),
    .b(\u2_Display/n1997 [11]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2018 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2583 (
    .a(\u2_Display/n1982 ),
    .b(\u2_Display/n1997 [12]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2017 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2584 (
    .a(\u2_Display/n1981 ),
    .b(\u2_Display/n1997 [13]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2016 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2585 (
    .a(\u2_Display/n1980 ),
    .b(\u2_Display/n1997 [14]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2015 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2586 (
    .a(\u2_Display/n1979 ),
    .b(\u2_Display/n1997 [15]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2014 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2587 (
    .a(\u2_Display/n1978 ),
    .b(\u2_Display/n1997 [16]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2013 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2588 (
    .a(\u2_Display/n1977 ),
    .b(\u2_Display/n1997 [17]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2012 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2589 (
    .a(\u2_Display/n1976 ),
    .b(\u2_Display/n1997 [18]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2011 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2590 (
    .a(\u2_Display/n1975 ),
    .b(\u2_Display/n1997 [19]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2010 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2591 (
    .a(\u2_Display/n1974 ),
    .b(\u2_Display/n1997 [20]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2009 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2592 (
    .a(\u2_Display/n1973 ),
    .b(\u2_Display/n1997 [21]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2008 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2593 (
    .a(\u2_Display/n1972 ),
    .b(\u2_Display/n1997 [22]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2007 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2594 (
    .a(\u2_Display/n1971 ),
    .b(\u2_Display/n1997 [23]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2006 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2595 (
    .a(\u2_Display/n1970 ),
    .b(\u2_Display/n1997 [24]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2005 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2596 (
    .a(\u2_Display/n1969 ),
    .b(\u2_Display/n1997 [25]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2004 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2597 (
    .a(\u2_Display/n1968 ),
    .b(\u2_Display/n1997 [26]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2003 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2598 (
    .a(\u2_Display/n1967 ),
    .b(\u2_Display/n1997 [27]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2002 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2599 (
    .a(\u2_Display/n1966 ),
    .b(\u2_Display/n1997 [28]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2001 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2600 (
    .a(\u2_Display/n1965 ),
    .b(\u2_Display/n1997 [29]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n2000 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2601 (
    .a(\u2_Display/n1964 ),
    .b(\u2_Display/n1997 [30]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n1999 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2602 (
    .a(\u2_Display/n1963 ),
    .b(\u2_Display/n1997 [31]),
    .c(\u2_Display/n1995 ),
    .o(\u2_Display/n1998 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2603 (
    .a(\u2_Display/n3117 ),
    .b(\u2_Display/n3120 [0]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3152 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2604 (
    .a(\u2_Display/n3116 ),
    .b(\u2_Display/n3120 [1]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3151 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2605 (
    .a(\u2_Display/n3115 ),
    .b(\u2_Display/n3120 [2]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3150 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2606 (
    .a(\u2_Display/n3114 ),
    .b(\u2_Display/n3120 [3]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3149 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2607 (
    .a(\u2_Display/n3113 ),
    .b(\u2_Display/n3120 [4]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3148 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2608 (
    .a(\u2_Display/n3112 ),
    .b(\u2_Display/n3120 [5]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3147 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2609 (
    .a(\u2_Display/n3111 ),
    .b(\u2_Display/n3120 [6]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3146 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2610 (
    .a(\u2_Display/n3110 ),
    .b(\u2_Display/n3120 [7]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3145 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2611 (
    .a(\u2_Display/n3109 ),
    .b(\u2_Display/n3120 [8]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3144 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2612 (
    .a(\u2_Display/n3108 ),
    .b(\u2_Display/n3120 [9]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3143 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2613 (
    .a(\u2_Display/n3107 ),
    .b(\u2_Display/n3120 [10]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3142 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2614 (
    .a(\u2_Display/n3106 ),
    .b(\u2_Display/n3120 [11]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3141 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2615 (
    .a(\u2_Display/n3105 ),
    .b(\u2_Display/n3120 [12]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3140 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2616 (
    .a(\u2_Display/n3104 ),
    .b(\u2_Display/n3120 [13]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3139 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2617 (
    .a(\u2_Display/n3103 ),
    .b(\u2_Display/n3120 [14]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3138 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2618 (
    .a(\u2_Display/n3102 ),
    .b(\u2_Display/n3120 [15]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3137 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2619 (
    .a(\u2_Display/n3101 ),
    .b(\u2_Display/n3120 [16]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3136 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2620 (
    .a(\u2_Display/n3100 ),
    .b(\u2_Display/n3120 [17]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3135 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2621 (
    .a(\u2_Display/n3099 ),
    .b(\u2_Display/n3120 [18]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3134 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2622 (
    .a(\u2_Display/n3098 ),
    .b(\u2_Display/n3120 [19]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3133 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2623 (
    .a(\u2_Display/n3097 ),
    .b(\u2_Display/n3120 [20]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3132 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2624 (
    .a(\u2_Display/n3096 ),
    .b(\u2_Display/n3120 [21]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3131 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2625 (
    .a(\u2_Display/n3095 ),
    .b(\u2_Display/n3120 [22]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3130 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2626 (
    .a(\u2_Display/n3094 ),
    .b(\u2_Display/n3120 [23]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3129 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2627 (
    .a(\u2_Display/n3093 ),
    .b(\u2_Display/n3120 [24]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3128 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2628 (
    .a(\u2_Display/n3092 ),
    .b(\u2_Display/n3120 [25]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3127 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2629 (
    .a(\u2_Display/n3091 ),
    .b(\u2_Display/n3120 [26]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3126 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2630 (
    .a(\u2_Display/n3090 ),
    .b(\u2_Display/n3120 [27]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3125 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2631 (
    .a(\u2_Display/n3089 ),
    .b(\u2_Display/n3120 [28]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3124 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2632 (
    .a(\u2_Display/n3088 ),
    .b(\u2_Display/n3120 [29]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3123 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2633 (
    .a(\u2_Display/n3087 ),
    .b(\u2_Display/n3120 [30]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3122 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2634 (
    .a(\u2_Display/n3086 ),
    .b(\u2_Display/n3120 [31]),
    .c(\u2_Display/n3118 ),
    .o(\u2_Display/n3121 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2635 (
    .a(\u2_Display/n4275 ),
    .b(\u2_Display/n4278 [0]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4310 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2636 (
    .a(\u2_Display/n4274 ),
    .b(\u2_Display/n4278 [1]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4309 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2637 (
    .a(\u2_Display/n4273 ),
    .b(\u2_Display/n4278 [2]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4308 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2638 (
    .a(\u2_Display/n4272 ),
    .b(\u2_Display/n4278 [3]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4307 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2639 (
    .a(\u2_Display/n4271 ),
    .b(\u2_Display/n4278 [4]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4306 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2640 (
    .a(\u2_Display/n4270 ),
    .b(\u2_Display/n4278 [5]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4305 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2641 (
    .a(\u2_Display/n4269 ),
    .b(\u2_Display/n4278 [6]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4304 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2642 (
    .a(\u2_Display/n4268 ),
    .b(\u2_Display/n4278 [7]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4303 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2643 (
    .a(\u2_Display/n4267 ),
    .b(\u2_Display/n4278 [8]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4302 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2644 (
    .a(\u2_Display/n4266 ),
    .b(\u2_Display/n4278 [9]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4301 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2645 (
    .a(\u2_Display/n4265 ),
    .b(\u2_Display/n4278 [10]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4300 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2646 (
    .a(\u2_Display/n4264 ),
    .b(\u2_Display/n4278 [11]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4299 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2647 (
    .a(\u2_Display/n4263 ),
    .b(\u2_Display/n4278 [12]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4298 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2648 (
    .a(\u2_Display/n4262 ),
    .b(\u2_Display/n4278 [13]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4297 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2649 (
    .a(\u2_Display/n4261 ),
    .b(\u2_Display/n4278 [14]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4296 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2650 (
    .a(\u2_Display/n4260 ),
    .b(\u2_Display/n4278 [15]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4295 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2651 (
    .a(\u2_Display/n4259 ),
    .b(\u2_Display/n4278 [16]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4294 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2652 (
    .a(\u2_Display/n4258 ),
    .b(\u2_Display/n4278 [17]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4293 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2653 (
    .a(\u2_Display/n4257 ),
    .b(\u2_Display/n4278 [18]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4292 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2654 (
    .a(\u2_Display/n4256 ),
    .b(\u2_Display/n4278 [19]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4291 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2655 (
    .a(\u2_Display/n4255 ),
    .b(\u2_Display/n4278 [20]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4290 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2656 (
    .a(\u2_Display/n4254 ),
    .b(\u2_Display/n4278 [21]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4289 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2657 (
    .a(\u2_Display/n4253 ),
    .b(\u2_Display/n4278 [22]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4288 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2658 (
    .a(\u2_Display/n4252 ),
    .b(\u2_Display/n4278 [23]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4287 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2659 (
    .a(\u2_Display/n4251 ),
    .b(\u2_Display/n4278 [24]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4286 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2660 (
    .a(\u2_Display/n4250 ),
    .b(\u2_Display/n4278 [25]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4285 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2661 (
    .a(\u2_Display/n4249 ),
    .b(\u2_Display/n4278 [26]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4284 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2662 (
    .a(\u2_Display/n4248 ),
    .b(\u2_Display/n4278 [27]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4283 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2663 (
    .a(\u2_Display/n4247 ),
    .b(\u2_Display/n4278 [28]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4282 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2664 (
    .a(\u2_Display/n4246 ),
    .b(\u2_Display/n4278 [29]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4281 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2665 (
    .a(\u2_Display/n4245 ),
    .b(\u2_Display/n4278 [30]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4280 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2666 (
    .a(\u2_Display/n4244 ),
    .b(\u2_Display/n4278 [31]),
    .c(\u2_Display/n4276 ),
    .o(\u2_Display/n4279 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2667 (
    .a(\u2_Display/n5398 ),
    .b(\u2_Display/n5401 [0]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5433 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2668 (
    .a(\u2_Display/n5397 ),
    .b(\u2_Display/n5401 [1]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5432 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2669 (
    .a(\u2_Display/n5396 ),
    .b(\u2_Display/n5401 [2]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5431 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2670 (
    .a(\u2_Display/n5395 ),
    .b(\u2_Display/n5401 [3]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5430 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2671 (
    .a(\u2_Display/n5394 ),
    .b(\u2_Display/n5401 [4]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5429 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2672 (
    .a(\u2_Display/n5393 ),
    .b(\u2_Display/n5401 [5]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5428 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2673 (
    .a(\u2_Display/n5392 ),
    .b(\u2_Display/n5401 [6]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5427 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2674 (
    .a(\u2_Display/n5391 ),
    .b(\u2_Display/n5401 [7]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5426 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2675 (
    .a(\u2_Display/n5390 ),
    .b(\u2_Display/n5401 [8]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5425 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2676 (
    .a(\u2_Display/n5389 ),
    .b(\u2_Display/n5401 [9]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5424 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2677 (
    .a(\u2_Display/n5388 ),
    .b(\u2_Display/n5401 [10]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5423 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2678 (
    .a(\u2_Display/n5387 ),
    .b(\u2_Display/n5401 [11]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5422 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2679 (
    .a(\u2_Display/n5386 ),
    .b(\u2_Display/n5401 [12]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5421 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2680 (
    .a(\u2_Display/n5385 ),
    .b(\u2_Display/n5401 [13]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5420 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2681 (
    .a(\u2_Display/n5384 ),
    .b(\u2_Display/n5401 [14]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5419 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2682 (
    .a(\u2_Display/n5383 ),
    .b(\u2_Display/n5401 [15]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5418 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2683 (
    .a(\u2_Display/n5382 ),
    .b(\u2_Display/n5401 [16]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5417 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2684 (
    .a(\u2_Display/n5381 ),
    .b(\u2_Display/n5401 [17]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5416 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2685 (
    .a(\u2_Display/n5380 ),
    .b(\u2_Display/n5401 [18]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5415 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2686 (
    .a(\u2_Display/n5379 ),
    .b(\u2_Display/n5401 [19]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5414 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2687 (
    .a(\u2_Display/n5378 ),
    .b(\u2_Display/n5401 [20]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5413 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2688 (
    .a(\u2_Display/n5377 ),
    .b(\u2_Display/n5401 [21]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5412 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2689 (
    .a(\u2_Display/n5376 ),
    .b(\u2_Display/n5401 [22]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5411 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2690 (
    .a(\u2_Display/n5375 ),
    .b(\u2_Display/n5401 [23]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5410 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2691 (
    .a(\u2_Display/n5374 ),
    .b(\u2_Display/n5401 [24]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5409 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2692 (
    .a(\u2_Display/n5373 ),
    .b(\u2_Display/n5401 [25]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5408 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2693 (
    .a(\u2_Display/n5372 ),
    .b(\u2_Display/n5401 [26]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5407 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2694 (
    .a(\u2_Display/n5371 ),
    .b(\u2_Display/n5401 [27]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5406 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2695 (
    .a(\u2_Display/n5370 ),
    .b(\u2_Display/n5401 [28]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5405 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2696 (
    .a(\u2_Display/n5369 ),
    .b(\u2_Display/n5401 [29]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5404 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2697 (
    .a(\u2_Display/n5368 ),
    .b(\u2_Display/n5401 [30]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5403 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2698 (
    .a(\u2_Display/n5367 ),
    .b(\u2_Display/n5401 [31]),
    .c(\u2_Display/n5399 ),
    .o(\u2_Display/n5402 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2699 (
    .a(\u2_Display/n906 ),
    .b(\u2_Display/n909 [0]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n941 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2700 (
    .a(\u2_Display/n905 ),
    .b(\u2_Display/n909 [1]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n940 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2701 (
    .a(\u2_Display/n904 ),
    .b(\u2_Display/n909 [2]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n939 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2702 (
    .a(\u2_Display/n903 ),
    .b(\u2_Display/n909 [3]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n938 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2703 (
    .a(\u2_Display/n902 ),
    .b(\u2_Display/n909 [4]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n937 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2704 (
    .a(\u2_Display/n901 ),
    .b(\u2_Display/n909 [5]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n936 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2705 (
    .a(\u2_Display/n900 ),
    .b(\u2_Display/n909 [6]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n935 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2706 (
    .a(\u2_Display/n899 ),
    .b(\u2_Display/n909 [7]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n934 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2707 (
    .a(\u2_Display/n898 ),
    .b(\u2_Display/n909 [8]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n933 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2708 (
    .a(\u2_Display/n897 ),
    .b(\u2_Display/n909 [9]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n932 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2709 (
    .a(\u2_Display/n896 ),
    .b(\u2_Display/n909 [10]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n931 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2710 (
    .a(\u2_Display/n895 ),
    .b(\u2_Display/n909 [11]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n930 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2711 (
    .a(\u2_Display/n894 ),
    .b(\u2_Display/n909 [12]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n929 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2712 (
    .a(\u2_Display/n893 ),
    .b(\u2_Display/n909 [13]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n928 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2713 (
    .a(\u2_Display/n892 ),
    .b(\u2_Display/n909 [14]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n927 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2714 (
    .a(\u2_Display/n891 ),
    .b(\u2_Display/n909 [15]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n926 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2715 (
    .a(\u2_Display/n890 ),
    .b(\u2_Display/n909 [16]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n925 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2716 (
    .a(\u2_Display/n889 ),
    .b(\u2_Display/n909 [17]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n924 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2717 (
    .a(\u2_Display/n888 ),
    .b(\u2_Display/n909 [18]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n923 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2718 (
    .a(\u2_Display/n887 ),
    .b(\u2_Display/n909 [19]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n922 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2719 (
    .a(\u2_Display/n886 ),
    .b(\u2_Display/n909 [20]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n921 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2720 (
    .a(\u2_Display/n885 ),
    .b(\u2_Display/n909 [21]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n920 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2721 (
    .a(\u2_Display/n884 ),
    .b(\u2_Display/n909 [22]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n919 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2722 (
    .a(\u2_Display/n883 ),
    .b(\u2_Display/n909 [23]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n918 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2723 (
    .a(\u2_Display/n882 ),
    .b(\u2_Display/n909 [24]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n917 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2724 (
    .a(\u2_Display/n881 ),
    .b(\u2_Display/n909 [25]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n916 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2725 (
    .a(\u2_Display/n880 ),
    .b(\u2_Display/n909 [26]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n915 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2726 (
    .a(\u2_Display/n879 ),
    .b(\u2_Display/n909 [27]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n914 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2727 (
    .a(\u2_Display/n878 ),
    .b(\u2_Display/n909 [28]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n913 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2728 (
    .a(\u2_Display/n877 ),
    .b(\u2_Display/n909 [29]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n912 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2729 (
    .a(\u2_Display/n876 ),
    .b(\u2_Display/n909 [30]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n911 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2730 (
    .a(\u2_Display/n875 ),
    .b(\u2_Display/n909 [31]),
    .c(\u2_Display/n907 ),
    .o(\u2_Display/n910 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2731 (
    .a(\u2_Display/n2029 ),
    .b(\u2_Display/n2032 [0]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2064 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2732 (
    .a(\u2_Display/n2028 ),
    .b(\u2_Display/n2032 [1]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2063 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2733 (
    .a(\u2_Display/n2027 ),
    .b(\u2_Display/n2032 [2]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2062 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2734 (
    .a(\u2_Display/n2026 ),
    .b(\u2_Display/n2032 [3]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2061 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2735 (
    .a(\u2_Display/n2025 ),
    .b(\u2_Display/n2032 [4]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2060 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2736 (
    .a(\u2_Display/n2024 ),
    .b(\u2_Display/n2032 [5]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2059 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2737 (
    .a(\u2_Display/n2023 ),
    .b(\u2_Display/n2032 [6]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2058 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2738 (
    .a(\u2_Display/n2022 ),
    .b(\u2_Display/n2032 [7]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2057 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2739 (
    .a(\u2_Display/n2021 ),
    .b(\u2_Display/n2032 [8]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2056 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2740 (
    .a(\u2_Display/n2020 ),
    .b(\u2_Display/n2032 [9]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2055 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2741 (
    .a(\u2_Display/n2019 ),
    .b(\u2_Display/n2032 [10]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2054 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2742 (
    .a(\u2_Display/n2018 ),
    .b(\u2_Display/n2032 [11]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2053 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2743 (
    .a(\u2_Display/n2017 ),
    .b(\u2_Display/n2032 [12]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2052 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2744 (
    .a(\u2_Display/n2016 ),
    .b(\u2_Display/n2032 [13]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2051 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2745 (
    .a(\u2_Display/n2015 ),
    .b(\u2_Display/n2032 [14]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2050 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2746 (
    .a(\u2_Display/n2014 ),
    .b(\u2_Display/n2032 [15]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2049 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2747 (
    .a(\u2_Display/n2013 ),
    .b(\u2_Display/n2032 [16]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2048 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2748 (
    .a(\u2_Display/n2012 ),
    .b(\u2_Display/n2032 [17]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2047 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2749 (
    .a(\u2_Display/n2011 ),
    .b(\u2_Display/n2032 [18]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2046 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2750 (
    .a(\u2_Display/n2010 ),
    .b(\u2_Display/n2032 [19]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2045 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2751 (
    .a(\u2_Display/n2009 ),
    .b(\u2_Display/n2032 [20]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2044 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2752 (
    .a(\u2_Display/n2008 ),
    .b(\u2_Display/n2032 [21]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2043 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2753 (
    .a(\u2_Display/n2007 ),
    .b(\u2_Display/n2032 [22]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2042 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2754 (
    .a(\u2_Display/n2006 ),
    .b(\u2_Display/n2032 [23]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2041 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2755 (
    .a(\u2_Display/n2005 ),
    .b(\u2_Display/n2032 [24]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2040 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2756 (
    .a(\u2_Display/n2004 ),
    .b(\u2_Display/n2032 [25]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2039 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2757 (
    .a(\u2_Display/n2003 ),
    .b(\u2_Display/n2032 [26]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2038 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2758 (
    .a(\u2_Display/n2002 ),
    .b(\u2_Display/n2032 [27]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2037 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2759 (
    .a(\u2_Display/n2001 ),
    .b(\u2_Display/n2032 [28]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2036 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2760 (
    .a(\u2_Display/n2000 ),
    .b(\u2_Display/n2032 [29]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2035 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2761 (
    .a(\u2_Display/n1999 ),
    .b(\u2_Display/n2032 [30]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2034 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2762 (
    .a(\u2_Display/n1998 ),
    .b(\u2_Display/n2032 [31]),
    .c(\u2_Display/n2030 ),
    .o(\u2_Display/n2033 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2763 (
    .a(\u2_Display/n3152 ),
    .b(\u2_Display/n3155 [0]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3187 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2764 (
    .a(\u2_Display/n3151 ),
    .b(\u2_Display/n3155 [1]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3186 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2765 (
    .a(\u2_Display/n3150 ),
    .b(\u2_Display/n3155 [2]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3185 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2766 (
    .a(\u2_Display/n3149 ),
    .b(\u2_Display/n3155 [3]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3184 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2767 (
    .a(\u2_Display/n3148 ),
    .b(\u2_Display/n3155 [4]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3183 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2768 (
    .a(\u2_Display/n3147 ),
    .b(\u2_Display/n3155 [5]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3182 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2769 (
    .a(\u2_Display/n3146 ),
    .b(\u2_Display/n3155 [6]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3181 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2770 (
    .a(\u2_Display/n3145 ),
    .b(\u2_Display/n3155 [7]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3180 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2771 (
    .a(\u2_Display/n3144 ),
    .b(\u2_Display/n3155 [8]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3179 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2772 (
    .a(\u2_Display/n3143 ),
    .b(\u2_Display/n3155 [9]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3178 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2773 (
    .a(\u2_Display/n3142 ),
    .b(\u2_Display/n3155 [10]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3177 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2774 (
    .a(\u2_Display/n3141 ),
    .b(\u2_Display/n3155 [11]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3176 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2775 (
    .a(\u2_Display/n3140 ),
    .b(\u2_Display/n3155 [12]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3175 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2776 (
    .a(\u2_Display/n3139 ),
    .b(\u2_Display/n3155 [13]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3174 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2777 (
    .a(\u2_Display/n3138 ),
    .b(\u2_Display/n3155 [14]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3173 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2778 (
    .a(\u2_Display/n3137 ),
    .b(\u2_Display/n3155 [15]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3172 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2779 (
    .a(\u2_Display/n3136 ),
    .b(\u2_Display/n3155 [16]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3171 ));
  EG_PHY_PAD #(
    //.LOCATION("K14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u278 (
    .ipad(clk_24m),
    .di(clk_24m_pad));  // source/rtl/VGA_Demo.v(4)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2780 (
    .a(\u2_Display/n3135 ),
    .b(\u2_Display/n3155 [17]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3170 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2781 (
    .a(\u2_Display/n3134 ),
    .b(\u2_Display/n3155 [18]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3169 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2782 (
    .a(\u2_Display/n3133 ),
    .b(\u2_Display/n3155 [19]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3168 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2783 (
    .a(\u2_Display/n3132 ),
    .b(\u2_Display/n3155 [20]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3167 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2784 (
    .a(\u2_Display/n3131 ),
    .b(\u2_Display/n3155 [21]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3166 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2785 (
    .a(\u2_Display/n3130 ),
    .b(\u2_Display/n3155 [22]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3165 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2786 (
    .a(\u2_Display/n3129 ),
    .b(\u2_Display/n3155 [23]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3164 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2787 (
    .a(\u2_Display/n3128 ),
    .b(\u2_Display/n3155 [24]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3163 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2788 (
    .a(\u2_Display/n3127 ),
    .b(\u2_Display/n3155 [25]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3162 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2789 (
    .a(\u2_Display/n3126 ),
    .b(\u2_Display/n3155 [26]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3161 ));
  EG_PHY_PAD #(
    //.LOCATION("P8"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u279 (
    .ipad(on_off[7]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2790 (
    .a(\u2_Display/n3125 ),
    .b(\u2_Display/n3155 [27]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3160 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2791 (
    .a(\u2_Display/n3124 ),
    .b(\u2_Display/n3155 [28]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3159 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2792 (
    .a(\u2_Display/n3123 ),
    .b(\u2_Display/n3155 [29]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3158 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2793 (
    .a(\u2_Display/n3122 ),
    .b(\u2_Display/n3155 [30]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3157 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2794 (
    .a(\u2_Display/n3121 ),
    .b(\u2_Display/n3155 [31]),
    .c(\u2_Display/n3153 ),
    .o(\u2_Display/n3156 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2795 (
    .a(\u2_Display/n4310 ),
    .b(\u2_Display/n4313 [0]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4345 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2796 (
    .a(\u2_Display/n4309 ),
    .b(\u2_Display/n4313 [1]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4344 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2797 (
    .a(\u2_Display/n4308 ),
    .b(\u2_Display/n4313 [2]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4343 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2798 (
    .a(\u2_Display/n4307 ),
    .b(\u2_Display/n4313 [3]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4342 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2799 (
    .a(\u2_Display/n4306 ),
    .b(\u2_Display/n4313 [4]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4341 ));
  EG_PHY_PAD #(
    //.LOCATION("N6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u280 (
    .ipad(on_off[6]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2800 (
    .a(\u2_Display/n4305 ),
    .b(\u2_Display/n4313 [5]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4340 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2801 (
    .a(\u2_Display/n4304 ),
    .b(\u2_Display/n4313 [6]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4339 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2802 (
    .a(\u2_Display/n4303 ),
    .b(\u2_Display/n4313 [7]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4338 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2803 (
    .a(\u2_Display/n4302 ),
    .b(\u2_Display/n4313 [8]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4337 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2804 (
    .a(\u2_Display/n4301 ),
    .b(\u2_Display/n4313 [9]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4336 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2805 (
    .a(\u2_Display/n4300 ),
    .b(\u2_Display/n4313 [10]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4335 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2806 (
    .a(\u2_Display/n4299 ),
    .b(\u2_Display/n4313 [11]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4334 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2807 (
    .a(\u2_Display/n4298 ),
    .b(\u2_Display/n4313 [12]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4333 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2808 (
    .a(\u2_Display/n4297 ),
    .b(\u2_Display/n4313 [13]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4332 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2809 (
    .a(\u2_Display/n4296 ),
    .b(\u2_Display/n4313 [14]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4331 ));
  EG_PHY_PAD #(
    //.LOCATION("P6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u281 (
    .ipad(on_off[5]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2810 (
    .a(\u2_Display/n4295 ),
    .b(\u2_Display/n4313 [15]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4330 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2811 (
    .a(\u2_Display/n4294 ),
    .b(\u2_Display/n4313 [16]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4329 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2812 (
    .a(\u2_Display/n4293 ),
    .b(\u2_Display/n4313 [17]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4328 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2813 (
    .a(\u2_Display/n4292 ),
    .b(\u2_Display/n4313 [18]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4327 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2814 (
    .a(\u2_Display/n4291 ),
    .b(\u2_Display/n4313 [19]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4326 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2815 (
    .a(\u2_Display/n4290 ),
    .b(\u2_Display/n4313 [20]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4325 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2816 (
    .a(\u2_Display/n4289 ),
    .b(\u2_Display/n4313 [21]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4324 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2817 (
    .a(\u2_Display/n4288 ),
    .b(\u2_Display/n4313 [22]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4323 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2818 (
    .a(\u2_Display/n4287 ),
    .b(\u2_Display/n4313 [23]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4322 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2819 (
    .a(\u2_Display/n4286 ),
    .b(\u2_Display/n4313 [24]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4321 ));
  EG_PHY_PAD #(
    //.LOCATION("M6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u282 (
    .ipad(on_off[4]),
    .di(on_off_pad[4]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2820 (
    .a(\u2_Display/n4285 ),
    .b(\u2_Display/n4313 [25]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4320 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2821 (
    .a(\u2_Display/n4284 ),
    .b(\u2_Display/n4313 [26]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4319 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2822 (
    .a(\u2_Display/n4283 ),
    .b(\u2_Display/n4313 [27]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4318 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2823 (
    .a(\u2_Display/n4282 ),
    .b(\u2_Display/n4313 [28]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4317 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2824 (
    .a(\u2_Display/n4281 ),
    .b(\u2_Display/n4313 [29]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4316 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2825 (
    .a(\u2_Display/n4280 ),
    .b(\u2_Display/n4313 [30]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4315 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2826 (
    .a(\u2_Display/n4279 ),
    .b(\u2_Display/n4313 [31]),
    .c(\u2_Display/n4311 ),
    .o(\u2_Display/n4314 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2827 (
    .a(\u2_Display/n5433 ),
    .b(\u2_Display/n5436 [0]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5468 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2828 (
    .a(\u2_Display/n5432 ),
    .b(\u2_Display/n5436 [1]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5467 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2829 (
    .a(\u2_Display/n5431 ),
    .b(\u2_Display/n5436 [2]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5466 ));
  EG_PHY_PAD #(
    //.LOCATION("T6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u283 (
    .ipad(on_off[3]),
    .di(on_off_pad[3]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2830 (
    .a(\u2_Display/n5430 ),
    .b(\u2_Display/n5436 [3]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5465 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2831 (
    .a(\u2_Display/n5429 ),
    .b(\u2_Display/n5436 [4]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5464 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2832 (
    .a(\u2_Display/n5428 ),
    .b(\u2_Display/n5436 [5]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5463 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2833 (
    .a(\u2_Display/n5427 ),
    .b(\u2_Display/n5436 [6]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5462 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2834 (
    .a(\u2_Display/n5426 ),
    .b(\u2_Display/n5436 [7]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5461 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2835 (
    .a(\u2_Display/n5425 ),
    .b(\u2_Display/n5436 [8]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5460 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2836 (
    .a(\u2_Display/n5424 ),
    .b(\u2_Display/n5436 [9]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5459 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2837 (
    .a(\u2_Display/n5423 ),
    .b(\u2_Display/n5436 [10]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5458 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2838 (
    .a(\u2_Display/n5422 ),
    .b(\u2_Display/n5436 [11]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5457 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2839 (
    .a(\u2_Display/n5421 ),
    .b(\u2_Display/n5436 [12]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5456 ));
  EG_PHY_PAD #(
    //.LOCATION("T5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u284 (
    .ipad(on_off[2]),
    .di(on_off_pad[2]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2840 (
    .a(\u2_Display/n5420 ),
    .b(\u2_Display/n5436 [13]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5455 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2841 (
    .a(\u2_Display/n5419 ),
    .b(\u2_Display/n5436 [14]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5454 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2842 (
    .a(\u2_Display/n5418 ),
    .b(\u2_Display/n5436 [15]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5453 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2843 (
    .a(\u2_Display/n5417 ),
    .b(\u2_Display/n5436 [16]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5452 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2844 (
    .a(\u2_Display/n5416 ),
    .b(\u2_Display/n5436 [17]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5451 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2845 (
    .a(\u2_Display/n5415 ),
    .b(\u2_Display/n5436 [18]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5450 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2846 (
    .a(\u2_Display/n5414 ),
    .b(\u2_Display/n5436 [19]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5449 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2847 (
    .a(\u2_Display/n5413 ),
    .b(\u2_Display/n5436 [20]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5448 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2848 (
    .a(\u2_Display/n5412 ),
    .b(\u2_Display/n5436 [21]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5447 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2849 (
    .a(\u2_Display/n5411 ),
    .b(\u2_Display/n5436 [22]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5446 ));
  EG_PHY_PAD #(
    //.LOCATION("R5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u285 (
    .ipad(on_off[1]),
    .di(on_off_pad[1]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2850 (
    .a(\u2_Display/n5410 ),
    .b(\u2_Display/n5436 [23]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5445 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2851 (
    .a(\u2_Display/n5409 ),
    .b(\u2_Display/n5436 [24]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5444 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2852 (
    .a(\u2_Display/n5408 ),
    .b(\u2_Display/n5436 [25]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5443 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2853 (
    .a(\u2_Display/n5407 ),
    .b(\u2_Display/n5436 [26]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5442 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2854 (
    .a(\u2_Display/n5406 ),
    .b(\u2_Display/n5436 [27]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5441 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2855 (
    .a(\u2_Display/n5405 ),
    .b(\u2_Display/n5436 [28]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5440 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2856 (
    .a(\u2_Display/n5404 ),
    .b(\u2_Display/n5436 [29]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5439 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2857 (
    .a(\u2_Display/n5403 ),
    .b(\u2_Display/n5436 [30]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5438 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2858 (
    .a(\u2_Display/n5402 ),
    .b(\u2_Display/n5436 [31]),
    .c(\u2_Display/n5434 ),
    .o(\u2_Display/n5437 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2859 (
    .a(\u2_Display/n941 ),
    .b(\u2_Display/n944 [0]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n976 ));
  EG_PHY_PAD #(
    //.LOCATION("T4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u286 (
    .ipad(on_off[0]),
    .di(on_off_pad[0]));  // source/rtl/VGA_Demo.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2860 (
    .a(\u2_Display/n940 ),
    .b(\u2_Display/n944 [1]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n975 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2861 (
    .a(\u2_Display/n939 ),
    .b(\u2_Display/n944 [2]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n974 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2862 (
    .a(\u2_Display/n938 ),
    .b(\u2_Display/n944 [3]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n973 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2863 (
    .a(\u2_Display/n937 ),
    .b(\u2_Display/n944 [4]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n972 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2864 (
    .a(\u2_Display/n936 ),
    .b(\u2_Display/n944 [5]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n971 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2865 (
    .a(\u2_Display/n935 ),
    .b(\u2_Display/n944 [6]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n970 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2866 (
    .a(\u2_Display/n934 ),
    .b(\u2_Display/n944 [7]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n969 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2867 (
    .a(\u2_Display/n933 ),
    .b(\u2_Display/n944 [8]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n968 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2868 (
    .a(\u2_Display/n932 ),
    .b(\u2_Display/n944 [9]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n967 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2869 (
    .a(\u2_Display/n931 ),
    .b(\u2_Display/n944 [10]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n966 ));
  EG_PHY_PAD #(
    //.LOCATION("G11"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u287 (
    .ipad(rst_n),
    .di(rst_n_pad));  // source/rtl/VGA_Demo.v(5)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2870 (
    .a(\u2_Display/n930 ),
    .b(\u2_Display/n944 [11]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n965 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2871 (
    .a(\u2_Display/n929 ),
    .b(\u2_Display/n944 [12]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n964 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2872 (
    .a(\u2_Display/n928 ),
    .b(\u2_Display/n944 [13]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n963 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2873 (
    .a(\u2_Display/n927 ),
    .b(\u2_Display/n944 [14]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n962 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2874 (
    .a(\u2_Display/n926 ),
    .b(\u2_Display/n944 [15]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n961 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2875 (
    .a(\u2_Display/n925 ),
    .b(\u2_Display/n944 [16]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n960 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2876 (
    .a(\u2_Display/n924 ),
    .b(\u2_Display/n944 [17]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n959 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2877 (
    .a(\u2_Display/n923 ),
    .b(\u2_Display/n944 [18]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n958 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2878 (
    .a(\u2_Display/n922 ),
    .b(\u2_Display/n944 [19]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n957 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2879 (
    .a(\u2_Display/n921 ),
    .b(\u2_Display/n944 [20]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n956 ));
  EG_PHY_PAD #(
    //.LOCATION("C1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u288 (
    .do({open_n174,open_n175,open_n176,vga_b_pad[0]}),
    .opad(vga_b[7]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2880 (
    .a(\u2_Display/n920 ),
    .b(\u2_Display/n944 [21]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n955 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2881 (
    .a(\u2_Display/n919 ),
    .b(\u2_Display/n944 [22]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n954 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2882 (
    .a(\u2_Display/n918 ),
    .b(\u2_Display/n944 [23]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n953 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2883 (
    .a(\u2_Display/n917 ),
    .b(\u2_Display/n944 [24]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n952 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2884 (
    .a(\u2_Display/n916 ),
    .b(\u2_Display/n944 [25]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n951 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2885 (
    .a(\u2_Display/n915 ),
    .b(\u2_Display/n944 [26]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n950 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2886 (
    .a(\u2_Display/n914 ),
    .b(\u2_Display/n944 [27]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n949 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2887 (
    .a(\u2_Display/n913 ),
    .b(\u2_Display/n944 [28]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n948 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2888 (
    .a(\u2_Display/n912 ),
    .b(\u2_Display/n944 [29]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n947 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2889 (
    .a(\u2_Display/n911 ),
    .b(\u2_Display/n944 [30]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n946 ));
  EG_PHY_PAD #(
    //.LOCATION("D1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u289 (
    .do({open_n191,open_n192,open_n193,vga_b_pad[0]}),
    .opad(vga_b[6]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2890 (
    .a(\u2_Display/n910 ),
    .b(\u2_Display/n944 [31]),
    .c(\u2_Display/n942 ),
    .o(\u2_Display/n945 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2891 (
    .a(\u2_Display/n2064 ),
    .b(\u2_Display/n2067 [0]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2099 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2892 (
    .a(\u2_Display/n2063 ),
    .b(\u2_Display/n2067 [1]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2098 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2893 (
    .a(\u2_Display/n2062 ),
    .b(\u2_Display/n2067 [2]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2097 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2894 (
    .a(\u2_Display/n2061 ),
    .b(\u2_Display/n2067 [3]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2096 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2895 (
    .a(\u2_Display/n2060 ),
    .b(\u2_Display/n2067 [4]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2095 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2896 (
    .a(\u2_Display/n2059 ),
    .b(\u2_Display/n2067 [5]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2094 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2897 (
    .a(\u2_Display/n2058 ),
    .b(\u2_Display/n2067 [6]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2093 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2898 (
    .a(\u2_Display/n2057 ),
    .b(\u2_Display/n2067 [7]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2092 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2899 (
    .a(\u2_Display/n2056 ),
    .b(\u2_Display/n2067 [8]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2091 ));
  EG_PHY_PAD #(
    //.LOCATION("E2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u290 (
    .do({open_n208,open_n209,open_n210,vga_b_pad[0]}),
    .opad(vga_b[5]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2900 (
    .a(\u2_Display/n2055 ),
    .b(\u2_Display/n2067 [9]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2090 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2901 (
    .a(\u2_Display/n2054 ),
    .b(\u2_Display/n2067 [10]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2089 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2902 (
    .a(\u2_Display/n2053 ),
    .b(\u2_Display/n2067 [11]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2088 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2903 (
    .a(\u2_Display/n2052 ),
    .b(\u2_Display/n2067 [12]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2087 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2904 (
    .a(\u2_Display/n2051 ),
    .b(\u2_Display/n2067 [13]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2086 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2905 (
    .a(\u2_Display/n2050 ),
    .b(\u2_Display/n2067 [14]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2085 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2906 (
    .a(\u2_Display/n2049 ),
    .b(\u2_Display/n2067 [15]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2084 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2907 (
    .a(\u2_Display/n2048 ),
    .b(\u2_Display/n2067 [16]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2083 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2908 (
    .a(\u2_Display/n2047 ),
    .b(\u2_Display/n2067 [17]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2082 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2909 (
    .a(\u2_Display/n2046 ),
    .b(\u2_Display/n2067 [18]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2081 ));
  EG_PHY_PAD #(
    //.LOCATION("G3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u291 (
    .do({open_n225,open_n226,open_n227,vga_b_pad[0]}),
    .opad(vga_b[4]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2910 (
    .a(\u2_Display/n2045 ),
    .b(\u2_Display/n2067 [19]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2080 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2911 (
    .a(\u2_Display/n2044 ),
    .b(\u2_Display/n2067 [20]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2079 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2912 (
    .a(\u2_Display/n2043 ),
    .b(\u2_Display/n2067 [21]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2078 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2913 (
    .a(\u2_Display/n2042 ),
    .b(\u2_Display/n2067 [22]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2077 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2914 (
    .a(\u2_Display/n2041 ),
    .b(\u2_Display/n2067 [23]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2076 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2915 (
    .a(\u2_Display/n2040 ),
    .b(\u2_Display/n2067 [24]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2075 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2916 (
    .a(\u2_Display/n2039 ),
    .b(\u2_Display/n2067 [25]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2074 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2917 (
    .a(\u2_Display/n2038 ),
    .b(\u2_Display/n2067 [26]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2073 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2918 (
    .a(\u2_Display/n2037 ),
    .b(\u2_Display/n2067 [27]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2072 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2919 (
    .a(\u2_Display/n2036 ),
    .b(\u2_Display/n2067 [28]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2071 ));
  EG_PHY_PAD #(
    //.LOCATION("E1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u292 (
    .do({open_n242,open_n243,open_n244,vga_b_pad[0]}),
    .opad(vga_b[3]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2920 (
    .a(\u2_Display/n2035 ),
    .b(\u2_Display/n2067 [29]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2070 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2921 (
    .a(\u2_Display/n2034 ),
    .b(\u2_Display/n2067 [30]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2069 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2922 (
    .a(\u2_Display/n2033 ),
    .b(\u2_Display/n2067 [31]),
    .c(\u2_Display/n2065 ),
    .o(\u2_Display/n2068 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2923 (
    .a(\u2_Display/n3187 ),
    .b(\u2_Display/n3190 [0]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3222 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2924 (
    .a(\u2_Display/n3186 ),
    .b(\u2_Display/n3190 [1]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3221 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2925 (
    .a(\u2_Display/n3185 ),
    .b(\u2_Display/n3190 [2]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3220 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2926 (
    .a(\u2_Display/n3184 ),
    .b(\u2_Display/n3190 [3]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3219 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2927 (
    .a(\u2_Display/n3183 ),
    .b(\u2_Display/n3190 [4]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3218 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2928 (
    .a(\u2_Display/n3182 ),
    .b(\u2_Display/n3190 [5]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3217 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2929 (
    .a(\u2_Display/n3181 ),
    .b(\u2_Display/n3190 [6]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3216 ));
  EG_PHY_PAD #(
    //.LOCATION("F2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u293 (
    .do({open_n259,open_n260,open_n261,vga_b_pad[0]}),
    .opad(vga_b[2]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2930 (
    .a(\u2_Display/n3180 ),
    .b(\u2_Display/n3190 [7]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3215 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2931 (
    .a(\u2_Display/n3179 ),
    .b(\u2_Display/n3190 [8]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3214 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2932 (
    .a(\u2_Display/n3178 ),
    .b(\u2_Display/n3190 [9]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3213 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2933 (
    .a(\u2_Display/n3177 ),
    .b(\u2_Display/n3190 [10]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3212 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2934 (
    .a(\u2_Display/n3176 ),
    .b(\u2_Display/n3190 [11]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3211 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2935 (
    .a(\u2_Display/n3175 ),
    .b(\u2_Display/n3190 [12]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3210 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2936 (
    .a(\u2_Display/n3174 ),
    .b(\u2_Display/n3190 [13]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3209 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2937 (
    .a(\u2_Display/n3173 ),
    .b(\u2_Display/n3190 [14]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3208 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2938 (
    .a(\u2_Display/n3172 ),
    .b(\u2_Display/n3190 [15]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3207 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2939 (
    .a(\u2_Display/n3171 ),
    .b(\u2_Display/n3190 [16]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3206 ));
  EG_PHY_PAD #(
    //.LOCATION("F1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u294 (
    .do({open_n276,open_n277,open_n278,vga_b_pad[0]}),
    .opad(vga_b[1]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2940 (
    .a(\u2_Display/n3170 ),
    .b(\u2_Display/n3190 [17]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3205 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2941 (
    .a(\u2_Display/n3169 ),
    .b(\u2_Display/n3190 [18]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3204 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2942 (
    .a(\u2_Display/n3168 ),
    .b(\u2_Display/n3190 [19]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3203 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2943 (
    .a(\u2_Display/n3167 ),
    .b(\u2_Display/n3190 [20]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3202 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2944 (
    .a(\u2_Display/n3166 ),
    .b(\u2_Display/n3190 [21]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3201 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2945 (
    .a(\u2_Display/n3165 ),
    .b(\u2_Display/n3190 [22]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3200 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2946 (
    .a(\u2_Display/n3164 ),
    .b(\u2_Display/n3190 [23]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3199 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2947 (
    .a(\u2_Display/n3163 ),
    .b(\u2_Display/n3190 [24]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3198 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2948 (
    .a(\u2_Display/n3162 ),
    .b(\u2_Display/n3190 [25]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3197 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2949 (
    .a(\u2_Display/n3161 ),
    .b(\u2_Display/n3190 [26]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3196 ));
  EG_PHY_PAD #(
    //.LOCATION("G1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u295 (
    .do({open_n293,open_n294,open_n295,vga_b_pad[0]}),
    .opad(vga_b[0]));  // source/rtl/VGA_Demo.v(17)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2950 (
    .a(\u2_Display/n3160 ),
    .b(\u2_Display/n3190 [27]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3195 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2951 (
    .a(\u2_Display/n3159 ),
    .b(\u2_Display/n3190 [28]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3194 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2952 (
    .a(\u2_Display/n3158 ),
    .b(\u2_Display/n3190 [29]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3193 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2953 (
    .a(\u2_Display/n3157 ),
    .b(\u2_Display/n3190 [30]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3192 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2954 (
    .a(\u2_Display/n3156 ),
    .b(\u2_Display/n3190 [31]),
    .c(\u2_Display/n3188 ),
    .o(\u2_Display/n3191 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2955 (
    .a(\u2_Display/n4345 ),
    .b(\u2_Display/n4348 [0]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4380 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2956 (
    .a(\u2_Display/n4344 ),
    .b(\u2_Display/n4348 [1]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4379 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2957 (
    .a(\u2_Display/n4343 ),
    .b(\u2_Display/n4348 [2]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4378 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2958 (
    .a(\u2_Display/n4342 ),
    .b(\u2_Display/n4348 [3]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4377 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2959 (
    .a(\u2_Display/n4341 ),
    .b(\u2_Display/n4348 [4]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4376 ));
  EG_PHY_PAD #(
    //.LOCATION("H2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u296 (
    .do({open_n310,open_n311,open_n312,vga_clk_pad}),
    .opad(vga_clk));  // source/rtl/VGA_Demo.v(9)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2960 (
    .a(\u2_Display/n4340 ),
    .b(\u2_Display/n4348 [5]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4375 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2961 (
    .a(\u2_Display/n4339 ),
    .b(\u2_Display/n4348 [6]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4374 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2962 (
    .a(\u2_Display/n4338 ),
    .b(\u2_Display/n4348 [7]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4373 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2963 (
    .a(\u2_Display/n4337 ),
    .b(\u2_Display/n4348 [8]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4372 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2964 (
    .a(\u2_Display/n4336 ),
    .b(\u2_Display/n4348 [9]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4371 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2965 (
    .a(\u2_Display/n4335 ),
    .b(\u2_Display/n4348 [10]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4370 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2966 (
    .a(\u2_Display/n4334 ),
    .b(\u2_Display/n4348 [11]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4369 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2967 (
    .a(\u2_Display/n4333 ),
    .b(\u2_Display/n4348 [12]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4368 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2968 (
    .a(\u2_Display/n4332 ),
    .b(\u2_Display/n4348 [13]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4367 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2969 (
    .a(\u2_Display/n4331 ),
    .b(\u2_Display/n4348 [14]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4366 ));
  EG_PHY_PAD #(
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u297 (
    .do({open_n327,open_n328,open_n329,vga_de_pad}),
    .opad(vga_de));  // source/rtl/VGA_Demo.v(13)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2970 (
    .a(\u2_Display/n4330 ),
    .b(\u2_Display/n4348 [15]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4365 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2971 (
    .a(\u2_Display/n4329 ),
    .b(\u2_Display/n4348 [16]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4364 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2972 (
    .a(\u2_Display/n4328 ),
    .b(\u2_Display/n4348 [17]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4363 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2973 (
    .a(\u2_Display/n4327 ),
    .b(\u2_Display/n4348 [18]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4362 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2974 (
    .a(\u2_Display/n4326 ),
    .b(\u2_Display/n4348 [19]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4361 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2975 (
    .a(\u2_Display/n4325 ),
    .b(\u2_Display/n4348 [20]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4360 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2976 (
    .a(\u2_Display/n4324 ),
    .b(\u2_Display/n4348 [21]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4359 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2977 (
    .a(\u2_Display/n4323 ),
    .b(\u2_Display/n4348 [22]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4358 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2978 (
    .a(\u2_Display/n4322 ),
    .b(\u2_Display/n4348 [23]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4357 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2979 (
    .a(\u2_Display/n4321 ),
    .b(\u2_Display/n4348 [24]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4356 ));
  EG_PHY_PAD #(
    //.LOCATION("H5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u298 (
    .do({open_n344,open_n345,open_n346,vga_b_pad[0]}),
    .opad(vga_g[7]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2980 (
    .a(\u2_Display/n4320 ),
    .b(\u2_Display/n4348 [25]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4355 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2981 (
    .a(\u2_Display/n4319 ),
    .b(\u2_Display/n4348 [26]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4354 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2982 (
    .a(\u2_Display/n4318 ),
    .b(\u2_Display/n4348 [27]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4353 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2983 (
    .a(\u2_Display/n4317 ),
    .b(\u2_Display/n4348 [28]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4352 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2984 (
    .a(\u2_Display/n4316 ),
    .b(\u2_Display/n4348 [29]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4351 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2985 (
    .a(\u2_Display/n4315 ),
    .b(\u2_Display/n4348 [30]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4350 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2986 (
    .a(\u2_Display/n4314 ),
    .b(\u2_Display/n4348 [31]),
    .c(\u2_Display/n4346 ),
    .o(\u2_Display/n4349 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2987 (
    .a(\u2_Display/n5468 ),
    .b(\u2_Display/n5471 [0]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5503 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2988 (
    .a(\u2_Display/n5467 ),
    .b(\u2_Display/n5471 [1]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5502 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2989 (
    .a(\u2_Display/n5466 ),
    .b(\u2_Display/n5471 [2]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5501 ));
  EG_PHY_PAD #(
    //.LOCATION("H1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u299 (
    .do({open_n361,open_n362,open_n363,vga_b_pad[0]}),
    .opad(vga_g[6]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2990 (
    .a(\u2_Display/n5465 ),
    .b(\u2_Display/n5471 [3]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5500 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2991 (
    .a(\u2_Display/n5464 ),
    .b(\u2_Display/n5471 [4]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5499 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2992 (
    .a(\u2_Display/n5463 ),
    .b(\u2_Display/n5471 [5]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5498 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2993 (
    .a(\u2_Display/n5462 ),
    .b(\u2_Display/n5471 [6]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5497 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2994 (
    .a(\u2_Display/n5461 ),
    .b(\u2_Display/n5471 [7]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5496 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2995 (
    .a(\u2_Display/n5460 ),
    .b(\u2_Display/n5471 [8]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5495 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2996 (
    .a(\u2_Display/n5459 ),
    .b(\u2_Display/n5471 [9]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5494 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2997 (
    .a(\u2_Display/n5458 ),
    .b(\u2_Display/n5471 [10]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5493 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2998 (
    .a(\u2_Display/n5457 ),
    .b(\u2_Display/n5471 [11]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5492 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u2999 (
    .a(\u2_Display/n5456 ),
    .b(\u2_Display/n5471 [12]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5491 ));
  EG_PHY_PAD #(
    //.LOCATION("J6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u300 (
    .do({open_n378,open_n379,open_n380,vga_b_pad[0]}),
    .opad(vga_g[5]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3000 (
    .a(\u2_Display/n5455 ),
    .b(\u2_Display/n5471 [13]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5490 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3001 (
    .a(\u2_Display/n5454 ),
    .b(\u2_Display/n5471 [14]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5489 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3002 (
    .a(\u2_Display/n5453 ),
    .b(\u2_Display/n5471 [15]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5488 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3003 (
    .a(\u2_Display/n5452 ),
    .b(\u2_Display/n5471 [16]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5487 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3004 (
    .a(\u2_Display/n5451 ),
    .b(\u2_Display/n5471 [17]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5486 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3005 (
    .a(\u2_Display/n5450 ),
    .b(\u2_Display/n5471 [18]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5485 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3006 (
    .a(\u2_Display/n5449 ),
    .b(\u2_Display/n5471 [19]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5484 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3007 (
    .a(\u2_Display/n5448 ),
    .b(\u2_Display/n5471 [20]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5483 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3008 (
    .a(\u2_Display/n5447 ),
    .b(\u2_Display/n5471 [21]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5482 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3009 (
    .a(\u2_Display/n5446 ),
    .b(\u2_Display/n5471 [22]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5481 ));
  EG_PHY_PAD #(
    //.LOCATION("H3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u301 (
    .do({open_n395,open_n396,open_n397,vga_b_pad[0]}),
    .opad(vga_g[4]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3010 (
    .a(\u2_Display/n5445 ),
    .b(\u2_Display/n5471 [23]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5480 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3011 (
    .a(\u2_Display/n5444 ),
    .b(\u2_Display/n5471 [24]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5479 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3012 (
    .a(\u2_Display/n5443 ),
    .b(\u2_Display/n5471 [25]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5478 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3013 (
    .a(\u2_Display/n5442 ),
    .b(\u2_Display/n5471 [26]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5477 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3014 (
    .a(\u2_Display/n5441 ),
    .b(\u2_Display/n5471 [27]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5476 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3015 (
    .a(\u2_Display/n5440 ),
    .b(\u2_Display/n5471 [28]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5475 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3016 (
    .a(\u2_Display/n5439 ),
    .b(\u2_Display/n5471 [29]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5474 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3017 (
    .a(\u2_Display/n5438 ),
    .b(\u2_Display/n5471 [30]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5473 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3018 (
    .a(\u2_Display/n5437 ),
    .b(\u2_Display/n5471 [31]),
    .c(\u2_Display/n5469 ),
    .o(\u2_Display/n5472 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3019 (
    .a(\u2_Display/n976 ),
    .b(\u2_Display/n979 [0]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1011 ));
  EG_PHY_PAD #(
    //.LOCATION("J1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u302 (
    .do({open_n412,open_n413,open_n414,vga_b_pad[0]}),
    .opad(vga_g[3]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3020 (
    .a(\u2_Display/n975 ),
    .b(\u2_Display/n979 [1]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1010 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3021 (
    .a(\u2_Display/n974 ),
    .b(\u2_Display/n979 [2]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1009 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3022 (
    .a(\u2_Display/n973 ),
    .b(\u2_Display/n979 [3]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1008 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3023 (
    .a(\u2_Display/n972 ),
    .b(\u2_Display/n979 [4]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1007 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3024 (
    .a(\u2_Display/n971 ),
    .b(\u2_Display/n979 [5]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1006 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3025 (
    .a(\u2_Display/n970 ),
    .b(\u2_Display/n979 [6]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1005 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3026 (
    .a(\u2_Display/n969 ),
    .b(\u2_Display/n979 [7]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1004 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3027 (
    .a(\u2_Display/n968 ),
    .b(\u2_Display/n979 [8]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1003 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3028 (
    .a(\u2_Display/n967 ),
    .b(\u2_Display/n979 [9]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1002 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3029 (
    .a(\u2_Display/n966 ),
    .b(\u2_Display/n979 [10]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1001 ));
  EG_PHY_PAD #(
    //.LOCATION("K1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u303 (
    .do({open_n429,open_n430,open_n431,vga_b_pad[0]}),
    .opad(vga_g[2]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3030 (
    .a(\u2_Display/n965 ),
    .b(\u2_Display/n979 [11]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n1000 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3031 (
    .a(\u2_Display/n964 ),
    .b(\u2_Display/n979 [12]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n999 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3032 (
    .a(\u2_Display/n963 ),
    .b(\u2_Display/n979 [13]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n998 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3033 (
    .a(\u2_Display/n962 ),
    .b(\u2_Display/n979 [14]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n997 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3034 (
    .a(\u2_Display/n961 ),
    .b(\u2_Display/n979 [15]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n996 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3035 (
    .a(\u2_Display/n960 ),
    .b(\u2_Display/n979 [16]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n995 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3036 (
    .a(\u2_Display/n959 ),
    .b(\u2_Display/n979 [17]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n994 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3037 (
    .a(\u2_Display/n958 ),
    .b(\u2_Display/n979 [18]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n993 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3038 (
    .a(\u2_Display/n957 ),
    .b(\u2_Display/n979 [19]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n992 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3039 (
    .a(\u2_Display/n956 ),
    .b(\u2_Display/n979 [20]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n991 ));
  EG_PHY_PAD #(
    //.LOCATION("K2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u304 (
    .do({open_n446,open_n447,open_n448,vga_b_pad[0]}),
    .opad(vga_g[1]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3040 (
    .a(\u2_Display/n955 ),
    .b(\u2_Display/n979 [21]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n990 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3041 (
    .a(\u2_Display/n954 ),
    .b(\u2_Display/n979 [22]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n989 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3042 (
    .a(\u2_Display/n953 ),
    .b(\u2_Display/n979 [23]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n988 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3043 (
    .a(\u2_Display/n952 ),
    .b(\u2_Display/n979 [24]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n987 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3044 (
    .a(\u2_Display/n951 ),
    .b(\u2_Display/n979 [25]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n986 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3045 (
    .a(\u2_Display/n950 ),
    .b(\u2_Display/n979 [26]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n985 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3046 (
    .a(\u2_Display/n949 ),
    .b(\u2_Display/n979 [27]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n984 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3047 (
    .a(\u2_Display/n948 ),
    .b(\u2_Display/n979 [28]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n983 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3048 (
    .a(\u2_Display/n947 ),
    .b(\u2_Display/n979 [29]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n982 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3049 (
    .a(\u2_Display/n946 ),
    .b(\u2_Display/n979 [30]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n981 ));
  EG_PHY_PAD #(
    //.LOCATION("L1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u305 (
    .do({open_n463,open_n464,open_n465,vga_b_pad[0]}),
    .opad(vga_g[0]));  // source/rtl/VGA_Demo.v(16)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3050 (
    .a(\u2_Display/n945 ),
    .b(\u2_Display/n979 [31]),
    .c(\u2_Display/n977 ),
    .o(\u2_Display/n980 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3051 (
    .a(\u2_Display/n2099 ),
    .b(\u2_Display/n2102 [0]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2134 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3052 (
    .a(\u2_Display/n2098 ),
    .b(\u2_Display/n2102 [1]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2133 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3053 (
    .a(\u2_Display/n2097 ),
    .b(\u2_Display/n2102 [2]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2132 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3054 (
    .a(\u2_Display/n2096 ),
    .b(\u2_Display/n2102 [3]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2131 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3055 (
    .a(\u2_Display/n2095 ),
    .b(\u2_Display/n2102 [4]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2130 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3056 (
    .a(\u2_Display/n2094 ),
    .b(\u2_Display/n2102 [5]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2129 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3057 (
    .a(\u2_Display/n2093 ),
    .b(\u2_Display/n2102 [6]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2128 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3058 (
    .a(\u2_Display/n2092 ),
    .b(\u2_Display/n2102 [7]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2127 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3059 (
    .a(\u2_Display/n2091 ),
    .b(\u2_Display/n2102 [8]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2126 ));
  EG_PHY_PAD #(
    //.LOCATION("J3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u306 (
    .do({open_n480,open_n481,open_n482,vga_hs_pad}),
    .opad(vga_hs));  // source/rtl/VGA_Demo.v(10)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3060 (
    .a(\u2_Display/n2090 ),
    .b(\u2_Display/n2102 [9]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2125 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3061 (
    .a(\u2_Display/n2089 ),
    .b(\u2_Display/n2102 [10]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2124 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3062 (
    .a(\u2_Display/n2088 ),
    .b(\u2_Display/n2102 [11]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2123 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3063 (
    .a(\u2_Display/n2087 ),
    .b(\u2_Display/n2102 [12]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2122 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3064 (
    .a(\u2_Display/n2086 ),
    .b(\u2_Display/n2102 [13]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2121 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3065 (
    .a(\u2_Display/n2085 ),
    .b(\u2_Display/n2102 [14]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2120 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3066 (
    .a(\u2_Display/n2084 ),
    .b(\u2_Display/n2102 [15]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2119 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3067 (
    .a(\u2_Display/n2083 ),
    .b(\u2_Display/n2102 [16]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2118 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3068 (
    .a(\u2_Display/n2082 ),
    .b(\u2_Display/n2102 [17]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2117 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3069 (
    .a(\u2_Display/n2081 ),
    .b(\u2_Display/n2102 [18]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2116 ));
  EG_PHY_PAD #(
    //.LOCATION("K6"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u307 (
    .do({open_n497,open_n498,open_n499,vga_b_pad[0]}),
    .opad(vga_r[7]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3070 (
    .a(\u2_Display/n2080 ),
    .b(\u2_Display/n2102 [19]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2115 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3071 (
    .a(\u2_Display/n2079 ),
    .b(\u2_Display/n2102 [20]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2114 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3072 (
    .a(\u2_Display/n2078 ),
    .b(\u2_Display/n2102 [21]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2113 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3073 (
    .a(\u2_Display/n2077 ),
    .b(\u2_Display/n2102 [22]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2112 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3074 (
    .a(\u2_Display/n2076 ),
    .b(\u2_Display/n2102 [23]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2111 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3075 (
    .a(\u2_Display/n2075 ),
    .b(\u2_Display/n2102 [24]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2110 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3076 (
    .a(\u2_Display/n2074 ),
    .b(\u2_Display/n2102 [25]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2109 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3077 (
    .a(\u2_Display/n2073 ),
    .b(\u2_Display/n2102 [26]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2108 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3078 (
    .a(\u2_Display/n2072 ),
    .b(\u2_Display/n2102 [27]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2107 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3079 (
    .a(\u2_Display/n2071 ),
    .b(\u2_Display/n2102 [28]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2106 ));
  EG_PHY_PAD #(
    //.LOCATION("K3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u308 (
    .do({open_n514,open_n515,open_n516,vga_b_pad[0]}),
    .opad(vga_r[6]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3080 (
    .a(\u2_Display/n2070 ),
    .b(\u2_Display/n2102 [29]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2105 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3081 (
    .a(\u2_Display/n2069 ),
    .b(\u2_Display/n2102 [30]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2104 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3082 (
    .a(\u2_Display/n2068 ),
    .b(\u2_Display/n2102 [31]),
    .c(\u2_Display/n2100 ),
    .o(\u2_Display/n2103 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3083 (
    .a(\u2_Display/n3222 ),
    .b(\u2_Display/n3225 [0]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3257 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3084 (
    .a(\u2_Display/n3221 ),
    .b(\u2_Display/n3225 [1]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3256 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3085 (
    .a(\u2_Display/n3220 ),
    .b(\u2_Display/n3225 [2]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3255 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3086 (
    .a(\u2_Display/n3219 ),
    .b(\u2_Display/n3225 [3]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3254 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3087 (
    .a(\u2_Display/n3218 ),
    .b(\u2_Display/n3225 [4]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3253 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3088 (
    .a(\u2_Display/n3217 ),
    .b(\u2_Display/n3225 [5]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3252 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3089 (
    .a(\u2_Display/n3216 ),
    .b(\u2_Display/n3225 [6]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3251 ));
  EG_PHY_PAD #(
    //.LOCATION("K5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u309 (
    .do({open_n531,open_n532,open_n533,vga_b_pad[0]}),
    .opad(vga_r[5]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3090 (
    .a(\u2_Display/n3215 ),
    .b(\u2_Display/n3225 [7]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3250 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3091 (
    .a(\u2_Display/n3214 ),
    .b(\u2_Display/n3225 [8]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3249 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3092 (
    .a(\u2_Display/n3213 ),
    .b(\u2_Display/n3225 [9]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3248 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3093 (
    .a(\u2_Display/n3212 ),
    .b(\u2_Display/n3225 [10]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3247 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3094 (
    .a(\u2_Display/n3211 ),
    .b(\u2_Display/n3225 [11]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3246 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3095 (
    .a(\u2_Display/n3210 ),
    .b(\u2_Display/n3225 [12]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3245 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3096 (
    .a(\u2_Display/n3209 ),
    .b(\u2_Display/n3225 [13]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3244 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3097 (
    .a(\u2_Display/n3208 ),
    .b(\u2_Display/n3225 [14]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3243 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3098 (
    .a(\u2_Display/n3207 ),
    .b(\u2_Display/n3225 [15]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3242 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3099 (
    .a(\u2_Display/n3206 ),
    .b(\u2_Display/n3225 [16]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3241 ));
  EG_PHY_PAD #(
    //.LOCATION("L4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u310 (
    .do({open_n548,open_n549,open_n550,vga_b_pad[0]}),
    .opad(vga_r[4]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3100 (
    .a(\u2_Display/n3205 ),
    .b(\u2_Display/n3225 [17]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3240 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3101 (
    .a(\u2_Display/n3204 ),
    .b(\u2_Display/n3225 [18]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3239 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3102 (
    .a(\u2_Display/n3203 ),
    .b(\u2_Display/n3225 [19]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3238 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3103 (
    .a(\u2_Display/n3202 ),
    .b(\u2_Display/n3225 [20]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3237 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3104 (
    .a(\u2_Display/n3201 ),
    .b(\u2_Display/n3225 [21]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3236 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3105 (
    .a(\u2_Display/n3200 ),
    .b(\u2_Display/n3225 [22]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3235 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3106 (
    .a(\u2_Display/n3199 ),
    .b(\u2_Display/n3225 [23]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3234 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3107 (
    .a(\u2_Display/n3198 ),
    .b(\u2_Display/n3225 [24]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3233 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3108 (
    .a(\u2_Display/n3197 ),
    .b(\u2_Display/n3225 [25]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3232 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3109 (
    .a(\u2_Display/n3196 ),
    .b(\u2_Display/n3225 [26]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3231 ));
  EG_PHY_PAD #(
    //.LOCATION("M1"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u311 (
    .do({open_n565,open_n566,open_n567,vga_b_pad[0]}),
    .opad(vga_r[3]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3110 (
    .a(\u2_Display/n3195 ),
    .b(\u2_Display/n3225 [27]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3230 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3111 (
    .a(\u2_Display/n3194 ),
    .b(\u2_Display/n3225 [28]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3229 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3112 (
    .a(\u2_Display/n3193 ),
    .b(\u2_Display/n3225 [29]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3228 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3113 (
    .a(\u2_Display/n3192 ),
    .b(\u2_Display/n3225 [30]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3227 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3114 (
    .a(\u2_Display/n3191 ),
    .b(\u2_Display/n3225 [31]),
    .c(\u2_Display/n3223 ),
    .o(\u2_Display/n3226 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3115 (
    .a(\u2_Display/n4380 ),
    .b(\u2_Display/n4383 [0]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4415 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3116 (
    .a(\u2_Display/n4379 ),
    .b(\u2_Display/n4383 [1]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4414 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3117 (
    .a(\u2_Display/n4378 ),
    .b(\u2_Display/n4383 [2]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4413 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3118 (
    .a(\u2_Display/n4377 ),
    .b(\u2_Display/n4383 [3]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4412 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3119 (
    .a(\u2_Display/n4376 ),
    .b(\u2_Display/n4383 [4]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4411 ));
  EG_PHY_PAD #(
    //.LOCATION("M2"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u312 (
    .do({open_n582,open_n583,open_n584,vga_b_pad[0]}),
    .opad(vga_r[2]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3120 (
    .a(\u2_Display/n4375 ),
    .b(\u2_Display/n4383 [5]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4410 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3121 (
    .a(\u2_Display/n4374 ),
    .b(\u2_Display/n4383 [6]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4409 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3122 (
    .a(\u2_Display/n4373 ),
    .b(\u2_Display/n4383 [7]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4408 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3123 (
    .a(\u2_Display/n4372 ),
    .b(\u2_Display/n4383 [8]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4407 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3124 (
    .a(\u2_Display/n4371 ),
    .b(\u2_Display/n4383 [9]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4406 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3125 (
    .a(\u2_Display/n4370 ),
    .b(\u2_Display/n4383 [10]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4405 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3126 (
    .a(\u2_Display/n4369 ),
    .b(\u2_Display/n4383 [11]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4404 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3127 (
    .a(\u2_Display/n4368 ),
    .b(\u2_Display/n4383 [12]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4403 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3128 (
    .a(\u2_Display/n4367 ),
    .b(\u2_Display/n4383 [13]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4402 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3129 (
    .a(\u2_Display/n4366 ),
    .b(\u2_Display/n4383 [14]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4401 ));
  EG_PHY_PAD #(
    //.LOCATION("L3"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u313 (
    .do({open_n599,open_n600,open_n601,vga_b_pad[0]}),
    .opad(vga_r[1]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3130 (
    .a(\u2_Display/n4365 ),
    .b(\u2_Display/n4383 [15]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4400 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3131 (
    .a(\u2_Display/n4364 ),
    .b(\u2_Display/n4383 [16]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4399 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3132 (
    .a(\u2_Display/n4363 ),
    .b(\u2_Display/n4383 [17]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4398 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3133 (
    .a(\u2_Display/n4362 ),
    .b(\u2_Display/n4383 [18]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4397 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3134 (
    .a(\u2_Display/n4361 ),
    .b(\u2_Display/n4383 [19]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4396 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3135 (
    .a(\u2_Display/n4360 ),
    .b(\u2_Display/n4383 [20]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4395 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3136 (
    .a(\u2_Display/n4359 ),
    .b(\u2_Display/n4383 [21]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4394 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3137 (
    .a(\u2_Display/n4358 ),
    .b(\u2_Display/n4383 [22]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4393 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3138 (
    .a(\u2_Display/n4357 ),
    .b(\u2_Display/n4383 [23]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4392 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3139 (
    .a(\u2_Display/n4356 ),
    .b(\u2_Display/n4383 [24]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4391 ));
  EG_PHY_PAD #(
    //.LOCATION("L5"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u314 (
    .do({open_n616,open_n617,open_n618,vga_b_pad[0]}),
    .opad(vga_r[0]));  // source/rtl/VGA_Demo.v(15)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3140 (
    .a(\u2_Display/n4355 ),
    .b(\u2_Display/n4383 [25]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4390 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3141 (
    .a(\u2_Display/n4354 ),
    .b(\u2_Display/n4383 [26]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4389 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3142 (
    .a(\u2_Display/n4353 ),
    .b(\u2_Display/n4383 [27]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4388 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3143 (
    .a(\u2_Display/n4352 ),
    .b(\u2_Display/n4383 [28]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4387 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3144 (
    .a(\u2_Display/n4351 ),
    .b(\u2_Display/n4383 [29]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4386 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3145 (
    .a(\u2_Display/n4350 ),
    .b(\u2_Display/n4383 [30]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4385 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3146 (
    .a(\u2_Display/n4349 ),
    .b(\u2_Display/n4383 [31]),
    .c(\u2_Display/n4381 ),
    .o(\u2_Display/n4384 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3147 (
    .a(\u2_Display/n5503 ),
    .b(\u2_Display/n5506 [0]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5538 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3148 (
    .a(\u2_Display/n5502 ),
    .b(\u2_Display/n5506 [1]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5537 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3149 (
    .a(\u2_Display/n5501 ),
    .b(\u2_Display/n5506 [2]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5536 ));
  EG_PHY_PAD #(
    //.LOCATION("J4"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u315 (
    .do({open_n633,open_n634,open_n635,vga_vs_pad}),
    .opad(vga_vs));  // source/rtl/VGA_Demo.v(11)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3150 (
    .a(\u2_Display/n5500 ),
    .b(\u2_Display/n5506 [3]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5535 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3151 (
    .a(\u2_Display/n5499 ),
    .b(\u2_Display/n5506 [4]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5534 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3152 (
    .a(\u2_Display/n5498 ),
    .b(\u2_Display/n5506 [5]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5533 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3153 (
    .a(\u2_Display/n5497 ),
    .b(\u2_Display/n5506 [6]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5532 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3154 (
    .a(\u2_Display/n5496 ),
    .b(\u2_Display/n5506 [7]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5531 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3155 (
    .a(\u2_Display/n5495 ),
    .b(\u2_Display/n5506 [8]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5530 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3156 (
    .a(\u2_Display/n5494 ),
    .b(\u2_Display/n5506 [9]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5529 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3157 (
    .a(\u2_Display/n5493 ),
    .b(\u2_Display/n5506 [10]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5528 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3158 (
    .a(\u2_Display/n5492 ),
    .b(\u2_Display/n5506 [11]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5527 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3159 (
    .a(\u2_Display/n5491 ),
    .b(\u2_Display/n5506 [12]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5526 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u316 (
    .a(\u1_Driver/n2 [9]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3160 (
    .a(\u2_Display/n5490 ),
    .b(\u2_Display/n5506 [13]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5525 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3161 (
    .a(\u2_Display/n5489 ),
    .b(\u2_Display/n5506 [14]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5524 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3162 (
    .a(\u2_Display/n5488 ),
    .b(\u2_Display/n5506 [15]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5523 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3163 (
    .a(\u2_Display/n5487 ),
    .b(\u2_Display/n5506 [16]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5522 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3164 (
    .a(\u2_Display/n5486 ),
    .b(\u2_Display/n5506 [17]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5521 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3165 (
    .a(\u2_Display/n5485 ),
    .b(\u2_Display/n5506 [18]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5520 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3166 (
    .a(\u2_Display/n5484 ),
    .b(\u2_Display/n5506 [19]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5519 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3167 (
    .a(\u2_Display/n5483 ),
    .b(\u2_Display/n5506 [20]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5518 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3168 (
    .a(\u2_Display/n5482 ),
    .b(\u2_Display/n5506 [21]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5517 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3169 (
    .a(\u2_Display/n5481 ),
    .b(\u2_Display/n5506 [22]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5516 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u317 (
    .a(\u1_Driver/n2 [8]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3170 (
    .a(\u2_Display/n5480 ),
    .b(\u2_Display/n5506 [23]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5515 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3171 (
    .a(\u2_Display/n5479 ),
    .b(\u2_Display/n5506 [24]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5514 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3172 (
    .a(\u2_Display/n5478 ),
    .b(\u2_Display/n5506 [25]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5513 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3173 (
    .a(\u2_Display/n5477 ),
    .b(\u2_Display/n5506 [26]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5512 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3174 (
    .a(\u2_Display/n5476 ),
    .b(\u2_Display/n5506 [27]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5511 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3175 (
    .a(\u2_Display/n5475 ),
    .b(\u2_Display/n5506 [28]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5510 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3176 (
    .a(\u2_Display/n5474 ),
    .b(\u2_Display/n5506 [29]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5509 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3177 (
    .a(\u2_Display/n5473 ),
    .b(\u2_Display/n5506 [30]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5508 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3178 (
    .a(\u2_Display/n5472 ),
    .b(\u2_Display/n5506 [31]),
    .c(\u2_Display/n5504 ),
    .o(\u2_Display/n5507 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3179 (
    .a(\u2_Display/n1011 ),
    .b(\u2_Display/n1014 [0]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1046 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u318 (
    .a(\u1_Driver/n2 [7]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3180 (
    .a(\u2_Display/n1010 ),
    .b(\u2_Display/n1014 [1]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1045 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3181 (
    .a(\u2_Display/n1009 ),
    .b(\u2_Display/n1014 [2]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1044 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3182 (
    .a(\u2_Display/n1008 ),
    .b(\u2_Display/n1014 [3]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1043 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3183 (
    .a(\u2_Display/n1007 ),
    .b(\u2_Display/n1014 [4]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1042 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3184 (
    .a(\u2_Display/n1006 ),
    .b(\u2_Display/n1014 [5]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1041 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3185 (
    .a(\u2_Display/n1005 ),
    .b(\u2_Display/n1014 [6]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1040 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3186 (
    .a(\u2_Display/n1004 ),
    .b(\u2_Display/n1014 [7]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1039 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3187 (
    .a(\u2_Display/n1003 ),
    .b(\u2_Display/n1014 [8]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1038 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3188 (
    .a(\u2_Display/n1002 ),
    .b(\u2_Display/n1014 [9]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1037 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3189 (
    .a(\u2_Display/n1001 ),
    .b(\u2_Display/n1014 [10]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1036 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u319 (
    .a(\u1_Driver/n2 [6]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3190 (
    .a(\u2_Display/n1000 ),
    .b(\u2_Display/n1014 [11]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1035 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3191 (
    .a(\u2_Display/n999 ),
    .b(\u2_Display/n1014 [12]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1034 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3192 (
    .a(\u2_Display/n998 ),
    .b(\u2_Display/n1014 [13]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1033 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3193 (
    .a(\u2_Display/n997 ),
    .b(\u2_Display/n1014 [14]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1032 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3194 (
    .a(\u2_Display/n996 ),
    .b(\u2_Display/n1014 [15]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1031 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3195 (
    .a(\u2_Display/n995 ),
    .b(\u2_Display/n1014 [16]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1030 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3196 (
    .a(\u2_Display/n994 ),
    .b(\u2_Display/n1014 [17]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1029 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3197 (
    .a(\u2_Display/n993 ),
    .b(\u2_Display/n1014 [18]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1028 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3198 (
    .a(\u2_Display/n992 ),
    .b(\u2_Display/n1014 [19]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1027 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3199 (
    .a(\u2_Display/n991 ),
    .b(\u2_Display/n1014 [20]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1026 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u320 (
    .a(\u1_Driver/n2 [5]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3200 (
    .a(\u2_Display/n990 ),
    .b(\u2_Display/n1014 [21]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1025 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3201 (
    .a(\u2_Display/n989 ),
    .b(\u2_Display/n1014 [22]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1024 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3202 (
    .a(\u2_Display/n988 ),
    .b(\u2_Display/n1014 [23]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1023 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3203 (
    .a(\u2_Display/n987 ),
    .b(\u2_Display/n1014 [24]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1022 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3204 (
    .a(\u2_Display/n986 ),
    .b(\u2_Display/n1014 [25]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1021 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3205 (
    .a(\u2_Display/n985 ),
    .b(\u2_Display/n1014 [26]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1020 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3206 (
    .a(\u2_Display/n984 ),
    .b(\u2_Display/n1014 [27]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1019 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3207 (
    .a(\u2_Display/n983 ),
    .b(\u2_Display/n1014 [28]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1018 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3208 (
    .a(\u2_Display/n982 ),
    .b(\u2_Display/n1014 [29]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1017 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3209 (
    .a(\u2_Display/n981 ),
    .b(\u2_Display/n1014 [30]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1016 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u321 (
    .a(\u1_Driver/n2 [4]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3210 (
    .a(\u2_Display/n980 ),
    .b(\u2_Display/n1014 [31]),
    .c(\u2_Display/n1012 ),
    .o(\u2_Display/n1015 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3211 (
    .a(\u2_Display/n2134 ),
    .b(\u2_Display/n2137 [0]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2169 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3212 (
    .a(\u2_Display/n2133 ),
    .b(\u2_Display/n2137 [1]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2168 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3213 (
    .a(\u2_Display/n2132 ),
    .b(\u2_Display/n2137 [2]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2167 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3214 (
    .a(\u2_Display/n2131 ),
    .b(\u2_Display/n2137 [3]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2166 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3215 (
    .a(\u2_Display/n2130 ),
    .b(\u2_Display/n2137 [4]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2165 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3216 (
    .a(\u2_Display/n2129 ),
    .b(\u2_Display/n2137 [5]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2164 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3217 (
    .a(\u2_Display/n2128 ),
    .b(\u2_Display/n2137 [6]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2163 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3218 (
    .a(\u2_Display/n2127 ),
    .b(\u2_Display/n2137 [7]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2162 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3219 (
    .a(\u2_Display/n2126 ),
    .b(\u2_Display/n2137 [8]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2161 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u322 (
    .a(\u1_Driver/n2 [3]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3220 (
    .a(\u2_Display/n2125 ),
    .b(\u2_Display/n2137 [9]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2160 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3221 (
    .a(\u2_Display/n2124 ),
    .b(\u2_Display/n2137 [10]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2159 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3222 (
    .a(\u2_Display/n2123 ),
    .b(\u2_Display/n2137 [11]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2158 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3223 (
    .a(\u2_Display/n2122 ),
    .b(\u2_Display/n2137 [12]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2157 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3224 (
    .a(\u2_Display/n2121 ),
    .b(\u2_Display/n2137 [13]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2156 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3225 (
    .a(\u2_Display/n2120 ),
    .b(\u2_Display/n2137 [14]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2155 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3226 (
    .a(\u2_Display/n2119 ),
    .b(\u2_Display/n2137 [15]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2154 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3227 (
    .a(\u2_Display/n2118 ),
    .b(\u2_Display/n2137 [16]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2153 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3228 (
    .a(\u2_Display/n2117 ),
    .b(\u2_Display/n2137 [17]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2152 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3229 (
    .a(\u2_Display/n2116 ),
    .b(\u2_Display/n2137 [18]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2151 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u323 (
    .a(\u1_Driver/n2 [2]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3230 (
    .a(\u2_Display/n2115 ),
    .b(\u2_Display/n2137 [19]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2150 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3231 (
    .a(\u2_Display/n2114 ),
    .b(\u2_Display/n2137 [20]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2149 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3232 (
    .a(\u2_Display/n2113 ),
    .b(\u2_Display/n2137 [21]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2148 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3233 (
    .a(\u2_Display/n2112 ),
    .b(\u2_Display/n2137 [22]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2147 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3234 (
    .a(\u2_Display/n2111 ),
    .b(\u2_Display/n2137 [23]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2146 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3235 (
    .a(\u2_Display/n2110 ),
    .b(\u2_Display/n2137 [24]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2145 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3236 (
    .a(\u2_Display/n2109 ),
    .b(\u2_Display/n2137 [25]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2144 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3237 (
    .a(\u2_Display/n2108 ),
    .b(\u2_Display/n2137 [26]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2143 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3238 (
    .a(\u2_Display/n2107 ),
    .b(\u2_Display/n2137 [27]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2142 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3239 (
    .a(\u2_Display/n2106 ),
    .b(\u2_Display/n2137 [28]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2141 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u324 (
    .a(\u1_Driver/n2 [11]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3240 (
    .a(\u2_Display/n2105 ),
    .b(\u2_Display/n2137 [29]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2140 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3241 (
    .a(\u2_Display/n2104 ),
    .b(\u2_Display/n2137 [30]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2139 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3242 (
    .a(\u2_Display/n2103 ),
    .b(\u2_Display/n2137 [31]),
    .c(\u2_Display/n2135 ),
    .o(\u2_Display/n2138 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3243 (
    .a(\u2_Display/n3257 ),
    .b(\u2_Display/n3260 [0]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3292 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3244 (
    .a(\u2_Display/n3256 ),
    .b(\u2_Display/n3260 [1]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3291 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3245 (
    .a(\u2_Display/n3255 ),
    .b(\u2_Display/n3260 [2]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3290 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3246 (
    .a(\u2_Display/n3254 ),
    .b(\u2_Display/n3260 [3]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3289 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3247 (
    .a(\u2_Display/n3253 ),
    .b(\u2_Display/n3260 [4]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3288 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3248 (
    .a(\u2_Display/n3252 ),
    .b(\u2_Display/n3260 [5]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3287 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3249 (
    .a(\u2_Display/n3251 ),
    .b(\u2_Display/n3260 [6]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3286 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u325 (
    .a(\u1_Driver/n2 [10]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3250 (
    .a(\u2_Display/n3250 ),
    .b(\u2_Display/n3260 [7]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3285 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3251 (
    .a(\u2_Display/n3249 ),
    .b(\u2_Display/n3260 [8]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3284 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3252 (
    .a(\u2_Display/n3248 ),
    .b(\u2_Display/n3260 [9]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3283 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3253 (
    .a(\u2_Display/n3247 ),
    .b(\u2_Display/n3260 [10]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3282 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3254 (
    .a(\u2_Display/n3246 ),
    .b(\u2_Display/n3260 [11]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3281 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3255 (
    .a(\u2_Display/n3245 ),
    .b(\u2_Display/n3260 [12]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3280 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3256 (
    .a(\u2_Display/n3244 ),
    .b(\u2_Display/n3260 [13]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3279 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3257 (
    .a(\u2_Display/n3243 ),
    .b(\u2_Display/n3260 [14]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3278 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3258 (
    .a(\u2_Display/n3242 ),
    .b(\u2_Display/n3260 [15]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3277 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3259 (
    .a(\u2_Display/n3241 ),
    .b(\u2_Display/n3260 [16]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3276 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u326 (
    .a(\u1_Driver/n2 [1]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3260 (
    .a(\u2_Display/n3240 ),
    .b(\u2_Display/n3260 [17]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3275 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3261 (
    .a(\u2_Display/n3239 ),
    .b(\u2_Display/n3260 [18]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3274 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3262 (
    .a(\u2_Display/n3238 ),
    .b(\u2_Display/n3260 [19]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3273 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3263 (
    .a(\u2_Display/n3237 ),
    .b(\u2_Display/n3260 [20]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3272 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3264 (
    .a(\u2_Display/n3236 ),
    .b(\u2_Display/n3260 [21]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3271 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3265 (
    .a(\u2_Display/n3235 ),
    .b(\u2_Display/n3260 [22]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3270 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3266 (
    .a(\u2_Display/n3234 ),
    .b(\u2_Display/n3260 [23]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3269 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3267 (
    .a(\u2_Display/n3233 ),
    .b(\u2_Display/n3260 [24]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3268 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3268 (
    .a(\u2_Display/n3232 ),
    .b(\u2_Display/n3260 [25]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3267 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3269 (
    .a(\u2_Display/n3231 ),
    .b(\u2_Display/n3260 [26]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3266 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u327 (
    .a(\u1_Driver/n2 [0]),
    .b(\u1_Driver/n1 ),
    .o(\u1_Driver/n3 [0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3270 (
    .a(\u2_Display/n3230 ),
    .b(\u2_Display/n3260 [27]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3265 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3271 (
    .a(\u2_Display/n3229 ),
    .b(\u2_Display/n3260 [28]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3264 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3272 (
    .a(\u2_Display/n3228 ),
    .b(\u2_Display/n3260 [29]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3263 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3273 (
    .a(\u2_Display/n3227 ),
    .b(\u2_Display/n3260 [30]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3262 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3274 (
    .a(\u2_Display/n3226 ),
    .b(\u2_Display/n3260 [31]),
    .c(\u2_Display/n3258 ),
    .o(\u2_Display/n3261 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3275 (
    .a(\u2_Display/n4415 ),
    .b(\u2_Display/n4418 [0]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4450 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3276 (
    .a(\u2_Display/n4414 ),
    .b(\u2_Display/n4418 [1]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4449 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3277 (
    .a(\u2_Display/n4413 ),
    .b(\u2_Display/n4418 [2]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4448 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3278 (
    .a(\u2_Display/n4412 ),
    .b(\u2_Display/n4418 [3]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4447 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3279 (
    .a(\u2_Display/n4411 ),
    .b(\u2_Display/n4418 [4]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4446 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u328 (
    .a(\u2_Display/i [10]),
    .b(\u2_Display/i [9]),
    .o(\u2_Display/add7_2_co ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3280 (
    .a(\u2_Display/n4410 ),
    .b(\u2_Display/n4418 [5]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4445 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3281 (
    .a(\u2_Display/n4409 ),
    .b(\u2_Display/n4418 [6]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4444 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3282 (
    .a(\u2_Display/n4408 ),
    .b(\u2_Display/n4418 [7]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4443 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3283 (
    .a(\u2_Display/n4407 ),
    .b(\u2_Display/n4418 [8]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4442 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3284 (
    .a(\u2_Display/n4406 ),
    .b(\u2_Display/n4418 [9]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4441 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3285 (
    .a(\u2_Display/n4405 ),
    .b(\u2_Display/n4418 [10]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4440 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3286 (
    .a(\u2_Display/n4404 ),
    .b(\u2_Display/n4418 [11]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4439 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3287 (
    .a(\u2_Display/n4403 ),
    .b(\u2_Display/n4418 [12]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4438 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3288 (
    .a(\u2_Display/n4402 ),
    .b(\u2_Display/n4418 [13]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4437 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3289 (
    .a(\u2_Display/n4401 ),
    .b(\u2_Display/n4418 [14]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4436 ));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u329 (
    .a(\u2_Display/i [10]),
    .b(\u2_Display/i [9]),
    .o(\u2_Display/n140 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3290 (
    .a(\u2_Display/n4400 ),
    .b(\u2_Display/n4418 [15]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4435 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3291 (
    .a(\u2_Display/n4399 ),
    .b(\u2_Display/n4418 [16]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4434 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3292 (
    .a(\u2_Display/n4398 ),
    .b(\u2_Display/n4418 [17]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4433 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3293 (
    .a(\u2_Display/n4397 ),
    .b(\u2_Display/n4418 [18]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4432 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3294 (
    .a(\u2_Display/n4396 ),
    .b(\u2_Display/n4418 [19]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4431 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3295 (
    .a(\u2_Display/n4395 ),
    .b(\u2_Display/n4418 [20]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4430 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3296 (
    .a(\u2_Display/n4394 ),
    .b(\u2_Display/n4418 [21]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4429 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3297 (
    .a(\u2_Display/n4393 ),
    .b(\u2_Display/n4418 [22]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4428 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3298 (
    .a(\u2_Display/n4392 ),
    .b(\u2_Display/n4418 [23]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4427 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3299 (
    .a(\u2_Display/n4391 ),
    .b(\u2_Display/n4418 [24]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4426 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u330 (
    .a(\u1_Driver/n11 ),
    .b(\u1_Driver/n12 ),
    .c(\u1_Driver/n14 ),
    .d(\u1_Driver/n15 ),
    .o(vga_de_pad));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3300 (
    .a(\u2_Display/n4390 ),
    .b(\u2_Display/n4418 [25]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4425 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3301 (
    .a(\u2_Display/n4389 ),
    .b(\u2_Display/n4418 [26]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4424 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3302 (
    .a(\u2_Display/n4388 ),
    .b(\u2_Display/n4418 [27]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4423 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3303 (
    .a(\u2_Display/n4387 ),
    .b(\u2_Display/n4418 [28]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4422 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3304 (
    .a(\u2_Display/n4386 ),
    .b(\u2_Display/n4418 [29]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4421 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3305 (
    .a(\u2_Display/n4385 ),
    .b(\u2_Display/n4418 [30]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4420 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3306 (
    .a(\u2_Display/n4384 ),
    .b(\u2_Display/n4418 [31]),
    .c(\u2_Display/n4416 ),
    .o(\u2_Display/n4419 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3307 (
    .a(\u2_Display/n5538 ),
    .b(\u2_Display/n5541 [0]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5573 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3308 (
    .a(\u2_Display/n5537 ),
    .b(\u2_Display/n5541 [1]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5572 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3309 (
    .a(\u2_Display/n5536 ),
    .b(\u2_Display/n5541 [2]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5571 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u331 (
    .a(\u2_Display/n3788 [0]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [0]),
    .o(\u2_Display/n3820 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3310 (
    .a(\u2_Display/n5535 ),
    .b(\u2_Display/n5541 [3]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5570 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3311 (
    .a(\u2_Display/n5534 ),
    .b(\u2_Display/n5541 [4]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5569 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3312 (
    .a(\u2_Display/n5533 ),
    .b(\u2_Display/n5541 [5]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5568 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3313 (
    .a(\u2_Display/n5532 ),
    .b(\u2_Display/n5541 [6]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5567 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3314 (
    .a(\u2_Display/n5531 ),
    .b(\u2_Display/n5541 [7]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5566 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3315 (
    .a(\u2_Display/n5530 ),
    .b(\u2_Display/n5541 [8]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5565 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3316 (
    .a(\u2_Display/n5529 ),
    .b(\u2_Display/n5541 [9]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5564 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3317 (
    .a(\u2_Display/n5528 ),
    .b(\u2_Display/n5541 [10]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5563 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3318 (
    .a(\u2_Display/n5527 ),
    .b(\u2_Display/n5541 [11]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5562 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3319 (
    .a(\u2_Display/n5526 ),
    .b(\u2_Display/n5541 [12]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5561 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u332 (
    .a(\u2_Display/n3788 [1]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [1]),
    .o(\u2_Display/n3819 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3320 (
    .a(\u2_Display/n5525 ),
    .b(\u2_Display/n5541 [13]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5560 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3321 (
    .a(\u2_Display/n5524 ),
    .b(\u2_Display/n5541 [14]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5559 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3322 (
    .a(\u2_Display/n5523 ),
    .b(\u2_Display/n5541 [15]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5558 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3323 (
    .a(\u2_Display/n5522 ),
    .b(\u2_Display/n5541 [16]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5557 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3324 (
    .a(\u2_Display/n5521 ),
    .b(\u2_Display/n5541 [17]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5556 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3325 (
    .a(\u2_Display/n5520 ),
    .b(\u2_Display/n5541 [18]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5555 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3326 (
    .a(\u2_Display/n5519 ),
    .b(\u2_Display/n5541 [19]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5554 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3327 (
    .a(\u2_Display/n5518 ),
    .b(\u2_Display/n5541 [20]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5553 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3328 (
    .a(\u2_Display/n5517 ),
    .b(\u2_Display/n5541 [21]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5552 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3329 (
    .a(\u2_Display/n5516 ),
    .b(\u2_Display/n5541 [22]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5551 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u333 (
    .a(\u2_Display/n3788 [2]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [2]),
    .o(\u2_Display/n3818 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3330 (
    .a(\u2_Display/n5515 ),
    .b(\u2_Display/n5541 [23]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5550 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3331 (
    .a(\u2_Display/n5514 ),
    .b(\u2_Display/n5541 [24]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5549 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3332 (
    .a(\u2_Display/n5513 ),
    .b(\u2_Display/n5541 [25]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5548 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3333 (
    .a(\u2_Display/n5512 ),
    .b(\u2_Display/n5541 [26]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5547 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3334 (
    .a(\u2_Display/n5511 ),
    .b(\u2_Display/n5541 [27]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5546 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3335 (
    .a(\u2_Display/n5510 ),
    .b(\u2_Display/n5541 [28]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5545 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3336 (
    .a(\u2_Display/n5509 ),
    .b(\u2_Display/n5541 [29]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5544 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3337 (
    .a(\u2_Display/n5508 ),
    .b(\u2_Display/n5541 [30]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5543 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3338 (
    .a(\u2_Display/n5507 ),
    .b(\u2_Display/n5541 [31]),
    .c(\u2_Display/n5539 ),
    .o(\u2_Display/n5542 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3339 (
    .a(\u2_Display/n1046 ),
    .b(\u2_Display/n1049 [0]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1081 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u334 (
    .a(\u2_Display/n3788 [3]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [3]),
    .o(\u2_Display/n3817 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3340 (
    .a(\u2_Display/n1045 ),
    .b(\u2_Display/n1049 [1]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1080 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3341 (
    .a(\u2_Display/n1044 ),
    .b(\u2_Display/n1049 [2]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1079 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3342 (
    .a(\u2_Display/n1043 ),
    .b(\u2_Display/n1049 [3]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1078 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3343 (
    .a(\u2_Display/n1042 ),
    .b(\u2_Display/n1049 [4]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1077 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3344 (
    .a(\u2_Display/n1041 ),
    .b(\u2_Display/n1049 [5]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1076 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3345 (
    .a(\u2_Display/n1040 ),
    .b(\u2_Display/n1049 [6]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1075 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3346 (
    .a(\u2_Display/n1039 ),
    .b(\u2_Display/n1049 [7]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1074 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3347 (
    .a(\u2_Display/n1038 ),
    .b(\u2_Display/n1049 [8]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1073 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3348 (
    .a(\u2_Display/n1037 ),
    .b(\u2_Display/n1049 [9]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1072 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3349 (
    .a(\u2_Display/n1036 ),
    .b(\u2_Display/n1049 [10]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1071 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u335 (
    .a(\u2_Display/n3788 [4]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [4]),
    .o(\u2_Display/n3816 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3350 (
    .a(\u2_Display/n1035 ),
    .b(\u2_Display/n1049 [11]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1070 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3351 (
    .a(\u2_Display/n1034 ),
    .b(\u2_Display/n1049 [12]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1069 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3352 (
    .a(\u2_Display/n1033 ),
    .b(\u2_Display/n1049 [13]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1068 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3353 (
    .a(\u2_Display/n1032 ),
    .b(\u2_Display/n1049 [14]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1067 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3354 (
    .a(\u2_Display/n1031 ),
    .b(\u2_Display/n1049 [15]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1066 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3355 (
    .a(\u2_Display/n1030 ),
    .b(\u2_Display/n1049 [16]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1065 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3356 (
    .a(\u2_Display/n1029 ),
    .b(\u2_Display/n1049 [17]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1064 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3357 (
    .a(\u2_Display/n1028 ),
    .b(\u2_Display/n1049 [18]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1063 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3358 (
    .a(\u2_Display/n1027 ),
    .b(\u2_Display/n1049 [19]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1062 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3359 (
    .a(\u2_Display/n1026 ),
    .b(\u2_Display/n1049 [20]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1061 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u336 (
    .a(\u2_Display/n3788 [5]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [5]),
    .o(\u2_Display/n3815 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3360 (
    .a(\u2_Display/n1025 ),
    .b(\u2_Display/n1049 [21]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1060 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3361 (
    .a(\u2_Display/n1024 ),
    .b(\u2_Display/n1049 [22]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1059 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3362 (
    .a(\u2_Display/n1023 ),
    .b(\u2_Display/n1049 [23]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1058 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3363 (
    .a(\u2_Display/n1022 ),
    .b(\u2_Display/n1049 [24]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1057 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3364 (
    .a(\u2_Display/n1021 ),
    .b(\u2_Display/n1049 [25]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1056 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3365 (
    .a(\u2_Display/n1020 ),
    .b(\u2_Display/n1049 [26]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1055 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3366 (
    .a(\u2_Display/n1019 ),
    .b(\u2_Display/n1049 [27]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1054 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3367 (
    .a(\u2_Display/n1018 ),
    .b(\u2_Display/n1049 [28]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1053 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3368 (
    .a(\u2_Display/n1017 ),
    .b(\u2_Display/n1049 [29]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1052 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3369 (
    .a(\u2_Display/n1016 ),
    .b(\u2_Display/n1049 [30]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1051 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u337 (
    .a(\u2_Display/n3788 [6]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [6]),
    .o(\u2_Display/n3814 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3370 (
    .a(\u2_Display/n1015 ),
    .b(\u2_Display/n1049 [31]),
    .c(\u2_Display/n1047 ),
    .o(\u2_Display/n1050 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3371 (
    .a(\u2_Display/n2169 ),
    .b(\u2_Display/n2172 [0]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2204 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3372 (
    .a(\u2_Display/n2168 ),
    .b(\u2_Display/n2172 [1]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2203 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3373 (
    .a(\u2_Display/n2167 ),
    .b(\u2_Display/n2172 [2]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2202 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3374 (
    .a(\u2_Display/n2166 ),
    .b(\u2_Display/n2172 [3]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2201 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3375 (
    .a(\u2_Display/n2165 ),
    .b(\u2_Display/n2172 [4]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2200 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3376 (
    .a(\u2_Display/n2164 ),
    .b(\u2_Display/n2172 [5]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2199 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3377 (
    .a(\u2_Display/n2163 ),
    .b(\u2_Display/n2172 [6]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2198 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3378 (
    .a(\u2_Display/n2162 ),
    .b(\u2_Display/n2172 [7]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2197 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3379 (
    .a(\u2_Display/n2161 ),
    .b(\u2_Display/n2172 [8]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2196 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u338 (
    .a(\u2_Display/n3788 [7]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [7]),
    .o(\u2_Display/n3813 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3380 (
    .a(\u2_Display/n2160 ),
    .b(\u2_Display/n2172 [9]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2195 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3381 (
    .a(\u2_Display/n2159 ),
    .b(\u2_Display/n2172 [10]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2194 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3382 (
    .a(\u2_Display/n2158 ),
    .b(\u2_Display/n2172 [11]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2193 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3383 (
    .a(\u2_Display/n2157 ),
    .b(\u2_Display/n2172 [12]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2192 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3384 (
    .a(\u2_Display/n2156 ),
    .b(\u2_Display/n2172 [13]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2191 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3385 (
    .a(\u2_Display/n2155 ),
    .b(\u2_Display/n2172 [14]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2190 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3386 (
    .a(\u2_Display/n2154 ),
    .b(\u2_Display/n2172 [15]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2189 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3387 (
    .a(\u2_Display/n2153 ),
    .b(\u2_Display/n2172 [16]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2188 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3388 (
    .a(\u2_Display/n2152 ),
    .b(\u2_Display/n2172 [17]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2187 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3389 (
    .a(\u2_Display/n2151 ),
    .b(\u2_Display/n2172 [18]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2186 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u339 (
    .a(\u2_Display/n3788 [8]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [8]),
    .o(\u2_Display/n3812 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3390 (
    .a(\u2_Display/n2150 ),
    .b(\u2_Display/n2172 [19]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2185 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3391 (
    .a(\u2_Display/n2149 ),
    .b(\u2_Display/n2172 [20]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2184 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3392 (
    .a(\u2_Display/n2148 ),
    .b(\u2_Display/n2172 [21]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2183 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3393 (
    .a(\u2_Display/n2147 ),
    .b(\u2_Display/n2172 [22]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2182 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3394 (
    .a(\u2_Display/n2146 ),
    .b(\u2_Display/n2172 [23]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2181 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3395 (
    .a(\u2_Display/n2145 ),
    .b(\u2_Display/n2172 [24]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2180 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3396 (
    .a(\u2_Display/n2144 ),
    .b(\u2_Display/n2172 [25]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2179 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3397 (
    .a(\u2_Display/n2143 ),
    .b(\u2_Display/n2172 [26]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2178 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3398 (
    .a(\u2_Display/n2142 ),
    .b(\u2_Display/n2172 [27]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2177 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3399 (
    .a(\u2_Display/n2141 ),
    .b(\u2_Display/n2172 [28]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2176 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u340 (
    .a(\u2_Display/n3788 [9]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [9]),
    .o(\u2_Display/n3811 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3400 (
    .a(\u2_Display/n2140 ),
    .b(\u2_Display/n2172 [29]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2175 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3401 (
    .a(\u2_Display/n2139 ),
    .b(\u2_Display/n2172 [30]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2174 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3402 (
    .a(\u2_Display/n2138 ),
    .b(\u2_Display/n2172 [31]),
    .c(\u2_Display/n2170 ),
    .o(\u2_Display/n2173 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3403 (
    .a(\u2_Display/n3292 ),
    .b(\u2_Display/n3295 [0]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3327 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3404 (
    .a(\u2_Display/n3291 ),
    .b(\u2_Display/n3295 [1]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3326 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3405 (
    .a(\u2_Display/n3290 ),
    .b(\u2_Display/n3295 [2]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3325 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3406 (
    .a(\u2_Display/n3289 ),
    .b(\u2_Display/n3295 [3]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3324 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3407 (
    .a(\u2_Display/n3288 ),
    .b(\u2_Display/n3295 [4]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3323 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3408 (
    .a(\u2_Display/n3287 ),
    .b(\u2_Display/n3295 [5]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3322 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3409 (
    .a(\u2_Display/n3286 ),
    .b(\u2_Display/n3295 [6]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3321 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u341 (
    .a(\u2_Display/n3788 [10]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [10]),
    .o(\u2_Display/n3810 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3410 (
    .a(\u2_Display/n3285 ),
    .b(\u2_Display/n3295 [7]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3320 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3411 (
    .a(\u2_Display/n3284 ),
    .b(\u2_Display/n3295 [8]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3319 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3412 (
    .a(\u2_Display/n3283 ),
    .b(\u2_Display/n3295 [9]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3318 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3413 (
    .a(\u2_Display/n3282 ),
    .b(\u2_Display/n3295 [10]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3317 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3414 (
    .a(\u2_Display/n3281 ),
    .b(\u2_Display/n3295 [11]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3316 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3415 (
    .a(\u2_Display/n3280 ),
    .b(\u2_Display/n3295 [12]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3315 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3416 (
    .a(\u2_Display/n3279 ),
    .b(\u2_Display/n3295 [13]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3314 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3417 (
    .a(\u2_Display/n3278 ),
    .b(\u2_Display/n3295 [14]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3313 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3418 (
    .a(\u2_Display/n3277 ),
    .b(\u2_Display/n3295 [15]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3312 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3419 (
    .a(\u2_Display/n3276 ),
    .b(\u2_Display/n3295 [16]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3311 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u342 (
    .a(\u2_Display/n3788 [11]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [11]),
    .o(\u2_Display/n3809 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3420 (
    .a(\u2_Display/n3275 ),
    .b(\u2_Display/n3295 [17]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3310 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3421 (
    .a(\u2_Display/n3274 ),
    .b(\u2_Display/n3295 [18]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3309 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3422 (
    .a(\u2_Display/n3273 ),
    .b(\u2_Display/n3295 [19]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3308 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3423 (
    .a(\u2_Display/n3272 ),
    .b(\u2_Display/n3295 [20]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3307 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3424 (
    .a(\u2_Display/n3271 ),
    .b(\u2_Display/n3295 [21]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3306 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3425 (
    .a(\u2_Display/n3270 ),
    .b(\u2_Display/n3295 [22]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3305 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3426 (
    .a(\u2_Display/n3269 ),
    .b(\u2_Display/n3295 [23]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3304 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3427 (
    .a(\u2_Display/n3268 ),
    .b(\u2_Display/n3295 [24]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3303 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3428 (
    .a(\u2_Display/n3267 ),
    .b(\u2_Display/n3295 [25]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3302 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3429 (
    .a(\u2_Display/n3266 ),
    .b(\u2_Display/n3295 [26]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3301 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u343 (
    .a(\u2_Display/n3788 [12]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [12]),
    .o(\u2_Display/n3808 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3430 (
    .a(\u2_Display/n3265 ),
    .b(\u2_Display/n3295 [27]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3300 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3431 (
    .a(\u2_Display/n3264 ),
    .b(\u2_Display/n3295 [28]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3299 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3432 (
    .a(\u2_Display/n3263 ),
    .b(\u2_Display/n3295 [29]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3298 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3433 (
    .a(\u2_Display/n3262 ),
    .b(\u2_Display/n3295 [30]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3297 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3434 (
    .a(\u2_Display/n3261 ),
    .b(\u2_Display/n3295 [31]),
    .c(\u2_Display/n3293 ),
    .o(\u2_Display/n3296 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3435 (
    .a(\u2_Display/n4450 ),
    .b(\u2_Display/n4453 [0]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4485 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3436 (
    .a(\u2_Display/n4449 ),
    .b(\u2_Display/n4453 [1]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4484 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3437 (
    .a(\u2_Display/n4448 ),
    .b(\u2_Display/n4453 [2]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4483 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3438 (
    .a(\u2_Display/n4447 ),
    .b(\u2_Display/n4453 [3]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4482 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3439 (
    .a(\u2_Display/n4446 ),
    .b(\u2_Display/n4453 [4]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4481 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u344 (
    .a(\u2_Display/n3788 [13]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [13]),
    .o(\u2_Display/n3807 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3440 (
    .a(\u2_Display/n4445 ),
    .b(\u2_Display/n4453 [5]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4480 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3441 (
    .a(\u2_Display/n4444 ),
    .b(\u2_Display/n4453 [6]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4479 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3442 (
    .a(\u2_Display/n4443 ),
    .b(\u2_Display/n4453 [7]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4478 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3443 (
    .a(\u2_Display/n4442 ),
    .b(\u2_Display/n4453 [8]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4477 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3444 (
    .a(\u2_Display/n4441 ),
    .b(\u2_Display/n4453 [9]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4476 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3445 (
    .a(\u2_Display/n4440 ),
    .b(\u2_Display/n4453 [10]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4475 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3446 (
    .a(\u2_Display/n4439 ),
    .b(\u2_Display/n4453 [11]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4474 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3447 (
    .a(\u2_Display/n4438 ),
    .b(\u2_Display/n4453 [12]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4473 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3448 (
    .a(\u2_Display/n4437 ),
    .b(\u2_Display/n4453 [13]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4472 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3449 (
    .a(\u2_Display/n4436 ),
    .b(\u2_Display/n4453 [14]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4471 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u345 (
    .a(\u2_Display/n3788 [14]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [14]),
    .o(\u2_Display/n3806 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3450 (
    .a(\u2_Display/n4435 ),
    .b(\u2_Display/n4453 [15]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4470 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3451 (
    .a(\u2_Display/n4434 ),
    .b(\u2_Display/n4453 [16]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4469 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3452 (
    .a(\u2_Display/n4433 ),
    .b(\u2_Display/n4453 [17]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4468 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3453 (
    .a(\u2_Display/n4432 ),
    .b(\u2_Display/n4453 [18]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4467 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3454 (
    .a(\u2_Display/n4431 ),
    .b(\u2_Display/n4453 [19]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4466 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3455 (
    .a(\u2_Display/n4430 ),
    .b(\u2_Display/n4453 [20]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4465 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3456 (
    .a(\u2_Display/n4429 ),
    .b(\u2_Display/n4453 [21]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4464 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3457 (
    .a(\u2_Display/n4428 ),
    .b(\u2_Display/n4453 [22]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4463 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3458 (
    .a(\u2_Display/n4427 ),
    .b(\u2_Display/n4453 [23]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4462 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3459 (
    .a(\u2_Display/n4426 ),
    .b(\u2_Display/n4453 [24]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4461 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u346 (
    .a(\u2_Display/n3788 [15]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [15]),
    .o(\u2_Display/n3805 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3460 (
    .a(\u2_Display/n4425 ),
    .b(\u2_Display/n4453 [25]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4460 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3461 (
    .a(\u2_Display/n4424 ),
    .b(\u2_Display/n4453 [26]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4459 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3462 (
    .a(\u2_Display/n4423 ),
    .b(\u2_Display/n4453 [27]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4458 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3463 (
    .a(\u2_Display/n4422 ),
    .b(\u2_Display/n4453 [28]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4457 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3464 (
    .a(\u2_Display/n4421 ),
    .b(\u2_Display/n4453 [29]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4456 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3465 (
    .a(\u2_Display/n4420 ),
    .b(\u2_Display/n4453 [30]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4455 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3466 (
    .a(\u2_Display/n4419 ),
    .b(\u2_Display/n4453 [31]),
    .c(\u2_Display/n4451 ),
    .o(\u2_Display/n4454 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3467 (
    .a(\u2_Display/n5573 ),
    .b(\u2_Display/n5576 [0]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5608 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3468 (
    .a(\u2_Display/n5572 ),
    .b(\u2_Display/n5576 [1]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5607 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3469 (
    .a(\u2_Display/n5571 ),
    .b(\u2_Display/n5576 [2]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5606 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u347 (
    .a(\u2_Display/n3788 [16]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [16]),
    .o(\u2_Display/n3804 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3470 (
    .a(\u2_Display/n5570 ),
    .b(\u2_Display/n5576 [3]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5605 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3471 (
    .a(\u2_Display/n5569 ),
    .b(\u2_Display/n5576 [4]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5604 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3472 (
    .a(\u2_Display/n5568 ),
    .b(\u2_Display/n5576 [5]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5603 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3473 (
    .a(\u2_Display/n5567 ),
    .b(\u2_Display/n5576 [6]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5602 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3474 (
    .a(\u2_Display/n5566 ),
    .b(\u2_Display/n5576 [7]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5601 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3475 (
    .a(\u2_Display/n5565 ),
    .b(\u2_Display/n5576 [8]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5600 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3476 (
    .a(\u2_Display/n5564 ),
    .b(\u2_Display/n5576 [9]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5599 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3477 (
    .a(\u2_Display/n5563 ),
    .b(\u2_Display/n5576 [10]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5598 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3478 (
    .a(\u2_Display/n5562 ),
    .b(\u2_Display/n5576 [11]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5597 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3479 (
    .a(\u2_Display/n5561 ),
    .b(\u2_Display/n5576 [12]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5596 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u348 (
    .a(\u2_Display/n3788 [17]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [17]),
    .o(\u2_Display/n3803 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3480 (
    .a(\u2_Display/n5560 ),
    .b(\u2_Display/n5576 [13]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5595 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3481 (
    .a(\u2_Display/n5559 ),
    .b(\u2_Display/n5576 [14]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5594 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3482 (
    .a(\u2_Display/n5558 ),
    .b(\u2_Display/n5576 [15]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5593 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3483 (
    .a(\u2_Display/n5557 ),
    .b(\u2_Display/n5576 [16]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5592 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3484 (
    .a(\u2_Display/n5556 ),
    .b(\u2_Display/n5576 [17]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5591 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3485 (
    .a(\u2_Display/n5555 ),
    .b(\u2_Display/n5576 [18]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5590 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3486 (
    .a(\u2_Display/n5554 ),
    .b(\u2_Display/n5576 [19]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5589 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3487 (
    .a(\u2_Display/n5553 ),
    .b(\u2_Display/n5576 [20]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5588 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3488 (
    .a(\u2_Display/n5552 ),
    .b(\u2_Display/n5576 [21]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5587 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3489 (
    .a(\u2_Display/n5551 ),
    .b(\u2_Display/n5576 [22]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5586 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u349 (
    .a(\u2_Display/n3788 [18]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [18]),
    .o(\u2_Display/n3802 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3490 (
    .a(\u2_Display/n5550 ),
    .b(\u2_Display/n5576 [23]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5585 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3491 (
    .a(\u2_Display/n5549 ),
    .b(\u2_Display/n5576 [24]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5584 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3492 (
    .a(\u2_Display/n5548 ),
    .b(\u2_Display/n5576 [25]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5583 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3493 (
    .a(\u2_Display/n5547 ),
    .b(\u2_Display/n5576 [26]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5582 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3494 (
    .a(\u2_Display/n5546 ),
    .b(\u2_Display/n5576 [27]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5581 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3495 (
    .a(\u2_Display/n5545 ),
    .b(\u2_Display/n5576 [28]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5580 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3496 (
    .a(\u2_Display/n5544 ),
    .b(\u2_Display/n5576 [29]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5579 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3497 (
    .a(\u2_Display/n5543 ),
    .b(\u2_Display/n5576 [30]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5578 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3498 (
    .a(\u2_Display/n5542 ),
    .b(\u2_Display/n5576 [31]),
    .c(\u2_Display/n5574 ),
    .o(\u2_Display/n5577 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3499 (
    .a(\u2_Display/n1081 ),
    .b(\u2_Display/n1084 [0]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1116 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u350 (
    .a(\u2_Display/n3788 [19]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [19]),
    .o(\u2_Display/n3801 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3500 (
    .a(\u2_Display/n1080 ),
    .b(\u2_Display/n1084 [1]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1115 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3501 (
    .a(\u2_Display/n1079 ),
    .b(\u2_Display/n1084 [2]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1114 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3502 (
    .a(\u2_Display/n1078 ),
    .b(\u2_Display/n1084 [3]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1113 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3503 (
    .a(\u2_Display/n1077 ),
    .b(\u2_Display/n1084 [4]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1112 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3504 (
    .a(\u2_Display/n1076 ),
    .b(\u2_Display/n1084 [5]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1111 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3505 (
    .a(\u2_Display/n1075 ),
    .b(\u2_Display/n1084 [6]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1110 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3506 (
    .a(\u2_Display/n1074 ),
    .b(\u2_Display/n1084 [7]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1109 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3507 (
    .a(\u2_Display/n1073 ),
    .b(\u2_Display/n1084 [8]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1108 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3508 (
    .a(\u2_Display/n1072 ),
    .b(\u2_Display/n1084 [9]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1107 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3509 (
    .a(\u2_Display/n1071 ),
    .b(\u2_Display/n1084 [10]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1106 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u351 (
    .a(\u2_Display/n3788 [20]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [20]),
    .o(\u2_Display/n3800 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3510 (
    .a(\u2_Display/n1070 ),
    .b(\u2_Display/n1084 [11]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1105 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3511 (
    .a(\u2_Display/n1069 ),
    .b(\u2_Display/n1084 [12]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1104 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3512 (
    .a(\u2_Display/n1068 ),
    .b(\u2_Display/n1084 [13]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1103 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3513 (
    .a(\u2_Display/n1067 ),
    .b(\u2_Display/n1084 [14]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1102 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3514 (
    .a(\u2_Display/n1066 ),
    .b(\u2_Display/n1084 [15]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1101 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3515 (
    .a(\u2_Display/n1065 ),
    .b(\u2_Display/n1084 [16]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1100 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3516 (
    .a(\u2_Display/n1064 ),
    .b(\u2_Display/n1084 [17]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1099 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3517 (
    .a(\u2_Display/n1063 ),
    .b(\u2_Display/n1084 [18]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1098 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3518 (
    .a(\u2_Display/n1062 ),
    .b(\u2_Display/n1084 [19]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1097 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3519 (
    .a(\u2_Display/n1061 ),
    .b(\u2_Display/n1084 [20]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1096 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u352 (
    .a(\u2_Display/n3788 [21]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [21]),
    .o(\u2_Display/n3799 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3520 (
    .a(\u2_Display/n1060 ),
    .b(\u2_Display/n1084 [21]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1095 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3521 (
    .a(\u2_Display/n1059 ),
    .b(\u2_Display/n1084 [22]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1094 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3522 (
    .a(\u2_Display/n1058 ),
    .b(\u2_Display/n1084 [23]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1093 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3523 (
    .a(\u2_Display/n1057 ),
    .b(\u2_Display/n1084 [24]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1092 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3524 (
    .a(\u2_Display/n1056 ),
    .b(\u2_Display/n1084 [25]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1091 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3525 (
    .a(\u2_Display/n1055 ),
    .b(\u2_Display/n1084 [26]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1090 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3526 (
    .a(\u2_Display/n1054 ),
    .b(\u2_Display/n1084 [27]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1089 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3527 (
    .a(\u2_Display/n1053 ),
    .b(\u2_Display/n1084 [28]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1088 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3528 (
    .a(\u2_Display/n1052 ),
    .b(\u2_Display/n1084 [29]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1087 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3529 (
    .a(\u2_Display/n1051 ),
    .b(\u2_Display/n1084 [30]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1086 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u353 (
    .a(\u2_Display/n3788 [22]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [22]),
    .o(\u2_Display/n3798 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3530 (
    .a(\u2_Display/n1050 ),
    .b(\u2_Display/n1084 [31]),
    .c(\u2_Display/n1082 ),
    .o(\u2_Display/n1085 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3531 (
    .a(\u2_Display/n2204 ),
    .b(\u2_Display/n2207 [0]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2239 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3532 (
    .a(\u2_Display/n2203 ),
    .b(\u2_Display/n2207 [1]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2238 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3533 (
    .a(\u2_Display/n2202 ),
    .b(\u2_Display/n2207 [2]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2237 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3534 (
    .a(\u2_Display/n2201 ),
    .b(\u2_Display/n2207 [3]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2236 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3535 (
    .a(\u2_Display/n2200 ),
    .b(\u2_Display/n2207 [4]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2235 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3536 (
    .a(\u2_Display/n2199 ),
    .b(\u2_Display/n2207 [5]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2234 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3537 (
    .a(\u2_Display/n2198 ),
    .b(\u2_Display/n2207 [6]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2233 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3538 (
    .a(\u2_Display/n2197 ),
    .b(\u2_Display/n2207 [7]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2232 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3539 (
    .a(\u2_Display/n2196 ),
    .b(\u2_Display/n2207 [8]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2231 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u354 (
    .a(\u2_Display/n3788 [23]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [23]),
    .o(\u2_Display/n3797 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3540 (
    .a(\u2_Display/n2195 ),
    .b(\u2_Display/n2207 [9]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2230 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3541 (
    .a(\u2_Display/n2194 ),
    .b(\u2_Display/n2207 [10]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2229 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3542 (
    .a(\u2_Display/n2193 ),
    .b(\u2_Display/n2207 [11]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2228 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3543 (
    .a(\u2_Display/n2192 ),
    .b(\u2_Display/n2207 [12]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2227 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3544 (
    .a(\u2_Display/n2191 ),
    .b(\u2_Display/n2207 [13]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2226 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3545 (
    .a(\u2_Display/n2190 ),
    .b(\u2_Display/n2207 [14]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2225 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3546 (
    .a(\u2_Display/n2189 ),
    .b(\u2_Display/n2207 [15]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2224 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3547 (
    .a(\u2_Display/n2188 ),
    .b(\u2_Display/n2207 [16]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2223 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3548 (
    .a(\u2_Display/n2187 ),
    .b(\u2_Display/n2207 [17]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2222 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3549 (
    .a(\u2_Display/n2186 ),
    .b(\u2_Display/n2207 [18]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2221 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u355 (
    .a(\u2_Display/n3788 [24]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [24]),
    .o(\u2_Display/n3796 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3550 (
    .a(\u2_Display/n2185 ),
    .b(\u2_Display/n2207 [19]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2220 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3551 (
    .a(\u2_Display/n2184 ),
    .b(\u2_Display/n2207 [20]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2219 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3552 (
    .a(\u2_Display/n2183 ),
    .b(\u2_Display/n2207 [21]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2218 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3553 (
    .a(\u2_Display/n2182 ),
    .b(\u2_Display/n2207 [22]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2217 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3554 (
    .a(\u2_Display/n2181 ),
    .b(\u2_Display/n2207 [23]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2216 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3555 (
    .a(\u2_Display/n2180 ),
    .b(\u2_Display/n2207 [24]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2215 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3556 (
    .a(\u2_Display/n2179 ),
    .b(\u2_Display/n2207 [25]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2214 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3557 (
    .a(\u2_Display/n2178 ),
    .b(\u2_Display/n2207 [26]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2213 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3558 (
    .a(\u2_Display/n2177 ),
    .b(\u2_Display/n2207 [27]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2212 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3559 (
    .a(\u2_Display/n2176 ),
    .b(\u2_Display/n2207 [28]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2211 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u356 (
    .a(\u2_Display/n3788 [25]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [25]),
    .o(\u2_Display/n3795 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3560 (
    .a(\u2_Display/n2175 ),
    .b(\u2_Display/n2207 [29]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2210 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3561 (
    .a(\u2_Display/n2174 ),
    .b(\u2_Display/n2207 [30]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2209 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3562 (
    .a(\u2_Display/n2173 ),
    .b(\u2_Display/n2207 [31]),
    .c(\u2_Display/n2205 ),
    .o(\u2_Display/n2208 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3563 (
    .a(\u2_Display/n3327 ),
    .b(\u2_Display/n3330 [0]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3362 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3564 (
    .a(\u2_Display/n3326 ),
    .b(\u2_Display/n3330 [1]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3361 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3565 (
    .a(\u2_Display/n3325 ),
    .b(\u2_Display/n3330 [2]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3360 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3566 (
    .a(\u2_Display/n3324 ),
    .b(\u2_Display/n3330 [3]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3359 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3567 (
    .a(\u2_Display/n3323 ),
    .b(\u2_Display/n3330 [4]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3358 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3568 (
    .a(\u2_Display/n3322 ),
    .b(\u2_Display/n3330 [5]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3357 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3569 (
    .a(\u2_Display/n3321 ),
    .b(\u2_Display/n3330 [6]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3356 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u357 (
    .a(\u2_Display/n3788 [26]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [26]),
    .o(\u2_Display/n3794 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3570 (
    .a(\u2_Display/n3320 ),
    .b(\u2_Display/n3330 [7]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3355 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3571 (
    .a(\u2_Display/n3319 ),
    .b(\u2_Display/n3330 [8]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3354 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3572 (
    .a(\u2_Display/n3318 ),
    .b(\u2_Display/n3330 [9]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3353 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3573 (
    .a(\u2_Display/n3317 ),
    .b(\u2_Display/n3330 [10]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3352 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3574 (
    .a(\u2_Display/n3316 ),
    .b(\u2_Display/n3330 [11]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3351 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3575 (
    .a(\u2_Display/n3315 ),
    .b(\u2_Display/n3330 [12]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3350 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3576 (
    .a(\u2_Display/n3314 ),
    .b(\u2_Display/n3330 [13]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3349 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3577 (
    .a(\u2_Display/n3313 ),
    .b(\u2_Display/n3330 [14]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3348 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3578 (
    .a(\u2_Display/n3312 ),
    .b(\u2_Display/n3330 [15]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3347 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3579 (
    .a(\u2_Display/n3311 ),
    .b(\u2_Display/n3330 [16]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3346 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u358 (
    .a(\u2_Display/n3788 [27]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [27]),
    .o(\u2_Display/n3793 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3580 (
    .a(\u2_Display/n3310 ),
    .b(\u2_Display/n3330 [17]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3345 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3581 (
    .a(\u2_Display/n3309 ),
    .b(\u2_Display/n3330 [18]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3344 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3582 (
    .a(\u2_Display/n3308 ),
    .b(\u2_Display/n3330 [19]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3343 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3583 (
    .a(\u2_Display/n3307 ),
    .b(\u2_Display/n3330 [20]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3342 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3584 (
    .a(\u2_Display/n3306 ),
    .b(\u2_Display/n3330 [21]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3341 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3585 (
    .a(\u2_Display/n3305 ),
    .b(\u2_Display/n3330 [22]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3340 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3586 (
    .a(\u2_Display/n3304 ),
    .b(\u2_Display/n3330 [23]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3339 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3587 (
    .a(\u2_Display/n3303 ),
    .b(\u2_Display/n3330 [24]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3338 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3588 (
    .a(\u2_Display/n3302 ),
    .b(\u2_Display/n3330 [25]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3337 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3589 (
    .a(\u2_Display/n3301 ),
    .b(\u2_Display/n3330 [26]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3336 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u359 (
    .a(\u2_Display/n3788 [28]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [28]),
    .o(\u2_Display/n3792 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3590 (
    .a(\u2_Display/n3300 ),
    .b(\u2_Display/n3330 [27]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3335 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3591 (
    .a(\u2_Display/n3299 ),
    .b(\u2_Display/n3330 [28]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3334 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3592 (
    .a(\u2_Display/n3298 ),
    .b(\u2_Display/n3330 [29]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3333 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3593 (
    .a(\u2_Display/n3297 ),
    .b(\u2_Display/n3330 [30]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3332 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3594 (
    .a(\u2_Display/n3296 ),
    .b(\u2_Display/n3330 [31]),
    .c(\u2_Display/n3328 ),
    .o(\u2_Display/n3331 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3595 (
    .a(\u2_Display/n4485 ),
    .b(\u2_Display/n4488 [0]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4520 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3596 (
    .a(\u2_Display/n4484 ),
    .b(\u2_Display/n4488 [1]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4519 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3597 (
    .a(\u2_Display/n4483 ),
    .b(\u2_Display/n4488 [2]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4518 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3598 (
    .a(\u2_Display/n4482 ),
    .b(\u2_Display/n4488 [3]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4517 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3599 (
    .a(\u2_Display/n4481 ),
    .b(\u2_Display/n4488 [4]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4516 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u360 (
    .a(\u2_Display/n3788 [29]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [29]),
    .o(\u2_Display/n3791 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3600 (
    .a(\u2_Display/n4480 ),
    .b(\u2_Display/n4488 [5]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4515 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3601 (
    .a(\u2_Display/n4479 ),
    .b(\u2_Display/n4488 [6]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4514 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3602 (
    .a(\u2_Display/n4478 ),
    .b(\u2_Display/n4488 [7]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4513 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3603 (
    .a(\u2_Display/n4477 ),
    .b(\u2_Display/n4488 [8]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4512 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3604 (
    .a(\u2_Display/n4476 ),
    .b(\u2_Display/n4488 [9]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4511 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3605 (
    .a(\u2_Display/n4475 ),
    .b(\u2_Display/n4488 [10]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4510 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3606 (
    .a(\u2_Display/n4474 ),
    .b(\u2_Display/n4488 [11]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4509 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3607 (
    .a(\u2_Display/n4473 ),
    .b(\u2_Display/n4488 [12]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4508 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3608 (
    .a(\u2_Display/n4472 ),
    .b(\u2_Display/n4488 [13]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4507 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3609 (
    .a(\u2_Display/n4471 ),
    .b(\u2_Display/n4488 [14]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4506 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u361 (
    .a(\u2_Display/n3788 [30]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [30]),
    .o(\u2_Display/n3790 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3610 (
    .a(\u2_Display/n4470 ),
    .b(\u2_Display/n4488 [15]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4505 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3611 (
    .a(\u2_Display/n4469 ),
    .b(\u2_Display/n4488 [16]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4504 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3612 (
    .a(\u2_Display/n4468 ),
    .b(\u2_Display/n4488 [17]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4503 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3613 (
    .a(\u2_Display/n4467 ),
    .b(\u2_Display/n4488 [18]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4502 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3614 (
    .a(\u2_Display/n4466 ),
    .b(\u2_Display/n4488 [19]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4501 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3615 (
    .a(\u2_Display/n4465 ),
    .b(\u2_Display/n4488 [20]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4500 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3616 (
    .a(\u2_Display/n4464 ),
    .b(\u2_Display/n4488 [21]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4499 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3617 (
    .a(\u2_Display/n4463 ),
    .b(\u2_Display/n4488 [22]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4498 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3618 (
    .a(\u2_Display/n4462 ),
    .b(\u2_Display/n4488 [23]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4497 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3619 (
    .a(\u2_Display/n4461 ),
    .b(\u2_Display/n4488 [24]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4496 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u362 (
    .a(\u2_Display/n3788 [31]),
    .b(\u2_Display/n3786 ),
    .c(\u2_Display/counta [31]),
    .o(\u2_Display/n3789 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3620 (
    .a(\u2_Display/n4460 ),
    .b(\u2_Display/n4488 [25]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4495 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3621 (
    .a(\u2_Display/n4459 ),
    .b(\u2_Display/n4488 [26]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4494 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3622 (
    .a(\u2_Display/n4458 ),
    .b(\u2_Display/n4488 [27]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4493 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3623 (
    .a(\u2_Display/n4457 ),
    .b(\u2_Display/n4488 [28]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4492 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3624 (
    .a(\u2_Display/n4456 ),
    .b(\u2_Display/n4488 [29]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4491 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3625 (
    .a(\u2_Display/n4455 ),
    .b(\u2_Display/n4488 [30]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4490 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3626 (
    .a(\u2_Display/n4454 ),
    .b(\u2_Display/n4488 [31]),
    .c(\u2_Display/n4486 ),
    .o(\u2_Display/n4489 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3627 (
    .a(\u2_Display/n5608 ),
    .b(\u2_Display/n5611 [0]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5643 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3628 (
    .a(\u2_Display/n5607 ),
    .b(\u2_Display/n5611 [1]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5642 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3629 (
    .a(\u2_Display/n5606 ),
    .b(\u2_Display/n5611 [2]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5641 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u363 (
    .a(\u2_Display/n4911 [0]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [0]),
    .o(\u2_Display/n6101 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3630 (
    .a(\u2_Display/n5605 ),
    .b(\u2_Display/n5611 [3]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5640 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3631 (
    .a(\u2_Display/n5604 ),
    .b(\u2_Display/n5611 [4]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5639 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3632 (
    .a(\u2_Display/n5603 ),
    .b(\u2_Display/n5611 [5]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5638 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3633 (
    .a(\u2_Display/n5602 ),
    .b(\u2_Display/n5611 [6]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5637 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3634 (
    .a(\u2_Display/n5601 ),
    .b(\u2_Display/n5611 [7]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5636 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3635 (
    .a(\u2_Display/n5600 ),
    .b(\u2_Display/n5611 [8]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5635 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3636 (
    .a(\u2_Display/n5599 ),
    .b(\u2_Display/n5611 [9]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5634 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3637 (
    .a(\u2_Display/n5598 ),
    .b(\u2_Display/n5611 [10]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5633 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3638 (
    .a(\u2_Display/n5597 ),
    .b(\u2_Display/n5611 [11]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5632 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3639 (
    .a(\u2_Display/n5596 ),
    .b(\u2_Display/n5611 [12]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5631 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u364 (
    .a(\u2_Display/n4911 [1]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [1]),
    .o(\u2_Display/n6100 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3640 (
    .a(\u2_Display/n5595 ),
    .b(\u2_Display/n5611 [13]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5630 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3641 (
    .a(\u2_Display/n5594 ),
    .b(\u2_Display/n5611 [14]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5629 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3642 (
    .a(\u2_Display/n5593 ),
    .b(\u2_Display/n5611 [15]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5628 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3643 (
    .a(\u2_Display/n5592 ),
    .b(\u2_Display/n5611 [16]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5627 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3644 (
    .a(\u2_Display/n5591 ),
    .b(\u2_Display/n5611 [17]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5626 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3645 (
    .a(\u2_Display/n5590 ),
    .b(\u2_Display/n5611 [18]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5625 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3646 (
    .a(\u2_Display/n5589 ),
    .b(\u2_Display/n5611 [19]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5624 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3647 (
    .a(\u2_Display/n5588 ),
    .b(\u2_Display/n5611 [20]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5623 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3648 (
    .a(\u2_Display/n5587 ),
    .b(\u2_Display/n5611 [21]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5622 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3649 (
    .a(\u2_Display/n5586 ),
    .b(\u2_Display/n5611 [22]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5621 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u365 (
    .a(\u2_Display/n4911 [2]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [2]),
    .o(\u2_Display/n6099 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3650 (
    .a(\u2_Display/n5585 ),
    .b(\u2_Display/n5611 [23]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5620 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3651 (
    .a(\u2_Display/n5584 ),
    .b(\u2_Display/n5611 [24]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5619 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3652 (
    .a(\u2_Display/n5583 ),
    .b(\u2_Display/n5611 [25]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5618 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3653 (
    .a(\u2_Display/n5582 ),
    .b(\u2_Display/n5611 [26]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5617 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3654 (
    .a(\u2_Display/n5581 ),
    .b(\u2_Display/n5611 [27]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5616 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3655 (
    .a(\u2_Display/n5580 ),
    .b(\u2_Display/n5611 [28]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5615 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3656 (
    .a(\u2_Display/n5579 ),
    .b(\u2_Display/n5611 [29]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5614 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3657 (
    .a(\u2_Display/n5578 ),
    .b(\u2_Display/n5611 [30]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5613 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3658 (
    .a(\u2_Display/n5577 ),
    .b(\u2_Display/n5611 [31]),
    .c(\u2_Display/n5609 ),
    .o(\u2_Display/n5612 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3659 (
    .a(\u2_Display/n1116 ),
    .b(\u2_Display/n1119 [0]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1151 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u366 (
    .a(\u2_Display/n4911 [3]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [3]),
    .o(\u2_Display/n6098 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3660 (
    .a(\u2_Display/n1115 ),
    .b(\u2_Display/n1119 [1]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1150 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3661 (
    .a(\u2_Display/n1114 ),
    .b(\u2_Display/n1119 [2]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1149 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3662 (
    .a(\u2_Display/n1113 ),
    .b(\u2_Display/n1119 [3]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1148 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3663 (
    .a(\u2_Display/n1112 ),
    .b(\u2_Display/n1119 [4]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1147 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3664 (
    .a(\u2_Display/n1111 ),
    .b(\u2_Display/n1119 [5]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1146 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3665 (
    .a(\u2_Display/n1110 ),
    .b(\u2_Display/n1119 [6]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1145 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3666 (
    .a(\u2_Display/n1109 ),
    .b(\u2_Display/n1119 [7]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1144 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3667 (
    .a(\u2_Display/n1108 ),
    .b(\u2_Display/n1119 [8]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1143 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3668 (
    .a(\u2_Display/n1107 ),
    .b(\u2_Display/n1119 [9]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1142 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3669 (
    .a(\u2_Display/n1106 ),
    .b(\u2_Display/n1119 [10]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1141 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u367 (
    .a(\u2_Display/n4911 [4]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [4]),
    .o(\u2_Display/n6097 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3670 (
    .a(\u2_Display/n1105 ),
    .b(\u2_Display/n1119 [11]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1140 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3671 (
    .a(\u2_Display/n1104 ),
    .b(\u2_Display/n1119 [12]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1139 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3672 (
    .a(\u2_Display/n1103 ),
    .b(\u2_Display/n1119 [13]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1138 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3673 (
    .a(\u2_Display/n1102 ),
    .b(\u2_Display/n1119 [14]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1137 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3674 (
    .a(\u2_Display/n1101 ),
    .b(\u2_Display/n1119 [15]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1136 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3675 (
    .a(\u2_Display/n1100 ),
    .b(\u2_Display/n1119 [16]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1135 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3676 (
    .a(\u2_Display/n1099 ),
    .b(\u2_Display/n1119 [17]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1134 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3677 (
    .a(\u2_Display/n1098 ),
    .b(\u2_Display/n1119 [18]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1133 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3678 (
    .a(\u2_Display/n1097 ),
    .b(\u2_Display/n1119 [19]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1132 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3679 (
    .a(\u2_Display/n1096 ),
    .b(\u2_Display/n1119 [20]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1131 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u368 (
    .a(\u2_Display/n4911 [5]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [5]),
    .o(\u2_Display/n6096 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3680 (
    .a(\u2_Display/n1095 ),
    .b(\u2_Display/n1119 [21]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1130 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3681 (
    .a(\u2_Display/n1094 ),
    .b(\u2_Display/n1119 [22]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1129 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3682 (
    .a(\u2_Display/n1093 ),
    .b(\u2_Display/n1119 [23]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1128 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3683 (
    .a(\u2_Display/n1092 ),
    .b(\u2_Display/n1119 [24]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1127 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3684 (
    .a(\u2_Display/n1091 ),
    .b(\u2_Display/n1119 [25]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1126 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3685 (
    .a(\u2_Display/n1090 ),
    .b(\u2_Display/n1119 [26]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1125 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3686 (
    .a(\u2_Display/n1089 ),
    .b(\u2_Display/n1119 [27]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1124 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3687 (
    .a(\u2_Display/n1088 ),
    .b(\u2_Display/n1119 [28]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1123 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3688 (
    .a(\u2_Display/n1087 ),
    .b(\u2_Display/n1119 [29]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1122 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3689 (
    .a(\u2_Display/n1086 ),
    .b(\u2_Display/n1119 [30]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1121 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u369 (
    .a(\u2_Display/n4911 [6]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [6]),
    .o(\u2_Display/n6095 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3690 (
    .a(\u2_Display/n1085 ),
    .b(\u2_Display/n1119 [31]),
    .c(\u2_Display/n1117 ),
    .o(\u2_Display/n1120 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3691 (
    .a(\u2_Display/n2239 ),
    .b(\u2_Display/n2242 [0]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2274 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3692 (
    .a(\u2_Display/n2238 ),
    .b(\u2_Display/n2242 [1]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2273 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3693 (
    .a(\u2_Display/n2237 ),
    .b(\u2_Display/n2242 [2]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2272 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3694 (
    .a(\u2_Display/n2236 ),
    .b(\u2_Display/n2242 [3]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2271 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3695 (
    .a(\u2_Display/n2235 ),
    .b(\u2_Display/n2242 [4]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2270 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3696 (
    .a(\u2_Display/n2234 ),
    .b(\u2_Display/n2242 [5]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2269 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3697 (
    .a(\u2_Display/n2233 ),
    .b(\u2_Display/n2242 [6]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2268 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3698 (
    .a(\u2_Display/n2232 ),
    .b(\u2_Display/n2242 [7]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2267 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3699 (
    .a(\u2_Display/n2231 ),
    .b(\u2_Display/n2242 [8]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2266 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u370 (
    .a(\u2_Display/n4911 [7]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [7]),
    .o(\u2_Display/n6094 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3700 (
    .a(\u2_Display/n2230 ),
    .b(\u2_Display/n2242 [9]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2265 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3701 (
    .a(\u2_Display/n2229 ),
    .b(\u2_Display/n2242 [10]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2264 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3702 (
    .a(\u2_Display/n2228 ),
    .b(\u2_Display/n2242 [11]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2263 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3703 (
    .a(\u2_Display/n2227 ),
    .b(\u2_Display/n2242 [12]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2262 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3704 (
    .a(\u2_Display/n2226 ),
    .b(\u2_Display/n2242 [13]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2261 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3705 (
    .a(\u2_Display/n2225 ),
    .b(\u2_Display/n2242 [14]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2260 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3706 (
    .a(\u2_Display/n2224 ),
    .b(\u2_Display/n2242 [15]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2259 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3707 (
    .a(\u2_Display/n2223 ),
    .b(\u2_Display/n2242 [16]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2258 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3708 (
    .a(\u2_Display/n2222 ),
    .b(\u2_Display/n2242 [17]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2257 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3709 (
    .a(\u2_Display/n2221 ),
    .b(\u2_Display/n2242 [18]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2256 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u371 (
    .a(\u2_Display/n4911 [8]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [8]),
    .o(\u2_Display/n6093 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3710 (
    .a(\u2_Display/n2220 ),
    .b(\u2_Display/n2242 [19]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2255 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3711 (
    .a(\u2_Display/n2219 ),
    .b(\u2_Display/n2242 [20]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2254 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3712 (
    .a(\u2_Display/n2218 ),
    .b(\u2_Display/n2242 [21]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2253 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3713 (
    .a(\u2_Display/n2217 ),
    .b(\u2_Display/n2242 [22]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2252 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3714 (
    .a(\u2_Display/n2216 ),
    .b(\u2_Display/n2242 [23]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2251 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3715 (
    .a(\u2_Display/n2215 ),
    .b(\u2_Display/n2242 [24]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2250 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3716 (
    .a(\u2_Display/n2214 ),
    .b(\u2_Display/n2242 [25]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2249 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3717 (
    .a(\u2_Display/n2213 ),
    .b(\u2_Display/n2242 [26]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2248 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3718 (
    .a(\u2_Display/n2212 ),
    .b(\u2_Display/n2242 [27]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2247 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3719 (
    .a(\u2_Display/n2211 ),
    .b(\u2_Display/n2242 [28]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2246 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u372 (
    .a(\u2_Display/n4911 [9]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [9]),
    .o(\u2_Display/n6092 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3720 (
    .a(\u2_Display/n2210 ),
    .b(\u2_Display/n2242 [29]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2245 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3721 (
    .a(\u2_Display/n2209 ),
    .b(\u2_Display/n2242 [30]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2244 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3722 (
    .a(\u2_Display/n2208 ),
    .b(\u2_Display/n2242 [31]),
    .c(\u2_Display/n2240 ),
    .o(\u2_Display/n2243 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3723 (
    .a(\u2_Display/n3362 ),
    .b(\u2_Display/n3365 [0]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3397 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3724 (
    .a(\u2_Display/n3361 ),
    .b(\u2_Display/n3365 [1]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3396 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3725 (
    .a(\u2_Display/n3360 ),
    .b(\u2_Display/n3365 [2]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3395 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3726 (
    .a(\u2_Display/n3359 ),
    .b(\u2_Display/n3365 [3]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3394 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3727 (
    .a(\u2_Display/n3358 ),
    .b(\u2_Display/n3365 [4]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3393 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3728 (
    .a(\u2_Display/n3357 ),
    .b(\u2_Display/n3365 [5]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3392 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3729 (
    .a(\u2_Display/n3356 ),
    .b(\u2_Display/n3365 [6]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3391 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u373 (
    .a(\u2_Display/n4911 [10]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [10]),
    .o(\u2_Display/n6091 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3730 (
    .a(\u2_Display/n3355 ),
    .b(\u2_Display/n3365 [7]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3390 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3731 (
    .a(\u2_Display/n3354 ),
    .b(\u2_Display/n3365 [8]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3389 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3732 (
    .a(\u2_Display/n3353 ),
    .b(\u2_Display/n3365 [9]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3388 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3733 (
    .a(\u2_Display/n3352 ),
    .b(\u2_Display/n3365 [10]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3387 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3734 (
    .a(\u2_Display/n3351 ),
    .b(\u2_Display/n3365 [11]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3386 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3735 (
    .a(\u2_Display/n3350 ),
    .b(\u2_Display/n3365 [12]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3385 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3736 (
    .a(\u2_Display/n3349 ),
    .b(\u2_Display/n3365 [13]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3384 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3737 (
    .a(\u2_Display/n3348 ),
    .b(\u2_Display/n3365 [14]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3383 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3738 (
    .a(\u2_Display/n3347 ),
    .b(\u2_Display/n3365 [15]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3382 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3739 (
    .a(\u2_Display/n3346 ),
    .b(\u2_Display/n3365 [16]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3381 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u374 (
    .a(\u2_Display/n4911 [11]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [11]),
    .o(\u2_Display/n6090 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3740 (
    .a(\u2_Display/n3345 ),
    .b(\u2_Display/n3365 [17]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3380 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3741 (
    .a(\u2_Display/n3344 ),
    .b(\u2_Display/n3365 [18]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3379 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3742 (
    .a(\u2_Display/n3343 ),
    .b(\u2_Display/n3365 [19]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3378 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3743 (
    .a(\u2_Display/n3342 ),
    .b(\u2_Display/n3365 [20]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3377 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3744 (
    .a(\u2_Display/n3341 ),
    .b(\u2_Display/n3365 [21]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3376 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3745 (
    .a(\u2_Display/n3340 ),
    .b(\u2_Display/n3365 [22]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3375 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3746 (
    .a(\u2_Display/n3339 ),
    .b(\u2_Display/n3365 [23]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3374 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3747 (
    .a(\u2_Display/n3338 ),
    .b(\u2_Display/n3365 [24]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3373 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3748 (
    .a(\u2_Display/n3337 ),
    .b(\u2_Display/n3365 [25]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3372 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3749 (
    .a(\u2_Display/n3336 ),
    .b(\u2_Display/n3365 [26]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3371 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u375 (
    .a(\u2_Display/n4911 [12]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [12]),
    .o(\u2_Display/n6089 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3750 (
    .a(\u2_Display/n3335 ),
    .b(\u2_Display/n3365 [27]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3370 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3751 (
    .a(\u2_Display/n3334 ),
    .b(\u2_Display/n3365 [28]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3369 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3752 (
    .a(\u2_Display/n3333 ),
    .b(\u2_Display/n3365 [29]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3368 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3753 (
    .a(\u2_Display/n3332 ),
    .b(\u2_Display/n3365 [30]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3367 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3754 (
    .a(\u2_Display/n3331 ),
    .b(\u2_Display/n3365 [31]),
    .c(\u2_Display/n3363 ),
    .o(\u2_Display/n3366 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3755 (
    .a(\u2_Display/n4520 ),
    .b(\u2_Display/n4523 [0]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4555 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3756 (
    .a(\u2_Display/n4519 ),
    .b(\u2_Display/n4523 [1]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4554 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3757 (
    .a(\u2_Display/n4518 ),
    .b(\u2_Display/n4523 [2]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4553 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3758 (
    .a(\u2_Display/n4517 ),
    .b(\u2_Display/n4523 [3]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4552 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3759 (
    .a(\u2_Display/n4516 ),
    .b(\u2_Display/n4523 [4]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4551 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u376 (
    .a(\u2_Display/n4911 [13]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [13]),
    .o(\u2_Display/n6088 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3760 (
    .a(\u2_Display/n4515 ),
    .b(\u2_Display/n4523 [5]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4550 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3761 (
    .a(\u2_Display/n4514 ),
    .b(\u2_Display/n4523 [6]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4549 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3762 (
    .a(\u2_Display/n4513 ),
    .b(\u2_Display/n4523 [7]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4548 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3763 (
    .a(\u2_Display/n4512 ),
    .b(\u2_Display/n4523 [8]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4547 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3764 (
    .a(\u2_Display/n4511 ),
    .b(\u2_Display/n4523 [9]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4546 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3765 (
    .a(\u2_Display/n4510 ),
    .b(\u2_Display/n4523 [10]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4545 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3766 (
    .a(\u2_Display/n4509 ),
    .b(\u2_Display/n4523 [11]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4544 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3767 (
    .a(\u2_Display/n4508 ),
    .b(\u2_Display/n4523 [12]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4543 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3768 (
    .a(\u2_Display/n4507 ),
    .b(\u2_Display/n4523 [13]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4542 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3769 (
    .a(\u2_Display/n4506 ),
    .b(\u2_Display/n4523 [14]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4541 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u377 (
    .a(\u2_Display/n4911 [14]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [14]),
    .o(\u2_Display/n6087 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3770 (
    .a(\u2_Display/n4505 ),
    .b(\u2_Display/n4523 [15]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4540 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3771 (
    .a(\u2_Display/n4504 ),
    .b(\u2_Display/n4523 [16]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4539 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3772 (
    .a(\u2_Display/n4503 ),
    .b(\u2_Display/n4523 [17]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4538 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3773 (
    .a(\u2_Display/n4502 ),
    .b(\u2_Display/n4523 [18]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4537 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3774 (
    .a(\u2_Display/n4501 ),
    .b(\u2_Display/n4523 [19]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4536 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3775 (
    .a(\u2_Display/n4500 ),
    .b(\u2_Display/n4523 [20]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4535 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3776 (
    .a(\u2_Display/n4499 ),
    .b(\u2_Display/n4523 [21]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4534 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3777 (
    .a(\u2_Display/n4498 ),
    .b(\u2_Display/n4523 [22]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4533 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3778 (
    .a(\u2_Display/n4497 ),
    .b(\u2_Display/n4523 [23]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4532 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3779 (
    .a(\u2_Display/n4496 ),
    .b(\u2_Display/n4523 [24]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4531 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u378 (
    .a(\u2_Display/n4911 [15]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [15]),
    .o(\u2_Display/n6086 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3780 (
    .a(\u2_Display/n4495 ),
    .b(\u2_Display/n4523 [25]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4530 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3781 (
    .a(\u2_Display/n4494 ),
    .b(\u2_Display/n4523 [26]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4529 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3782 (
    .a(\u2_Display/n4493 ),
    .b(\u2_Display/n4523 [27]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4528 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3783 (
    .a(\u2_Display/n4492 ),
    .b(\u2_Display/n4523 [28]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4527 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3784 (
    .a(\u2_Display/n4491 ),
    .b(\u2_Display/n4523 [29]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4526 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3785 (
    .a(\u2_Display/n4490 ),
    .b(\u2_Display/n4523 [30]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4525 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3786 (
    .a(\u2_Display/n4489 ),
    .b(\u2_Display/n4523 [31]),
    .c(\u2_Display/n4521 ),
    .o(\u2_Display/n4524 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3787 (
    .a(\u2_Display/n5643 ),
    .b(\u2_Display/n5646 [0]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5678 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3788 (
    .a(\u2_Display/n5642 ),
    .b(\u2_Display/n5646 [1]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5677 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3789 (
    .a(\u2_Display/n5641 ),
    .b(\u2_Display/n5646 [2]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5676 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u379 (
    .a(\u2_Display/n4911 [16]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [16]),
    .o(\u2_Display/n6085 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3790 (
    .a(\u2_Display/n5640 ),
    .b(\u2_Display/n5646 [3]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5675 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3791 (
    .a(\u2_Display/n5639 ),
    .b(\u2_Display/n5646 [4]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5674 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3792 (
    .a(\u2_Display/n5638 ),
    .b(\u2_Display/n5646 [5]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5673 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3793 (
    .a(\u2_Display/n5637 ),
    .b(\u2_Display/n5646 [6]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5672 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3794 (
    .a(\u2_Display/n5636 ),
    .b(\u2_Display/n5646 [7]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5671 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3795 (
    .a(\u2_Display/n5635 ),
    .b(\u2_Display/n5646 [8]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5670 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3796 (
    .a(\u2_Display/n5634 ),
    .b(\u2_Display/n5646 [9]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5669 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3797 (
    .a(\u2_Display/n5633 ),
    .b(\u2_Display/n5646 [10]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5668 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3798 (
    .a(\u2_Display/n5632 ),
    .b(\u2_Display/n5646 [11]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5667 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3799 (
    .a(\u2_Display/n5631 ),
    .b(\u2_Display/n5646 [12]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5666 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u380 (
    .a(\u2_Display/n4911 [17]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [17]),
    .o(\u2_Display/n6084 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3800 (
    .a(\u2_Display/n5630 ),
    .b(\u2_Display/n5646 [13]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5665 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3801 (
    .a(\u2_Display/n5629 ),
    .b(\u2_Display/n5646 [14]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5664 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3802 (
    .a(\u2_Display/n5628 ),
    .b(\u2_Display/n5646 [15]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5663 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3803 (
    .a(\u2_Display/n5627 ),
    .b(\u2_Display/n5646 [16]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5662 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3804 (
    .a(\u2_Display/n5626 ),
    .b(\u2_Display/n5646 [17]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5661 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3805 (
    .a(\u2_Display/n5625 ),
    .b(\u2_Display/n5646 [18]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5660 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3806 (
    .a(\u2_Display/n5624 ),
    .b(\u2_Display/n5646 [19]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5659 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3807 (
    .a(\u2_Display/n5623 ),
    .b(\u2_Display/n5646 [20]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5658 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3808 (
    .a(\u2_Display/n5622 ),
    .b(\u2_Display/n5646 [21]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5657 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3809 (
    .a(\u2_Display/n5621 ),
    .b(\u2_Display/n5646 [22]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5656 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u381 (
    .a(\u2_Display/n4911 [18]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [18]),
    .o(\u2_Display/n6083 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3810 (
    .a(\u2_Display/n5620 ),
    .b(\u2_Display/n5646 [23]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5655 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3811 (
    .a(\u2_Display/n5619 ),
    .b(\u2_Display/n5646 [24]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5654 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3812 (
    .a(\u2_Display/n5618 ),
    .b(\u2_Display/n5646 [25]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5653 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3813 (
    .a(\u2_Display/n5617 ),
    .b(\u2_Display/n5646 [26]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5652 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3814 (
    .a(\u2_Display/n5616 ),
    .b(\u2_Display/n5646 [27]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5651 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3815 (
    .a(\u2_Display/n5615 ),
    .b(\u2_Display/n5646 [28]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5650 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3816 (
    .a(\u2_Display/n5614 ),
    .b(\u2_Display/n5646 [29]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5649 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3817 (
    .a(\u2_Display/n5613 ),
    .b(\u2_Display/n5646 [30]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5648 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3818 (
    .a(\u2_Display/n5612 ),
    .b(\u2_Display/n5646 [31]),
    .c(\u2_Display/n5644 ),
    .o(\u2_Display/n5647 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3819 (
    .a(\u2_Display/n1151 ),
    .b(\u2_Display/n1154 [0]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1186 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u382 (
    .a(\u2_Display/n4911 [19]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [19]),
    .o(\u2_Display/n6082 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3820 (
    .a(\u2_Display/n1150 ),
    .b(\u2_Display/n1154 [1]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1185 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3821 (
    .a(\u2_Display/n1149 ),
    .b(\u2_Display/n1154 [2]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1184 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3822 (
    .a(\u2_Display/n1148 ),
    .b(\u2_Display/n1154 [3]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1183 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3823 (
    .a(\u2_Display/n1147 ),
    .b(\u2_Display/n1154 [4]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1182 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3824 (
    .a(\u2_Display/n1146 ),
    .b(\u2_Display/n1154 [5]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1181 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3825 (
    .a(\u2_Display/n1145 ),
    .b(\u2_Display/n1154 [6]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1180 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3826 (
    .a(\u2_Display/n1144 ),
    .b(\u2_Display/n1154 [7]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1179 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3827 (
    .a(\u2_Display/n1143 ),
    .b(\u2_Display/n1154 [8]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1178 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3828 (
    .a(\u2_Display/n1142 ),
    .b(\u2_Display/n1154 [9]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1177 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3829 (
    .a(\u2_Display/n1141 ),
    .b(\u2_Display/n1154 [10]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1176 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u383 (
    .a(\u2_Display/n4911 [20]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [20]),
    .o(\u2_Display/n6081 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3830 (
    .a(\u2_Display/n1140 ),
    .b(\u2_Display/n1154 [11]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1175 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3831 (
    .a(\u2_Display/n1139 ),
    .b(\u2_Display/n1154 [12]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1174 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3832 (
    .a(\u2_Display/n1138 ),
    .b(\u2_Display/n1154 [13]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1173 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3833 (
    .a(\u2_Display/n1137 ),
    .b(\u2_Display/n1154 [14]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1172 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3834 (
    .a(\u2_Display/n1136 ),
    .b(\u2_Display/n1154 [15]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1171 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3835 (
    .a(\u2_Display/n1135 ),
    .b(\u2_Display/n1154 [16]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1170 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3836 (
    .a(\u2_Display/n1134 ),
    .b(\u2_Display/n1154 [17]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1169 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3837 (
    .a(\u2_Display/n1133 ),
    .b(\u2_Display/n1154 [18]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1168 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3838 (
    .a(\u2_Display/n1132 ),
    .b(\u2_Display/n1154 [19]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1167 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3839 (
    .a(\u2_Display/n1131 ),
    .b(\u2_Display/n1154 [20]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1166 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u384 (
    .a(\u2_Display/n4911 [21]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [21]),
    .o(\u2_Display/n6080 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3840 (
    .a(\u2_Display/n1130 ),
    .b(\u2_Display/n1154 [21]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1165 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3841 (
    .a(\u2_Display/n1129 ),
    .b(\u2_Display/n1154 [22]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1164 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3842 (
    .a(\u2_Display/n1128 ),
    .b(\u2_Display/n1154 [23]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1163 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3843 (
    .a(\u2_Display/n1127 ),
    .b(\u2_Display/n1154 [24]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1162 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3844 (
    .a(\u2_Display/n1126 ),
    .b(\u2_Display/n1154 [25]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1161 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3845 (
    .a(\u2_Display/n1125 ),
    .b(\u2_Display/n1154 [26]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1160 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3846 (
    .a(\u2_Display/n1124 ),
    .b(\u2_Display/n1154 [27]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1159 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3847 (
    .a(\u2_Display/n1123 ),
    .b(\u2_Display/n1154 [28]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1158 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3848 (
    .a(\u2_Display/n1122 ),
    .b(\u2_Display/n1154 [29]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1157 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3849 (
    .a(\u2_Display/n1121 ),
    .b(\u2_Display/n1154 [30]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1156 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u385 (
    .a(\u2_Display/n4911 [22]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [22]),
    .o(\u2_Display/n6079 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3850 (
    .a(\u2_Display/n1120 ),
    .b(\u2_Display/n1154 [31]),
    .c(\u2_Display/n1152 ),
    .o(\u2_Display/n1155 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3851 (
    .a(\u2_Display/n2274 ),
    .b(\u2_Display/n2277 [0]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2309 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3852 (
    .a(\u2_Display/n2273 ),
    .b(\u2_Display/n2277 [1]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2308 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3853 (
    .a(\u2_Display/n2272 ),
    .b(\u2_Display/n2277 [2]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2307 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3854 (
    .a(\u2_Display/n2271 ),
    .b(\u2_Display/n2277 [3]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2306 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3855 (
    .a(\u2_Display/n2270 ),
    .b(\u2_Display/n2277 [4]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2305 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3856 (
    .a(\u2_Display/n2269 ),
    .b(\u2_Display/n2277 [5]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2304 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3857 (
    .a(\u2_Display/n2268 ),
    .b(\u2_Display/n2277 [6]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2303 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3858 (
    .a(\u2_Display/n2267 ),
    .b(\u2_Display/n2277 [7]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2302 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3859 (
    .a(\u2_Display/n2266 ),
    .b(\u2_Display/n2277 [8]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2301 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u386 (
    .a(\u2_Display/n4911 [23]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [23]),
    .o(\u2_Display/n6078 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3860 (
    .a(\u2_Display/n2265 ),
    .b(\u2_Display/n2277 [9]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2300 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3861 (
    .a(\u2_Display/n2264 ),
    .b(\u2_Display/n2277 [10]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2299 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3862 (
    .a(\u2_Display/n2263 ),
    .b(\u2_Display/n2277 [11]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2298 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3863 (
    .a(\u2_Display/n2262 ),
    .b(\u2_Display/n2277 [12]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2297 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3864 (
    .a(\u2_Display/n2261 ),
    .b(\u2_Display/n2277 [13]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2296 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3865 (
    .a(\u2_Display/n2260 ),
    .b(\u2_Display/n2277 [14]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2295 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3866 (
    .a(\u2_Display/n2259 ),
    .b(\u2_Display/n2277 [15]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2294 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3867 (
    .a(\u2_Display/n2258 ),
    .b(\u2_Display/n2277 [16]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2293 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3868 (
    .a(\u2_Display/n2257 ),
    .b(\u2_Display/n2277 [17]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2292 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3869 (
    .a(\u2_Display/n2256 ),
    .b(\u2_Display/n2277 [18]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2291 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u387 (
    .a(\u2_Display/n4911 [24]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [24]),
    .o(\u2_Display/n6077 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3870 (
    .a(\u2_Display/n2255 ),
    .b(\u2_Display/n2277 [19]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2290 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3871 (
    .a(\u2_Display/n2254 ),
    .b(\u2_Display/n2277 [20]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2289 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3872 (
    .a(\u2_Display/n2253 ),
    .b(\u2_Display/n2277 [21]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2288 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3873 (
    .a(\u2_Display/n2252 ),
    .b(\u2_Display/n2277 [22]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2287 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3874 (
    .a(\u2_Display/n2251 ),
    .b(\u2_Display/n2277 [23]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2286 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3875 (
    .a(\u2_Display/n2250 ),
    .b(\u2_Display/n2277 [24]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2285 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3876 (
    .a(\u2_Display/n2249 ),
    .b(\u2_Display/n2277 [25]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2284 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3877 (
    .a(\u2_Display/n2248 ),
    .b(\u2_Display/n2277 [26]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2283 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3878 (
    .a(\u2_Display/n2247 ),
    .b(\u2_Display/n2277 [27]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2282 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3879 (
    .a(\u2_Display/n2246 ),
    .b(\u2_Display/n2277 [28]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2281 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u388 (
    .a(\u2_Display/n4911 [25]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [25]),
    .o(\u2_Display/n6076 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3880 (
    .a(\u2_Display/n2245 ),
    .b(\u2_Display/n2277 [29]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2280 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3881 (
    .a(\u2_Display/n2244 ),
    .b(\u2_Display/n2277 [30]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2279 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3882 (
    .a(\u2_Display/n2243 ),
    .b(\u2_Display/n2277 [31]),
    .c(\u2_Display/n2275 ),
    .o(\u2_Display/n2278 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3883 (
    .a(\u2_Display/n3397 ),
    .b(\u2_Display/n3400 [0]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3432 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3884 (
    .a(\u2_Display/n3396 ),
    .b(\u2_Display/n3400 [1]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3431 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3885 (
    .a(\u2_Display/n3395 ),
    .b(\u2_Display/n3400 [2]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3430 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3886 (
    .a(\u2_Display/n3394 ),
    .b(\u2_Display/n3400 [3]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3429 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3887 (
    .a(\u2_Display/n3393 ),
    .b(\u2_Display/n3400 [4]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3428 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3888 (
    .a(\u2_Display/n3392 ),
    .b(\u2_Display/n3400 [5]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3427 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3889 (
    .a(\u2_Display/n3391 ),
    .b(\u2_Display/n3400 [6]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3426 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u389 (
    .a(\u2_Display/n4911 [26]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [26]),
    .o(\u2_Display/n6075 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3890 (
    .a(\u2_Display/n3390 ),
    .b(\u2_Display/n3400 [7]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3425 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3891 (
    .a(\u2_Display/n3389 ),
    .b(\u2_Display/n3400 [8]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3424 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3892 (
    .a(\u2_Display/n3388 ),
    .b(\u2_Display/n3400 [9]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3423 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3893 (
    .a(\u2_Display/n3387 ),
    .b(\u2_Display/n3400 [10]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3422 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3894 (
    .a(\u2_Display/n3386 ),
    .b(\u2_Display/n3400 [11]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3421 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3895 (
    .a(\u2_Display/n3385 ),
    .b(\u2_Display/n3400 [12]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3420 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3896 (
    .a(\u2_Display/n3384 ),
    .b(\u2_Display/n3400 [13]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3419 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3897 (
    .a(\u2_Display/n3383 ),
    .b(\u2_Display/n3400 [14]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3418 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3898 (
    .a(\u2_Display/n3382 ),
    .b(\u2_Display/n3400 [15]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3417 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3899 (
    .a(\u2_Display/n3381 ),
    .b(\u2_Display/n3400 [16]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3416 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u390 (
    .a(\u2_Display/n4911 [27]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [27]),
    .o(\u2_Display/n6074 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3900 (
    .a(\u2_Display/n3380 ),
    .b(\u2_Display/n3400 [17]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3415 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3901 (
    .a(\u2_Display/n3379 ),
    .b(\u2_Display/n3400 [18]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3414 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3902 (
    .a(\u2_Display/n3378 ),
    .b(\u2_Display/n3400 [19]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3413 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3903 (
    .a(\u2_Display/n3377 ),
    .b(\u2_Display/n3400 [20]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3412 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3904 (
    .a(\u2_Display/n3376 ),
    .b(\u2_Display/n3400 [21]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3411 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3905 (
    .a(\u2_Display/n3375 ),
    .b(\u2_Display/n3400 [22]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3410 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3906 (
    .a(\u2_Display/n3374 ),
    .b(\u2_Display/n3400 [23]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3409 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3907 (
    .a(\u2_Display/n3373 ),
    .b(\u2_Display/n3400 [24]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3408 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3908 (
    .a(\u2_Display/n3372 ),
    .b(\u2_Display/n3400 [25]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3407 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3909 (
    .a(\u2_Display/n3371 ),
    .b(\u2_Display/n3400 [26]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3406 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u391 (
    .a(\u2_Display/n4911 [28]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [28]),
    .o(\u2_Display/n6073 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3910 (
    .a(\u2_Display/n3370 ),
    .b(\u2_Display/n3400 [27]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3405 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3911 (
    .a(\u2_Display/n3369 ),
    .b(\u2_Display/n3400 [28]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3404 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3912 (
    .a(\u2_Display/n3368 ),
    .b(\u2_Display/n3400 [29]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3403 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3913 (
    .a(\u2_Display/n3367 ),
    .b(\u2_Display/n3400 [30]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3402 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3914 (
    .a(\u2_Display/n3366 ),
    .b(\u2_Display/n3400 [31]),
    .c(\u2_Display/n3398 ),
    .o(\u2_Display/n3401 ));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*B)*~(C*A))"),
    .INIT(16'heca0))
    _al_u3915 (
    .a(\u2_Display/n5668 ),
    .b(_al_u1168_o),
    .c(on_off_pad[0]),
    .d(\u2_Display/i [10]),
    .o(\u2_Display/n238 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3916 (
    .a(\u2_Display/n3432 ),
    .b(\u2_Display/n3435 [0]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3916_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3917 (
    .a(\u2_Display/n1186 ),
    .b(\u2_Display/n1189 [0]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3917_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3918 (
    .a(_al_u3916_o),
    .b(_al_u3917_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [0]),
    .o(_al_u3918_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3919 (
    .a(_al_u3918_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [0]),
    .o(\u2_Display/n239 [0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u392 (
    .a(\u2_Display/n4911 [29]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [29]),
    .o(\u2_Display/n6072 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3920 (
    .a(\u2_Display/n3431 ),
    .b(\u2_Display/n3435 [1]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3920_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3921 (
    .a(\u2_Display/n1185 ),
    .b(\u2_Display/n1189 [1]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3921_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3922 (
    .a(_al_u3920_o),
    .b(_al_u3921_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [1]),
    .o(_al_u3922_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3923 (
    .a(_al_u3922_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [1]),
    .o(\u2_Display/n239 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3924 (
    .a(\u2_Display/n1184 ),
    .b(\u2_Display/n1189 [2]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3924_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3925 (
    .a(\u2_Display/n3430 ),
    .b(\u2_Display/n3435 [2]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3925_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~((E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D))*~(C)+B*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*~(C)+~(B)*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*C+B*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*C)"),
    .INIT(32'hacfcac0c))
    _al_u3926 (
    .a(_al_u3924_o),
    .b(_al_u3925_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [2]),
    .o(_al_u3926_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u3927 (
    .a(_al_u3926_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [2]),
    .o(\u2_Display/n239 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3928 (
    .a(\u2_Display/n3429 ),
    .b(\u2_Display/n3435 [3]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3928_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3929 (
    .a(\u2_Display/n1183 ),
    .b(\u2_Display/n1189 [3]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3929_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u393 (
    .a(\u2_Display/n4911 [30]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [30]),
    .o(\u2_Display/n6071 ));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3930 (
    .a(_al_u3928_o),
    .b(_al_u3929_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [3]),
    .o(_al_u3930_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3931 (
    .a(_al_u3930_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [3]),
    .o(\u2_Display/n239 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3932 (
    .a(\u2_Display/n3428 ),
    .b(\u2_Display/n3435 [4]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3932_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3933 (
    .a(\u2_Display/n1182 ),
    .b(\u2_Display/n1189 [4]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3933_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3934 (
    .a(_al_u3932_o),
    .b(_al_u3933_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [4]),
    .o(_al_u3934_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3935 (
    .a(_al_u3934_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [4]),
    .o(\u2_Display/n239 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3936 (
    .a(\u2_Display/n3427 ),
    .b(\u2_Display/n3435 [5]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3936_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3937 (
    .a(\u2_Display/n1181 ),
    .b(\u2_Display/n1189 [5]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3937_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3938 (
    .a(_al_u3936_o),
    .b(_al_u3937_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [5]),
    .o(_al_u3938_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3939 (
    .a(_al_u3938_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [5]),
    .o(\u2_Display/n239 [5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u394 (
    .a(\u2_Display/n4911 [31]),
    .b(\u2_Display/n4909 ),
    .c(\u2_Display/counta [31]),
    .o(\u2_Display/n6070 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3940 (
    .a(\u2_Display/n1180 ),
    .b(\u2_Display/n1189 [6]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3940_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3941 (
    .a(\u2_Display/n3426 ),
    .b(\u2_Display/n3435 [6]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3941_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~((E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D))*~(C)+B*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*~(C)+~(B)*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*C+B*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*C)"),
    .INIT(32'hacfcac0c))
    _al_u3942 (
    .a(_al_u3940_o),
    .b(_al_u3941_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [6]),
    .o(_al_u3942_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u3943 (
    .a(_al_u3942_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [6]),
    .o(\u2_Display/n239 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3944 (
    .a(\u2_Display/n3425 ),
    .b(\u2_Display/n3435 [7]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3944_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3945 (
    .a(\u2_Display/n1179 ),
    .b(\u2_Display/n1189 [7]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3945_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3946 (
    .a(_al_u3944_o),
    .b(_al_u3945_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [7]),
    .o(_al_u3946_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h74))
    _al_u3947 (
    .a(_al_u3946_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [7]),
    .o(\u2_Display/n239 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3948 (
    .a(\u2_Display/n1178 ),
    .b(\u2_Display/n1189 [8]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3948_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3949 (
    .a(\u2_Display/n3424 ),
    .b(\u2_Display/n3435 [8]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3949_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u395 (
    .a(\u2_Display/n419 [0]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [0]),
    .o(\u2_Display/n451 ));
  AL_MAP_LUT5 #(
    .EQN("(B*~((E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D))*~(C)+B*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*~(C)+~(B)*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*C+B*(E*~(A)*~(D)+E*A*~(D)+~(E)*A*D+E*A*D)*C)"),
    .INIT(32'hacfcac0c))
    _al_u3950 (
    .a(_al_u3948_o),
    .b(_al_u3949_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [8]),
    .o(_al_u3950_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u3951 (
    .a(_al_u3950_o),
    .b(\u2_Display/mux19_b0_sel_is_0_o ),
    .c(\u2_Display/counta [8]),
    .o(\u2_Display/n239 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3952 (
    .a(\u2_Display/n3423 ),
    .b(\u2_Display/n3435 [9]),
    .c(\u2_Display/n3433 ),
    .o(_al_u3952_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3953 (
    .a(\u2_Display/n1177 ),
    .b(\u2_Display/n1189 [9]),
    .c(\u2_Display/n1187 ),
    .o(_al_u3953_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D))*~(C)+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*~(C)+~(A)*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C+A*(E*~(B)*~(D)+E*B*~(D)+~(E)*B*D+E*B*D)*C)"),
    .INIT(32'h350535f5))
    _al_u3954 (
    .a(_al_u3952_o),
    .b(_al_u3953_o),
    .c(\u2_Display/mux11_b0_sel_is_0_o ),
    .d(on_off_pad[4]),
    .e(\u2_Display/j [9]),
    .o(_al_u3954_o));
  AL_MAP_LUT4 #(
    .EQN("((~B*~A)*~(D)*~(C)+(~B*~A)*D*~(C)+~((~B*~A))*D*C+(~B*~A)*D*C)"),
    .INIT(16'hf101))
    _al_u3955 (
    .a(_al_u3954_o),
    .b(on_off_pad[1]),
    .c(on_off_pad[0]),
    .d(\u2_Display/counta [9]),
    .o(\u2_Display/n239 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .INIT(16'haab8))
    _al_u3956 (
    .a(\u2_Display/n5678 ),
    .b(on_off_pad[0]),
    .c(\u2_Display/n5681 [0]),
    .d(\u2_Display/n5679 ),
    .o(_al_u3956_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3957 (
    .a(\u2_Display/n2309 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [0]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [0]),
    .o(_al_u3957_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*~(C)+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(C)+~(~A)*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C)"),
    .INIT(32'h3a3a0afa))
    _al_u3958 (
    .a(_al_u3957_o),
    .b(\u2_Display/n4555 ),
    .c(on_off_pad[2]),
    .d(\u2_Display/n4558 [0]),
    .e(\u2_Display/n4556 ),
    .o(_al_u3958_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u3959 (
    .a(_al_u3958_o),
    .b(_al_u3956_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u396 (
    .a(\u2_Display/n419 [1]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [1]),
    .o(\u2_Display/n450 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3960 (
    .a(\u2_Display/n2308 ),
    .b(\u2_Display/n2312 [1]),
    .c(\u2_Display/n2310 ),
    .o(_al_u3960_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3961 (
    .a(\u2_Display/n4554 ),
    .b(\u2_Display/n4558 [1]),
    .c(\u2_Display/n4556 ),
    .o(_al_u3961_o));
  AL_MAP_LUT5 #(
    .EQN("~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'h330533f5))
    _al_u3962 (
    .a(_al_u3960_o),
    .b(_al_u3961_o),
    .c(\u2_Display/mux5_b0_sel_is_0_o ),
    .d(on_off_pad[2]),
    .e(\u2_Display/i [1]),
    .o(_al_u3962_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h5757535f))
    _al_u3963 (
    .a(\u2_Display/n5677 ),
    .b(on_off_pad[1]),
    .c(on_off_pad[0]),
    .d(\u2_Display/n5681 [1]),
    .e(\u2_Display/n5679 ),
    .o(_al_u3963_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u3964 (
    .a(_al_u3962_o),
    .b(_al_u3963_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .INIT(16'haab8))
    _al_u3965 (
    .a(\u2_Display/n5676 ),
    .b(on_off_pad[0]),
    .c(\u2_Display/n5681 [2]),
    .d(\u2_Display/n5679 ),
    .o(_al_u3965_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3966 (
    .a(\u2_Display/n2307 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [2]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [2]),
    .o(_al_u3966_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*~(C)+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(C)+~(~A)*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C)"),
    .INIT(32'h3a3a0afa))
    _al_u3967 (
    .a(_al_u3966_o),
    .b(\u2_Display/n4553 ),
    .c(on_off_pad[2]),
    .d(\u2_Display/n4558 [2]),
    .e(\u2_Display/n4556 ),
    .o(_al_u3967_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u3968 (
    .a(_al_u3967_o),
    .b(_al_u3965_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3969 (
    .a(\u2_Display/n2306 ),
    .b(\u2_Display/n2312 [3]),
    .c(\u2_Display/n2310 ),
    .o(_al_u3969_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u397 (
    .a(\u2_Display/n419 [2]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [2]),
    .o(\u2_Display/n449 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3970 (
    .a(\u2_Display/n4552 ),
    .b(\u2_Display/n4558 [3]),
    .c(\u2_Display/n4556 ),
    .o(_al_u3970_o));
  AL_MAP_LUT5 #(
    .EQN("~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*~(B)*~(D)+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*~(D)+~((A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C))*B*D+(A*~(E)*~(C)+A*E*~(C)+~(A)*E*C+A*E*C)*B*D)"),
    .INIT(32'h330533f5))
    _al_u3971 (
    .a(_al_u3969_o),
    .b(_al_u3970_o),
    .c(\u2_Display/mux5_b0_sel_is_0_o ),
    .d(on_off_pad[2]),
    .e(\u2_Display/i [3]),
    .o(_al_u3971_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h5757535f))
    _al_u3972 (
    .a(\u2_Display/n5675 ),
    .b(on_off_pad[1]),
    .c(on_off_pad[0]),
    .d(\u2_Display/n5681 [3]),
    .e(\u2_Display/n5679 ),
    .o(_al_u3972_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C*~A))"),
    .INIT(8'h73))
    _al_u3973 (
    .a(_al_u3971_o),
    .b(_al_u3972_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3974 (
    .a(\u2_Display/n4551 ),
    .b(\u2_Display/n4558 [4]),
    .c(\u2_Display/n4556 ),
    .o(_al_u3974_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3975 (
    .a(\u2_Display/n2305 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [4]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [4]),
    .o(_al_u3975_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h5757535f))
    _al_u3976 (
    .a(\u2_Display/n5674 ),
    .b(on_off_pad[1]),
    .c(on_off_pad[0]),
    .d(\u2_Display/n5681 [4]),
    .e(\u2_Display/n5679 ),
    .o(_al_u3976_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*(~B*~(A)*~(E)+~B*A*~(E)+~(~B)*A*E+~B*A*E)))"),
    .INIT(32'haf0f3f0f))
    _al_u3977 (
    .a(_al_u3974_o),
    .b(_al_u3975_o),
    .c(_al_u3976_o),
    .d(\u2_Display/mux19_b0_sel_is_0_o ),
    .e(on_off_pad[2]),
    .o(\u2_Display/n238 [4]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hababafa3))
    _al_u3978 (
    .a(\u2_Display/n5673 ),
    .b(on_off_pad[1]),
    .c(on_off_pad[0]),
    .d(\u2_Display/n5681 [5]),
    .e(\u2_Display/n5679 ),
    .o(_al_u3978_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3979 (
    .a(\u2_Display/n2304 ),
    .b(\u2_Display/n2312 [5]),
    .c(\u2_Display/n2310 ),
    .o(_al_u3979_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u398 (
    .a(\u2_Display/n419 [3]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [3]),
    .o(\u2_Display/n448 ));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .INIT(16'h0e02))
    _al_u3980 (
    .a(_al_u3979_o),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(on_off_pad[2]),
    .d(\u2_Display/i [5]),
    .o(_al_u3980_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    .INIT(16'h88c0))
    _al_u3981 (
    .a(\u2_Display/n4550 ),
    .b(on_off_pad[2]),
    .c(\u2_Display/n4558 [5]),
    .d(\u2_Display/n4556 ),
    .o(_al_u3981_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*~A))"),
    .INIT(16'hc8cc))
    _al_u3982 (
    .a(_al_u3980_o),
    .b(_al_u3978_o),
    .c(_al_u3981_o),
    .d(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u3983 (
    .a(\u2_Display/n4549 ),
    .b(\u2_Display/n4558 [6]),
    .c(\u2_Display/n4556 ),
    .o(_al_u3983_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3984 (
    .a(\u2_Display/n2303 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [6]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [6]),
    .o(_al_u3984_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h5757535f))
    _al_u3985 (
    .a(\u2_Display/n5672 ),
    .b(on_off_pad[1]),
    .c(on_off_pad[0]),
    .d(\u2_Display/n5681 [6]),
    .e(\u2_Display/n5679 ),
    .o(_al_u3985_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*(~B*~(A)*~(E)+~B*A*~(E)+~(~B)*A*E+~B*A*E)))"),
    .INIT(32'haf0f3f0f))
    _al_u3986 (
    .a(_al_u3983_o),
    .b(_al_u3984_o),
    .c(_al_u3985_o),
    .d(\u2_Display/mux19_b0_sel_is_0_o ),
    .e(on_off_pad[2]),
    .o(\u2_Display/n238 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .INIT(16'haab8))
    _al_u3987 (
    .a(\u2_Display/n5671 ),
    .b(on_off_pad[0]),
    .c(\u2_Display/n5681 [7]),
    .d(\u2_Display/n5679 ),
    .o(_al_u3987_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3988 (
    .a(\u2_Display/n2302 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [7]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [7]),
    .o(_al_u3988_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*~(C)+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(C)+~(~A)*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C)"),
    .INIT(32'h3a3a0afa))
    _al_u3989 (
    .a(_al_u3988_o),
    .b(\u2_Display/n4548 ),
    .c(on_off_pad[2]),
    .d(\u2_Display/n4558 [7]),
    .e(\u2_Display/n4556 ),
    .o(_al_u3989_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u399 (
    .a(\u2_Display/n419 [4]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [4]),
    .o(\u2_Display/n447 ));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u3990 (
    .a(_al_u3989_o),
    .b(_al_u3987_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .INIT(16'haab8))
    _al_u3991 (
    .a(\u2_Display/n5670 ),
    .b(on_off_pad[0]),
    .c(\u2_Display/n5681 [8]),
    .d(\u2_Display/n5679 ),
    .o(_al_u3991_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3992 (
    .a(\u2_Display/n2301 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [8]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [8]),
    .o(_al_u3992_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*~(C)+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(C)+~(~A)*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C)"),
    .INIT(32'h3a3a0afa))
    _al_u3993 (
    .a(_al_u3992_o),
    .b(\u2_Display/n4547 ),
    .c(on_off_pad[2]),
    .d(\u2_Display/n4558 [8]),
    .e(\u2_Display/n4556 ),
    .o(_al_u3993_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u3994 (
    .a(_al_u3993_o),
    .b(_al_u3991_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C)*~((~D*~B))+A*C*~((~D*~B))+~(A)*C*(~D*~B)+A*C*(~D*~B))"),
    .INIT(16'haab8))
    _al_u3995 (
    .a(\u2_Display/n5669 ),
    .b(on_off_pad[0]),
    .c(\u2_Display/n5681 [9]),
    .d(\u2_Display/n5679 ),
    .o(_al_u3995_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(E)*~(B)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*~(B)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*E*B+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*E*B)"),
    .INIT(32'h1103ddcf))
    _al_u3996 (
    .a(\u2_Display/n2300 ),
    .b(\u2_Display/mux5_b0_sel_is_0_o ),
    .c(\u2_Display/n2312 [9]),
    .d(\u2_Display/n2310 ),
    .e(\u2_Display/i [9]),
    .o(_al_u3996_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E))*~(C)+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*~(C)+~(~A)*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C+~A*(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)*C)"),
    .INIT(32'h3a3a0afa))
    _al_u3997 (
    .a(_al_u3996_o),
    .b(\u2_Display/n4546 ),
    .c(on_off_pad[2]),
    .d(\u2_Display/n4558 [9]),
    .e(\u2_Display/n4556 ),
    .o(_al_u3997_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u3998 (
    .a(_al_u3997_o),
    .b(_al_u3995_o),
    .c(\u2_Display/mux19_b0_sel_is_0_o ),
    .o(\u2_Display/n238 [9]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u3999 (
    .a(rst_n_pad),
    .o(\u0_PLL/n0 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u400 (
    .a(\u2_Display/n419 [5]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [5]),
    .o(\u2_Display/n446 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u4000 (
    .a(clk_vga),
    .o(vga_clk_pad));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u4001 (
    .a(\u1_Driver/n4 ),
    .o(vga_hs_pad));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u4002 (
    .a(\u1_Driver/n10 ),
    .o(vga_vs_pad));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u4003 (
    .a(\u2_Display/clk1s ),
    .o(\u2_Display/n36 ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u4004 (
    .a(\u2_Display/i [9]),
    .o(\u2_Display/n140 [0]));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u4005 (
    .a(\u2_Display/j [9]),
    .o(\u2_Display/n99 [0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u401 (
    .a(\u2_Display/n419 [6]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [6]),
    .o(\u2_Display/n445 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u402 (
    .a(\u2_Display/n419 [7]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [7]),
    .o(\u2_Display/n444 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u403 (
    .a(\u2_Display/n419 [8]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [8]),
    .o(\u2_Display/n443 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u404 (
    .a(\u2_Display/n419 [9]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [9]),
    .o(\u2_Display/n442 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u405 (
    .a(\u2_Display/n419 [10]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [10]),
    .o(\u2_Display/n441 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u406 (
    .a(\u2_Display/n419 [11]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [11]),
    .o(\u2_Display/n440 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u407 (
    .a(\u2_Display/n419 [12]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [12]),
    .o(\u2_Display/n439 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u408 (
    .a(\u2_Display/n419 [13]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [13]),
    .o(\u2_Display/n438 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u409 (
    .a(\u2_Display/n419 [14]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [14]),
    .o(\u2_Display/n437 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u410 (
    .a(\u2_Display/n419 [15]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [15]),
    .o(\u2_Display/n436 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u411 (
    .a(\u2_Display/n419 [16]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [16]),
    .o(\u2_Display/n435 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u412 (
    .a(\u2_Display/n419 [17]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [17]),
    .o(\u2_Display/n434 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u413 (
    .a(\u2_Display/n419 [18]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [18]),
    .o(\u2_Display/n433 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u414 (
    .a(\u2_Display/n419 [19]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [19]),
    .o(\u2_Display/n432 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u415 (
    .a(\u2_Display/n419 [20]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [20]),
    .o(\u2_Display/n431 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u416 (
    .a(\u2_Display/n419 [21]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [21]),
    .o(\u2_Display/n430 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u417 (
    .a(\u2_Display/n419 [22]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [22]),
    .o(\u2_Display/n429 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u418 (
    .a(\u2_Display/n419 [23]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [23]),
    .o(\u2_Display/n428 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u419 (
    .a(\u2_Display/n419 [24]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [24]),
    .o(\u2_Display/n427 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u420 (
    .a(\u2_Display/n419 [25]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [25]),
    .o(\u2_Display/n426 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u421 (
    .a(\u2_Display/n419 [26]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [26]),
    .o(\u2_Display/n425 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u422 (
    .a(\u2_Display/n419 [27]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [27]),
    .o(\u2_Display/n424 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u423 (
    .a(\u2_Display/n419 [28]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [28]),
    .o(\u2_Display/n423 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u424 (
    .a(\u2_Display/n419 [29]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [29]),
    .o(\u2_Display/n422 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u425 (
    .a(\u2_Display/n419 [30]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [30]),
    .o(\u2_Display/n421 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u426 (
    .a(\u2_Display/n419 [31]),
    .b(\u2_Display/n417 ),
    .c(\u2_Display/counta [31]),
    .o(\u2_Display/n420 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u427 (
    .a(\u2_Display/n1542 [0]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [0]),
    .o(\u2_Display/n1574 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u428 (
    .a(\u2_Display/n1542 [1]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [1]),
    .o(\u2_Display/n1573 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u429 (
    .a(\u2_Display/n1542 [2]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [2]),
    .o(\u2_Display/n1572 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u430 (
    .a(\u2_Display/n1542 [3]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [3]),
    .o(\u2_Display/n1571 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u431 (
    .a(\u2_Display/n1542 [4]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [4]),
    .o(\u2_Display/n1570 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u432 (
    .a(\u2_Display/n1542 [5]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [5]),
    .o(\u2_Display/n1569 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u433 (
    .a(\u2_Display/n1542 [6]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [6]),
    .o(\u2_Display/n1568 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u434 (
    .a(\u2_Display/n1542 [7]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [7]),
    .o(\u2_Display/n1567 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u435 (
    .a(\u2_Display/n1542 [8]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [8]),
    .o(\u2_Display/n1566 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u436 (
    .a(\u2_Display/n1542 [9]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [9]),
    .o(\u2_Display/n1565 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u437 (
    .a(\u2_Display/n1542 [10]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [10]),
    .o(\u2_Display/n1564 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u438 (
    .a(\u2_Display/n1542 [11]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [11]),
    .o(\u2_Display/n1563 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u439 (
    .a(\u2_Display/n1542 [12]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [12]),
    .o(\u2_Display/n1562 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u440 (
    .a(\u2_Display/n1542 [13]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [13]),
    .o(\u2_Display/n1561 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u441 (
    .a(\u2_Display/n1542 [14]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [14]),
    .o(\u2_Display/n1560 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u442 (
    .a(\u2_Display/n1542 [15]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [15]),
    .o(\u2_Display/n1559 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u443 (
    .a(\u2_Display/n1542 [16]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [16]),
    .o(\u2_Display/n1558 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u444 (
    .a(\u2_Display/n1542 [17]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [17]),
    .o(\u2_Display/n1557 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u445 (
    .a(\u2_Display/n1542 [18]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [18]),
    .o(\u2_Display/n1556 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u446 (
    .a(\u2_Display/n1542 [19]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [19]),
    .o(\u2_Display/n1555 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u447 (
    .a(\u2_Display/n1542 [20]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [20]),
    .o(\u2_Display/n1554 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u448 (
    .a(\u2_Display/n1542 [21]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [21]),
    .o(\u2_Display/n1553 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u449 (
    .a(\u2_Display/n1542 [22]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [22]),
    .o(\u2_Display/n1552 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u450 (
    .a(\u2_Display/n1542 [23]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [23]),
    .o(\u2_Display/n1551 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u451 (
    .a(\u2_Display/n1542 [24]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [24]),
    .o(\u2_Display/n1550 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u452 (
    .a(\u2_Display/n1542 [25]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [25]),
    .o(\u2_Display/n1549 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u453 (
    .a(\u2_Display/n1542 [26]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [26]),
    .o(\u2_Display/n1548 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u454 (
    .a(\u2_Display/n1542 [27]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [27]),
    .o(\u2_Display/n1547 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u455 (
    .a(\u2_Display/n1542 [28]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [28]),
    .o(\u2_Display/n1546 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u456 (
    .a(\u2_Display/n1542 [29]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [29]),
    .o(\u2_Display/n1545 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u457 (
    .a(\u2_Display/n1542 [30]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [30]),
    .o(\u2_Display/n1544 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u458 (
    .a(\u2_Display/n1542 [31]),
    .b(\u2_Display/n1540 ),
    .c(\u2_Display/counta [31]),
    .o(\u2_Display/n1543 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u459 (
    .a(\u2_Display/n2665 [0]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [0]),
    .o(\u2_Display/n2697 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u460 (
    .a(\u2_Display/n2665 [1]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [1]),
    .o(\u2_Display/n2696 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u461 (
    .a(\u2_Display/n2665 [2]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [2]),
    .o(\u2_Display/n2695 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u462 (
    .a(\u2_Display/n2665 [3]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [3]),
    .o(\u2_Display/n2694 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u463 (
    .a(\u2_Display/n2665 [4]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [4]),
    .o(\u2_Display/n2693 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u464 (
    .a(\u2_Display/n2665 [5]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [5]),
    .o(\u2_Display/n2692 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u465 (
    .a(\u2_Display/n2665 [6]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [6]),
    .o(\u2_Display/n2691 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u466 (
    .a(\u2_Display/n2665 [7]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [7]),
    .o(\u2_Display/n2690 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u467 (
    .a(\u2_Display/n2665 [8]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [8]),
    .o(\u2_Display/n2689 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u468 (
    .a(\u2_Display/n2665 [9]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [9]),
    .o(\u2_Display/n2688 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u469 (
    .a(\u2_Display/n2665 [10]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [10]),
    .o(\u2_Display/n2687 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u470 (
    .a(\u2_Display/n2665 [11]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [11]),
    .o(\u2_Display/n2686 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u471 (
    .a(\u2_Display/n2665 [12]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [12]),
    .o(\u2_Display/n2685 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u472 (
    .a(\u2_Display/n2665 [13]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [13]),
    .o(\u2_Display/n2684 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u473 (
    .a(\u2_Display/n2665 [14]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [14]),
    .o(\u2_Display/n2683 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u474 (
    .a(\u2_Display/n2665 [15]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [15]),
    .o(\u2_Display/n2682 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u475 (
    .a(\u2_Display/n2665 [16]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [16]),
    .o(\u2_Display/n2681 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u476 (
    .a(\u2_Display/n2665 [17]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [17]),
    .o(\u2_Display/n2680 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u477 (
    .a(\u2_Display/n2665 [18]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [18]),
    .o(\u2_Display/n2679 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u478 (
    .a(\u2_Display/n2665 [19]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [19]),
    .o(\u2_Display/n2678 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u479 (
    .a(\u2_Display/n2665 [20]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [20]),
    .o(\u2_Display/n2677 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u480 (
    .a(\u2_Display/n2665 [21]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [21]),
    .o(\u2_Display/n2676 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u481 (
    .a(\u2_Display/n2665 [22]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [22]),
    .o(\u2_Display/n2675 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u482 (
    .a(\u2_Display/n2665 [23]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [23]),
    .o(\u2_Display/n2674 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u483 (
    .a(\u2_Display/n2665 [24]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [24]),
    .o(\u2_Display/n2673 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u484 (
    .a(\u2_Display/n2665 [25]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [25]),
    .o(\u2_Display/n2672 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u485 (
    .a(\u2_Display/n2665 [26]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [26]),
    .o(\u2_Display/n2671 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u486 (
    .a(\u2_Display/n2665 [27]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [27]),
    .o(\u2_Display/n2670 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u487 (
    .a(\u2_Display/n2665 [28]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [28]),
    .o(\u2_Display/n2669 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u488 (
    .a(\u2_Display/n2665 [29]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [29]),
    .o(\u2_Display/n2668 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u489 (
    .a(\u2_Display/n2665 [30]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [30]),
    .o(\u2_Display/n2667 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u490 (
    .a(\u2_Display/n2665 [31]),
    .b(\u2_Display/n2663 ),
    .c(\u2_Display/counta [31]),
    .o(\u2_Display/n2666 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u491 (
    .a(vga_de_pad),
    .b(lcd_data[23]),
    .o(vga_b_pad[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u492 (
    .a(\u1_Driver/n14 ),
    .b(\u1_Driver/n15 ),
    .c(\u1_Driver/n17 ),
    .d(\u1_Driver/n18 ),
    .o(\u1_Driver/lcd_request ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u493 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [9]),
    .o(lcd_ypos[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u494 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [8]),
    .o(lcd_ypos[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u495 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [7]),
    .o(lcd_ypos[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u496 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [6]),
    .o(lcd_ypos[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u497 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [5]),
    .o(lcd_ypos[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u498 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [4]),
    .o(lcd_ypos[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u499 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [3]),
    .o(lcd_ypos[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u500 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [2]),
    .o(lcd_ypos[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u501 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [11]),
    .o(lcd_ypos[11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u502 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [10]),
    .o(lcd_ypos[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u503 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [1]),
    .o(lcd_ypos[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u504 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n21 [0]),
    .o(lcd_ypos[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u505 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [9]),
    .o(lcd_xpos[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u506 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [8]),
    .o(lcd_xpos[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u507 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [7]),
    .o(lcd_xpos[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u508 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [6]),
    .o(lcd_xpos[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u509 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [5]),
    .o(lcd_xpos[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u510 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [4]),
    .o(lcd_xpos[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u511 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [3]),
    .o(lcd_xpos[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u512 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [2]),
    .o(lcd_xpos[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u513 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [11]),
    .o(lcd_xpos[11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u514 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [10]),
    .o(lcd_xpos[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u515 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [1]),
    .o(lcd_xpos[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u516 (
    .a(\u1_Driver/lcd_request ),
    .b(\u1_Driver/n20 [0]),
    .o(lcd_xpos[0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u517 (
    .a(\u2_Display/n3820 ),
    .b(\u2_Display/n3823 [0]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3855 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u518 (
    .a(\u2_Display/n3819 ),
    .b(\u2_Display/n3823 [1]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3854 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u519 (
    .a(\u2_Display/n3818 ),
    .b(\u2_Display/n3823 [2]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3853 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u520 (
    .a(\u2_Display/n3817 ),
    .b(\u2_Display/n3823 [3]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3852 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u521 (
    .a(\u2_Display/n3816 ),
    .b(\u2_Display/n3823 [4]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3851 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u522 (
    .a(\u2_Display/n3815 ),
    .b(\u2_Display/n3823 [5]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3850 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u523 (
    .a(\u2_Display/n3814 ),
    .b(\u2_Display/n3823 [6]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3849 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u524 (
    .a(\u2_Display/n3813 ),
    .b(\u2_Display/n3823 [7]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3848 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u525 (
    .a(\u2_Display/n3812 ),
    .b(\u2_Display/n3823 [8]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3847 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u526 (
    .a(\u2_Display/n3811 ),
    .b(\u2_Display/n3823 [9]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3846 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u527 (
    .a(\u2_Display/n3810 ),
    .b(\u2_Display/n3823 [10]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3845 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u528 (
    .a(\u2_Display/n3809 ),
    .b(\u2_Display/n3823 [11]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3844 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u529 (
    .a(\u2_Display/n3808 ),
    .b(\u2_Display/n3823 [12]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3843 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u530 (
    .a(\u2_Display/n3807 ),
    .b(\u2_Display/n3823 [13]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3842 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u531 (
    .a(\u2_Display/n3806 ),
    .b(\u2_Display/n3823 [14]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3841 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u532 (
    .a(\u2_Display/n3805 ),
    .b(\u2_Display/n3823 [15]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3840 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u533 (
    .a(\u2_Display/n3804 ),
    .b(\u2_Display/n3823 [16]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3839 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u534 (
    .a(\u2_Display/n3803 ),
    .b(\u2_Display/n3823 [17]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3838 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u535 (
    .a(\u2_Display/n3802 ),
    .b(\u2_Display/n3823 [18]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3837 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u536 (
    .a(\u2_Display/n3801 ),
    .b(\u2_Display/n3823 [19]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3836 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u537 (
    .a(\u2_Display/n3800 ),
    .b(\u2_Display/n3823 [20]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3835 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u538 (
    .a(\u2_Display/n3799 ),
    .b(\u2_Display/n3823 [21]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3834 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u539 (
    .a(\u2_Display/n3798 ),
    .b(\u2_Display/n3823 [22]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3833 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u540 (
    .a(\u2_Display/n3797 ),
    .b(\u2_Display/n3823 [23]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3832 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u541 (
    .a(\u2_Display/n3796 ),
    .b(\u2_Display/n3823 [24]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3831 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u542 (
    .a(\u2_Display/n3795 ),
    .b(\u2_Display/n3823 [25]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3830 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u543 (
    .a(\u2_Display/n3794 ),
    .b(\u2_Display/n3823 [26]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3829 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u544 (
    .a(\u2_Display/n3793 ),
    .b(\u2_Display/n3823 [27]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3828 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u545 (
    .a(\u2_Display/n3792 ),
    .b(\u2_Display/n3823 [28]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3827 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u546 (
    .a(\u2_Display/n3791 ),
    .b(\u2_Display/n3823 [29]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3826 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u547 (
    .a(\u2_Display/n3790 ),
    .b(\u2_Display/n3823 [30]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3825 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u548 (
    .a(\u2_Display/n3789 ),
    .b(\u2_Display/n3823 [31]),
    .c(\u2_Display/n3821 ),
    .o(\u2_Display/n3824 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u549 (
    .a(\u2_Display/n6101 ),
    .b(\u2_Display/n4946 [0]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6136 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u550 (
    .a(\u2_Display/n6100 ),
    .b(\u2_Display/n4946 [1]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6135 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u551 (
    .a(\u2_Display/n6099 ),
    .b(\u2_Display/n4946 [2]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6134 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u552 (
    .a(\u2_Display/n6098 ),
    .b(\u2_Display/n4946 [3]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6133 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u553 (
    .a(\u2_Display/n6097 ),
    .b(\u2_Display/n4946 [4]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6132 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u554 (
    .a(\u2_Display/n6096 ),
    .b(\u2_Display/n4946 [5]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6131 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u555 (
    .a(\u2_Display/n6095 ),
    .b(\u2_Display/n4946 [6]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6130 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u556 (
    .a(\u2_Display/n6094 ),
    .b(\u2_Display/n4946 [7]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6129 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u557 (
    .a(\u2_Display/n6093 ),
    .b(\u2_Display/n4946 [8]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6128 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u558 (
    .a(\u2_Display/n6092 ),
    .b(\u2_Display/n4946 [9]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6127 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u559 (
    .a(\u2_Display/n6091 ),
    .b(\u2_Display/n4946 [10]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6126 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u560 (
    .a(\u2_Display/n6090 ),
    .b(\u2_Display/n4946 [11]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6125 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u561 (
    .a(\u2_Display/n6089 ),
    .b(\u2_Display/n4946 [12]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6124 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u562 (
    .a(\u2_Display/n6088 ),
    .b(\u2_Display/n4946 [13]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6123 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u563 (
    .a(\u2_Display/n6087 ),
    .b(\u2_Display/n4946 [14]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6122 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u564 (
    .a(\u2_Display/n6086 ),
    .b(\u2_Display/n4946 [15]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6121 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u565 (
    .a(\u2_Display/n6085 ),
    .b(\u2_Display/n4946 [16]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6120 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u566 (
    .a(\u2_Display/n6084 ),
    .b(\u2_Display/n4946 [17]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6119 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u567 (
    .a(\u2_Display/n6083 ),
    .b(\u2_Display/n4946 [18]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6118 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u568 (
    .a(\u2_Display/n6082 ),
    .b(\u2_Display/n4946 [19]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6117 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u569 (
    .a(\u2_Display/n6081 ),
    .b(\u2_Display/n4946 [20]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6116 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u570 (
    .a(\u2_Display/n6080 ),
    .b(\u2_Display/n4946 [21]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6115 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u571 (
    .a(\u2_Display/n6079 ),
    .b(\u2_Display/n4946 [22]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6114 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u572 (
    .a(\u2_Display/n6078 ),
    .b(\u2_Display/n4946 [23]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6113 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u573 (
    .a(\u2_Display/n6077 ),
    .b(\u2_Display/n4946 [24]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6112 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u574 (
    .a(\u2_Display/n6076 ),
    .b(\u2_Display/n4946 [25]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6111 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u575 (
    .a(\u2_Display/n6075 ),
    .b(\u2_Display/n4946 [26]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6110 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u576 (
    .a(\u2_Display/n6074 ),
    .b(\u2_Display/n4946 [27]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6109 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u577 (
    .a(\u2_Display/n6073 ),
    .b(\u2_Display/n4946 [28]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6108 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u578 (
    .a(\u2_Display/n6072 ),
    .b(\u2_Display/n4946 [29]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6107 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u579 (
    .a(\u2_Display/n6071 ),
    .b(\u2_Display/n4946 [30]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6106 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u580 (
    .a(\u2_Display/n6070 ),
    .b(\u2_Display/n4946 [31]),
    .c(\u2_Display/n4944 ),
    .o(\u2_Display/n6105 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u581 (
    .a(\u2_Display/n451 ),
    .b(\u2_Display/n454 [0]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n486 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u582 (
    .a(\u2_Display/n450 ),
    .b(\u2_Display/n454 [1]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n485 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u583 (
    .a(\u2_Display/n449 ),
    .b(\u2_Display/n454 [2]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n484 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u584 (
    .a(\u2_Display/n448 ),
    .b(\u2_Display/n454 [3]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n483 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u585 (
    .a(\u2_Display/n447 ),
    .b(\u2_Display/n454 [4]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n482 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u586 (
    .a(\u2_Display/n446 ),
    .b(\u2_Display/n454 [5]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n481 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u587 (
    .a(\u2_Display/n445 ),
    .b(\u2_Display/n454 [6]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n480 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u588 (
    .a(\u2_Display/n444 ),
    .b(\u2_Display/n454 [7]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n479 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u589 (
    .a(\u2_Display/n443 ),
    .b(\u2_Display/n454 [8]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n478 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u590 (
    .a(\u2_Display/n442 ),
    .b(\u2_Display/n454 [9]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n477 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u591 (
    .a(\u2_Display/n441 ),
    .b(\u2_Display/n454 [10]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n476 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u592 (
    .a(\u2_Display/n440 ),
    .b(\u2_Display/n454 [11]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n475 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u593 (
    .a(\u2_Display/n439 ),
    .b(\u2_Display/n454 [12]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n474 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u594 (
    .a(\u2_Display/n438 ),
    .b(\u2_Display/n454 [13]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n473 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u595 (
    .a(\u2_Display/n437 ),
    .b(\u2_Display/n454 [14]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n472 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u596 (
    .a(\u2_Display/n436 ),
    .b(\u2_Display/n454 [15]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n471 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u597 (
    .a(\u2_Display/n435 ),
    .b(\u2_Display/n454 [16]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n470 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u598 (
    .a(\u2_Display/n434 ),
    .b(\u2_Display/n454 [17]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n469 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u599 (
    .a(\u2_Display/n433 ),
    .b(\u2_Display/n454 [18]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n468 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u600 (
    .a(\u2_Display/n432 ),
    .b(\u2_Display/n454 [19]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n467 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u601 (
    .a(\u2_Display/n431 ),
    .b(\u2_Display/n454 [20]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n466 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u602 (
    .a(\u2_Display/n430 ),
    .b(\u2_Display/n454 [21]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n465 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u603 (
    .a(\u2_Display/n429 ),
    .b(\u2_Display/n454 [22]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n464 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u604 (
    .a(\u2_Display/n428 ),
    .b(\u2_Display/n454 [23]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n463 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u605 (
    .a(\u2_Display/n427 ),
    .b(\u2_Display/n454 [24]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n462 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u606 (
    .a(\u2_Display/n426 ),
    .b(\u2_Display/n454 [25]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n461 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u607 (
    .a(\u2_Display/n425 ),
    .b(\u2_Display/n454 [26]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n460 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u608 (
    .a(\u2_Display/n424 ),
    .b(\u2_Display/n454 [27]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n459 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u609 (
    .a(\u2_Display/n423 ),
    .b(\u2_Display/n454 [28]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n458 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u610 (
    .a(\u2_Display/n422 ),
    .b(\u2_Display/n454 [29]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n457 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u611 (
    .a(\u2_Display/n421 ),
    .b(\u2_Display/n454 [30]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n456 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u612 (
    .a(\u2_Display/n420 ),
    .b(\u2_Display/n454 [31]),
    .c(\u2_Display/n452 ),
    .o(\u2_Display/n455 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u613 (
    .a(\u2_Display/n1574 ),
    .b(\u2_Display/n1577 [0]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1609 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u614 (
    .a(\u2_Display/n1573 ),
    .b(\u2_Display/n1577 [1]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1608 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u615 (
    .a(\u2_Display/n1572 ),
    .b(\u2_Display/n1577 [2]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1607 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u616 (
    .a(\u2_Display/n1571 ),
    .b(\u2_Display/n1577 [3]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1606 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u617 (
    .a(\u2_Display/n1570 ),
    .b(\u2_Display/n1577 [4]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1605 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u618 (
    .a(\u2_Display/n1569 ),
    .b(\u2_Display/n1577 [5]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1604 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u619 (
    .a(\u2_Display/n1568 ),
    .b(\u2_Display/n1577 [6]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1603 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u620 (
    .a(\u2_Display/n1567 ),
    .b(\u2_Display/n1577 [7]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1602 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u621 (
    .a(\u2_Display/n1566 ),
    .b(\u2_Display/n1577 [8]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1601 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u622 (
    .a(\u2_Display/n1565 ),
    .b(\u2_Display/n1577 [9]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1600 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u623 (
    .a(\u2_Display/n1564 ),
    .b(\u2_Display/n1577 [10]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1599 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u624 (
    .a(\u2_Display/n1563 ),
    .b(\u2_Display/n1577 [11]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1598 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u625 (
    .a(\u2_Display/n1562 ),
    .b(\u2_Display/n1577 [12]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1597 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u626 (
    .a(\u2_Display/n1561 ),
    .b(\u2_Display/n1577 [13]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1596 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u627 (
    .a(\u2_Display/n1560 ),
    .b(\u2_Display/n1577 [14]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1595 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u628 (
    .a(\u2_Display/n1559 ),
    .b(\u2_Display/n1577 [15]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1594 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u629 (
    .a(\u2_Display/n1558 ),
    .b(\u2_Display/n1577 [16]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1593 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u630 (
    .a(\u2_Display/n1557 ),
    .b(\u2_Display/n1577 [17]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1592 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u631 (
    .a(\u2_Display/n1556 ),
    .b(\u2_Display/n1577 [18]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1591 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u632 (
    .a(\u2_Display/n1555 ),
    .b(\u2_Display/n1577 [19]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1590 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u633 (
    .a(\u2_Display/n1554 ),
    .b(\u2_Display/n1577 [20]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1589 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u634 (
    .a(\u2_Display/n1553 ),
    .b(\u2_Display/n1577 [21]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1588 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u635 (
    .a(\u2_Display/n1552 ),
    .b(\u2_Display/n1577 [22]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1587 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u636 (
    .a(\u2_Display/n1551 ),
    .b(\u2_Display/n1577 [23]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1586 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u637 (
    .a(\u2_Display/n1550 ),
    .b(\u2_Display/n1577 [24]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1585 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u638 (
    .a(\u2_Display/n1549 ),
    .b(\u2_Display/n1577 [25]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1584 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u639 (
    .a(\u2_Display/n1548 ),
    .b(\u2_Display/n1577 [26]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1583 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u640 (
    .a(\u2_Display/n1547 ),
    .b(\u2_Display/n1577 [27]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1582 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u641 (
    .a(\u2_Display/n1546 ),
    .b(\u2_Display/n1577 [28]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1581 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u642 (
    .a(\u2_Display/n1545 ),
    .b(\u2_Display/n1577 [29]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1580 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u643 (
    .a(\u2_Display/n1544 ),
    .b(\u2_Display/n1577 [30]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1579 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u644 (
    .a(\u2_Display/n1543 ),
    .b(\u2_Display/n1577 [31]),
    .c(\u2_Display/n1575 ),
    .o(\u2_Display/n1578 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u645 (
    .a(\u2_Display/n2697 ),
    .b(\u2_Display/n2700 [0]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2732 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u646 (
    .a(\u2_Display/n2696 ),
    .b(\u2_Display/n2700 [1]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2731 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u647 (
    .a(\u2_Display/n2695 ),
    .b(\u2_Display/n2700 [2]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2730 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u648 (
    .a(\u2_Display/n2694 ),
    .b(\u2_Display/n2700 [3]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2729 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u649 (
    .a(\u2_Display/n2693 ),
    .b(\u2_Display/n2700 [4]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2728 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u650 (
    .a(\u2_Display/n2692 ),
    .b(\u2_Display/n2700 [5]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2727 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u651 (
    .a(\u2_Display/n2691 ),
    .b(\u2_Display/n2700 [6]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2726 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u652 (
    .a(\u2_Display/n2690 ),
    .b(\u2_Display/n2700 [7]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2725 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u653 (
    .a(\u2_Display/n2689 ),
    .b(\u2_Display/n2700 [8]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2724 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u654 (
    .a(\u2_Display/n2688 ),
    .b(\u2_Display/n2700 [9]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2723 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u655 (
    .a(\u2_Display/n2687 ),
    .b(\u2_Display/n2700 [10]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2722 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u656 (
    .a(\u2_Display/n2686 ),
    .b(\u2_Display/n2700 [11]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2721 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u657 (
    .a(\u2_Display/n2685 ),
    .b(\u2_Display/n2700 [12]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2720 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u658 (
    .a(\u2_Display/n2684 ),
    .b(\u2_Display/n2700 [13]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2719 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u659 (
    .a(\u2_Display/n2683 ),
    .b(\u2_Display/n2700 [14]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2718 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u660 (
    .a(\u2_Display/n2682 ),
    .b(\u2_Display/n2700 [15]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2717 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u661 (
    .a(\u2_Display/n2681 ),
    .b(\u2_Display/n2700 [16]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2716 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u662 (
    .a(\u2_Display/n2680 ),
    .b(\u2_Display/n2700 [17]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2715 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u663 (
    .a(\u2_Display/n2679 ),
    .b(\u2_Display/n2700 [18]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2714 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u664 (
    .a(\u2_Display/n2678 ),
    .b(\u2_Display/n2700 [19]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2713 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u665 (
    .a(\u2_Display/n2677 ),
    .b(\u2_Display/n2700 [20]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2712 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u666 (
    .a(\u2_Display/n2676 ),
    .b(\u2_Display/n2700 [21]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2711 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u667 (
    .a(\u2_Display/n2675 ),
    .b(\u2_Display/n2700 [22]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2710 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u668 (
    .a(\u2_Display/n2674 ),
    .b(\u2_Display/n2700 [23]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2709 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u669 (
    .a(\u2_Display/n2673 ),
    .b(\u2_Display/n2700 [24]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2708 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u670 (
    .a(\u2_Display/n2672 ),
    .b(\u2_Display/n2700 [25]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2707 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u671 (
    .a(\u2_Display/n2671 ),
    .b(\u2_Display/n2700 [26]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2706 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u672 (
    .a(\u2_Display/n2670 ),
    .b(\u2_Display/n2700 [27]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2705 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u673 (
    .a(\u2_Display/n2669 ),
    .b(\u2_Display/n2700 [28]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2704 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u674 (
    .a(\u2_Display/n2668 ),
    .b(\u2_Display/n2700 [29]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2703 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u675 (
    .a(\u2_Display/n2667 ),
    .b(\u2_Display/n2700 [30]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2702 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u676 (
    .a(\u2_Display/n2666 ),
    .b(\u2_Display/n2700 [31]),
    .c(\u2_Display/n2698 ),
    .o(\u2_Display/n2701 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u677 (
    .a(\u2_Display/n3855 ),
    .b(\u2_Display/n3858 [0]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3890 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u678 (
    .a(\u2_Display/n3854 ),
    .b(\u2_Display/n3858 [1]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3889 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u679 (
    .a(\u2_Display/n3853 ),
    .b(\u2_Display/n3858 [2]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3888 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u680 (
    .a(\u2_Display/n3852 ),
    .b(\u2_Display/n3858 [3]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3887 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u681 (
    .a(\u2_Display/n3851 ),
    .b(\u2_Display/n3858 [4]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3886 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u682 (
    .a(\u2_Display/n3850 ),
    .b(\u2_Display/n3858 [5]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3885 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u683 (
    .a(\u2_Display/n3849 ),
    .b(\u2_Display/n3858 [6]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3884 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u684 (
    .a(\u2_Display/n3848 ),
    .b(\u2_Display/n3858 [7]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3883 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u685 (
    .a(\u2_Display/n3847 ),
    .b(\u2_Display/n3858 [8]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3882 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u686 (
    .a(\u2_Display/n3846 ),
    .b(\u2_Display/n3858 [9]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3881 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u687 (
    .a(\u2_Display/n3845 ),
    .b(\u2_Display/n3858 [10]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3880 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u688 (
    .a(\u2_Display/n3844 ),
    .b(\u2_Display/n3858 [11]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3879 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u689 (
    .a(\u2_Display/n3843 ),
    .b(\u2_Display/n3858 [12]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3878 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u690 (
    .a(\u2_Display/n3842 ),
    .b(\u2_Display/n3858 [13]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3877 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u691 (
    .a(\u2_Display/n3841 ),
    .b(\u2_Display/n3858 [14]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3876 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u692 (
    .a(\u2_Display/n3840 ),
    .b(\u2_Display/n3858 [15]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3875 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u693 (
    .a(\u2_Display/n3839 ),
    .b(\u2_Display/n3858 [16]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3874 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u694 (
    .a(\u2_Display/n3838 ),
    .b(\u2_Display/n3858 [17]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3873 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u695 (
    .a(\u2_Display/n3837 ),
    .b(\u2_Display/n3858 [18]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3872 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u696 (
    .a(\u2_Display/n3836 ),
    .b(\u2_Display/n3858 [19]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3871 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u697 (
    .a(\u2_Display/n3835 ),
    .b(\u2_Display/n3858 [20]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3870 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u698 (
    .a(\u2_Display/n3834 ),
    .b(\u2_Display/n3858 [21]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3869 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u699 (
    .a(\u2_Display/n3833 ),
    .b(\u2_Display/n3858 [22]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3868 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u700 (
    .a(\u2_Display/n3832 ),
    .b(\u2_Display/n3858 [23]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3867 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u701 (
    .a(\u2_Display/n3831 ),
    .b(\u2_Display/n3858 [24]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3866 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u702 (
    .a(\u2_Display/n3830 ),
    .b(\u2_Display/n3858 [25]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3865 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u703 (
    .a(\u2_Display/n3829 ),
    .b(\u2_Display/n3858 [26]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3864 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u704 (
    .a(\u2_Display/n3828 ),
    .b(\u2_Display/n3858 [27]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3863 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u705 (
    .a(\u2_Display/n3827 ),
    .b(\u2_Display/n3858 [28]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3862 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u706 (
    .a(\u2_Display/n3826 ),
    .b(\u2_Display/n3858 [29]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3861 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u707 (
    .a(\u2_Display/n3825 ),
    .b(\u2_Display/n3858 [30]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3860 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u708 (
    .a(\u2_Display/n3824 ),
    .b(\u2_Display/n3858 [31]),
    .c(\u2_Display/n3856 ),
    .o(\u2_Display/n3859 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u709 (
    .a(\u2_Display/n6136 ),
    .b(\u2_Display/n4981 [0]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6171 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u710 (
    .a(\u2_Display/n6135 ),
    .b(\u2_Display/n4981 [1]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6170 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u711 (
    .a(\u2_Display/n6134 ),
    .b(\u2_Display/n4981 [2]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6169 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u712 (
    .a(\u2_Display/n6133 ),
    .b(\u2_Display/n4981 [3]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6168 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u713 (
    .a(\u2_Display/n6132 ),
    .b(\u2_Display/n4981 [4]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6167 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u714 (
    .a(\u2_Display/n6131 ),
    .b(\u2_Display/n4981 [5]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6166 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u715 (
    .a(\u2_Display/n6130 ),
    .b(\u2_Display/n4981 [6]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6165 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u716 (
    .a(\u2_Display/n6129 ),
    .b(\u2_Display/n4981 [7]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6164 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u717 (
    .a(\u2_Display/n6128 ),
    .b(\u2_Display/n4981 [8]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6163 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u718 (
    .a(\u2_Display/n6127 ),
    .b(\u2_Display/n4981 [9]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6162 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u719 (
    .a(\u2_Display/n6126 ),
    .b(\u2_Display/n4981 [10]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6161 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u720 (
    .a(\u2_Display/n6125 ),
    .b(\u2_Display/n4981 [11]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6160 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u721 (
    .a(\u2_Display/n6124 ),
    .b(\u2_Display/n4981 [12]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6159 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u722 (
    .a(\u2_Display/n6123 ),
    .b(\u2_Display/n4981 [13]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6158 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u723 (
    .a(\u2_Display/n6122 ),
    .b(\u2_Display/n4981 [14]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6157 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u724 (
    .a(\u2_Display/n6121 ),
    .b(\u2_Display/n4981 [15]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6156 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u725 (
    .a(\u2_Display/n6120 ),
    .b(\u2_Display/n4981 [16]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6155 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u726 (
    .a(\u2_Display/n6119 ),
    .b(\u2_Display/n4981 [17]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6154 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u727 (
    .a(\u2_Display/n6118 ),
    .b(\u2_Display/n4981 [18]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6153 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u728 (
    .a(\u2_Display/n6117 ),
    .b(\u2_Display/n4981 [19]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6152 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u729 (
    .a(\u2_Display/n6116 ),
    .b(\u2_Display/n4981 [20]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6151 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u730 (
    .a(\u2_Display/n6115 ),
    .b(\u2_Display/n4981 [21]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6150 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u731 (
    .a(\u2_Display/n6114 ),
    .b(\u2_Display/n4981 [22]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6149 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u732 (
    .a(\u2_Display/n6113 ),
    .b(\u2_Display/n4981 [23]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6148 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u733 (
    .a(\u2_Display/n6112 ),
    .b(\u2_Display/n4981 [24]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6147 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u734 (
    .a(\u2_Display/n6111 ),
    .b(\u2_Display/n4981 [25]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6146 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u735 (
    .a(\u2_Display/n6110 ),
    .b(\u2_Display/n4981 [26]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6145 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u736 (
    .a(\u2_Display/n6109 ),
    .b(\u2_Display/n4981 [27]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6144 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u737 (
    .a(\u2_Display/n6108 ),
    .b(\u2_Display/n4981 [28]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6143 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u738 (
    .a(\u2_Display/n6107 ),
    .b(\u2_Display/n4981 [29]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6142 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u739 (
    .a(\u2_Display/n6106 ),
    .b(\u2_Display/n4981 [30]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6141 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u740 (
    .a(\u2_Display/n6105 ),
    .b(\u2_Display/n4981 [31]),
    .c(\u2_Display/n4979 ),
    .o(\u2_Display/n6140 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u741 (
    .a(\u2_Display/n486 ),
    .b(\u2_Display/n489 [0]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n521 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u742 (
    .a(\u2_Display/n485 ),
    .b(\u2_Display/n489 [1]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n520 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u743 (
    .a(\u2_Display/n484 ),
    .b(\u2_Display/n489 [2]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n519 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u744 (
    .a(\u2_Display/n483 ),
    .b(\u2_Display/n489 [3]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n518 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u745 (
    .a(\u2_Display/n482 ),
    .b(\u2_Display/n489 [4]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n517 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u746 (
    .a(\u2_Display/n481 ),
    .b(\u2_Display/n489 [5]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n516 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u747 (
    .a(\u2_Display/n480 ),
    .b(\u2_Display/n489 [6]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n515 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u748 (
    .a(\u2_Display/n479 ),
    .b(\u2_Display/n489 [7]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n514 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u749 (
    .a(\u2_Display/n478 ),
    .b(\u2_Display/n489 [8]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n513 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u750 (
    .a(\u2_Display/n477 ),
    .b(\u2_Display/n489 [9]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n512 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u751 (
    .a(\u2_Display/n476 ),
    .b(\u2_Display/n489 [10]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n511 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u752 (
    .a(\u2_Display/n475 ),
    .b(\u2_Display/n489 [11]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n510 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u753 (
    .a(\u2_Display/n474 ),
    .b(\u2_Display/n489 [12]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n509 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u754 (
    .a(\u2_Display/n473 ),
    .b(\u2_Display/n489 [13]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n508 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u755 (
    .a(\u2_Display/n472 ),
    .b(\u2_Display/n489 [14]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n507 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u756 (
    .a(\u2_Display/n471 ),
    .b(\u2_Display/n489 [15]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n506 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u757 (
    .a(\u2_Display/n470 ),
    .b(\u2_Display/n489 [16]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n505 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u758 (
    .a(\u2_Display/n469 ),
    .b(\u2_Display/n489 [17]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n504 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u759 (
    .a(\u2_Display/n468 ),
    .b(\u2_Display/n489 [18]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n503 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u760 (
    .a(\u2_Display/n467 ),
    .b(\u2_Display/n489 [19]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n502 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u761 (
    .a(\u2_Display/n466 ),
    .b(\u2_Display/n489 [20]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n501 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u762 (
    .a(\u2_Display/n465 ),
    .b(\u2_Display/n489 [21]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n500 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u763 (
    .a(\u2_Display/n464 ),
    .b(\u2_Display/n489 [22]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n499 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u764 (
    .a(\u2_Display/n463 ),
    .b(\u2_Display/n489 [23]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n498 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u765 (
    .a(\u2_Display/n462 ),
    .b(\u2_Display/n489 [24]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n497 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u766 (
    .a(\u2_Display/n461 ),
    .b(\u2_Display/n489 [25]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n496 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u767 (
    .a(\u2_Display/n460 ),
    .b(\u2_Display/n489 [26]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n495 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u768 (
    .a(\u2_Display/n459 ),
    .b(\u2_Display/n489 [27]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n494 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u769 (
    .a(\u2_Display/n458 ),
    .b(\u2_Display/n489 [28]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n493 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u770 (
    .a(\u2_Display/n457 ),
    .b(\u2_Display/n489 [29]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n492 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u771 (
    .a(\u2_Display/n456 ),
    .b(\u2_Display/n489 [30]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n491 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u772 (
    .a(\u2_Display/n455 ),
    .b(\u2_Display/n489 [31]),
    .c(\u2_Display/n487 ),
    .o(\u2_Display/n490 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u773 (
    .a(\u2_Display/n1609 ),
    .b(\u2_Display/n1612 [0]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1644 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u774 (
    .a(\u2_Display/n1608 ),
    .b(\u2_Display/n1612 [1]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1643 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u775 (
    .a(\u2_Display/n1607 ),
    .b(\u2_Display/n1612 [2]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1642 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u776 (
    .a(\u2_Display/n1606 ),
    .b(\u2_Display/n1612 [3]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1641 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u777 (
    .a(\u2_Display/n1605 ),
    .b(\u2_Display/n1612 [4]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1640 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u778 (
    .a(\u2_Display/n1604 ),
    .b(\u2_Display/n1612 [5]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1639 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u779 (
    .a(\u2_Display/n1603 ),
    .b(\u2_Display/n1612 [6]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1638 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u780 (
    .a(\u2_Display/n1602 ),
    .b(\u2_Display/n1612 [7]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1637 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u781 (
    .a(\u2_Display/n1601 ),
    .b(\u2_Display/n1612 [8]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1636 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u782 (
    .a(\u2_Display/n1600 ),
    .b(\u2_Display/n1612 [9]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1635 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u783 (
    .a(\u2_Display/n1599 ),
    .b(\u2_Display/n1612 [10]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1634 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u784 (
    .a(\u2_Display/n1598 ),
    .b(\u2_Display/n1612 [11]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1633 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u785 (
    .a(\u2_Display/n1597 ),
    .b(\u2_Display/n1612 [12]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1632 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u786 (
    .a(\u2_Display/n1596 ),
    .b(\u2_Display/n1612 [13]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1631 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u787 (
    .a(\u2_Display/n1595 ),
    .b(\u2_Display/n1612 [14]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1630 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u788 (
    .a(\u2_Display/n1594 ),
    .b(\u2_Display/n1612 [15]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1629 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u789 (
    .a(\u2_Display/n1593 ),
    .b(\u2_Display/n1612 [16]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1628 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u790 (
    .a(\u2_Display/n1592 ),
    .b(\u2_Display/n1612 [17]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1627 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u791 (
    .a(\u2_Display/n1591 ),
    .b(\u2_Display/n1612 [18]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1626 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u792 (
    .a(\u2_Display/n1590 ),
    .b(\u2_Display/n1612 [19]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1625 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u793 (
    .a(\u2_Display/n1589 ),
    .b(\u2_Display/n1612 [20]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1624 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u794 (
    .a(\u2_Display/n1588 ),
    .b(\u2_Display/n1612 [21]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1623 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u795 (
    .a(\u2_Display/n1587 ),
    .b(\u2_Display/n1612 [22]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1622 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u796 (
    .a(\u2_Display/n1586 ),
    .b(\u2_Display/n1612 [23]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1621 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u797 (
    .a(\u2_Display/n1585 ),
    .b(\u2_Display/n1612 [24]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1620 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u798 (
    .a(\u2_Display/n1584 ),
    .b(\u2_Display/n1612 [25]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1619 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u799 (
    .a(\u2_Display/n1583 ),
    .b(\u2_Display/n1612 [26]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1618 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u800 (
    .a(\u2_Display/n1582 ),
    .b(\u2_Display/n1612 [27]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1617 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u801 (
    .a(\u2_Display/n1581 ),
    .b(\u2_Display/n1612 [28]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1616 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u802 (
    .a(\u2_Display/n1580 ),
    .b(\u2_Display/n1612 [29]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1615 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u803 (
    .a(\u2_Display/n1579 ),
    .b(\u2_Display/n1612 [30]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1614 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u804 (
    .a(\u2_Display/n1578 ),
    .b(\u2_Display/n1612 [31]),
    .c(\u2_Display/n1610 ),
    .o(\u2_Display/n1613 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u805 (
    .a(\u2_Display/n2732 ),
    .b(\u2_Display/n2735 [0]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2767 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u806 (
    .a(\u2_Display/n2731 ),
    .b(\u2_Display/n2735 [1]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2766 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u807 (
    .a(\u2_Display/n2730 ),
    .b(\u2_Display/n2735 [2]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2765 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u808 (
    .a(\u2_Display/n2729 ),
    .b(\u2_Display/n2735 [3]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2764 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u809 (
    .a(\u2_Display/n2728 ),
    .b(\u2_Display/n2735 [4]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2763 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u810 (
    .a(\u2_Display/n2727 ),
    .b(\u2_Display/n2735 [5]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2762 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u811 (
    .a(\u2_Display/n2726 ),
    .b(\u2_Display/n2735 [6]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2761 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u812 (
    .a(\u2_Display/n2725 ),
    .b(\u2_Display/n2735 [7]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2760 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u813 (
    .a(\u2_Display/n2724 ),
    .b(\u2_Display/n2735 [8]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2759 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u814 (
    .a(\u2_Display/n2723 ),
    .b(\u2_Display/n2735 [9]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2758 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u815 (
    .a(\u2_Display/n2722 ),
    .b(\u2_Display/n2735 [10]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2757 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u816 (
    .a(\u2_Display/n2721 ),
    .b(\u2_Display/n2735 [11]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2756 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u817 (
    .a(\u2_Display/n2720 ),
    .b(\u2_Display/n2735 [12]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2755 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u818 (
    .a(\u2_Display/n2719 ),
    .b(\u2_Display/n2735 [13]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2754 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u819 (
    .a(\u2_Display/n2718 ),
    .b(\u2_Display/n2735 [14]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2753 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u820 (
    .a(\u2_Display/n2717 ),
    .b(\u2_Display/n2735 [15]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2752 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u821 (
    .a(\u2_Display/n2716 ),
    .b(\u2_Display/n2735 [16]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2751 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u822 (
    .a(\u2_Display/n2715 ),
    .b(\u2_Display/n2735 [17]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2750 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u823 (
    .a(\u2_Display/n2714 ),
    .b(\u2_Display/n2735 [18]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2749 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u824 (
    .a(\u2_Display/n2713 ),
    .b(\u2_Display/n2735 [19]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2748 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u825 (
    .a(\u2_Display/n2712 ),
    .b(\u2_Display/n2735 [20]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2747 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u826 (
    .a(\u2_Display/n2711 ),
    .b(\u2_Display/n2735 [21]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2746 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u827 (
    .a(\u2_Display/n2710 ),
    .b(\u2_Display/n2735 [22]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2745 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u828 (
    .a(\u2_Display/n2709 ),
    .b(\u2_Display/n2735 [23]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2744 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u829 (
    .a(\u2_Display/n2708 ),
    .b(\u2_Display/n2735 [24]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2743 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u830 (
    .a(\u2_Display/n2707 ),
    .b(\u2_Display/n2735 [25]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2742 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u831 (
    .a(\u2_Display/n2706 ),
    .b(\u2_Display/n2735 [26]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2741 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u832 (
    .a(\u2_Display/n2705 ),
    .b(\u2_Display/n2735 [27]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2740 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u833 (
    .a(\u2_Display/n2704 ),
    .b(\u2_Display/n2735 [28]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2739 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u834 (
    .a(\u2_Display/n2703 ),
    .b(\u2_Display/n2735 [29]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2738 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u835 (
    .a(\u2_Display/n2702 ),
    .b(\u2_Display/n2735 [30]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2737 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u836 (
    .a(\u2_Display/n2701 ),
    .b(\u2_Display/n2735 [31]),
    .c(\u2_Display/n2733 ),
    .o(\u2_Display/n2736 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u837 (
    .a(\u2_Display/n3890 ),
    .b(\u2_Display/n3893 [0]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3925 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u838 (
    .a(\u2_Display/n3889 ),
    .b(\u2_Display/n3893 [1]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3924 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u839 (
    .a(\u2_Display/n3888 ),
    .b(\u2_Display/n3893 [2]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3923 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u840 (
    .a(\u2_Display/n3887 ),
    .b(\u2_Display/n3893 [3]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3922 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u841 (
    .a(\u2_Display/n3886 ),
    .b(\u2_Display/n3893 [4]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3921 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u842 (
    .a(\u2_Display/n3885 ),
    .b(\u2_Display/n3893 [5]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3920 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u843 (
    .a(\u2_Display/n3884 ),
    .b(\u2_Display/n3893 [6]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3919 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u844 (
    .a(\u2_Display/n3883 ),
    .b(\u2_Display/n3893 [7]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3918 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u845 (
    .a(\u2_Display/n3882 ),
    .b(\u2_Display/n3893 [8]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3917 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u846 (
    .a(\u2_Display/n3881 ),
    .b(\u2_Display/n3893 [9]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3916 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u847 (
    .a(\u2_Display/n3880 ),
    .b(\u2_Display/n3893 [10]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3915 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u848 (
    .a(\u2_Display/n3879 ),
    .b(\u2_Display/n3893 [11]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3914 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u849 (
    .a(\u2_Display/n3878 ),
    .b(\u2_Display/n3893 [12]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3913 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u850 (
    .a(\u2_Display/n3877 ),
    .b(\u2_Display/n3893 [13]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3912 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u851 (
    .a(\u2_Display/n3876 ),
    .b(\u2_Display/n3893 [14]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3911 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u852 (
    .a(\u2_Display/n3875 ),
    .b(\u2_Display/n3893 [15]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3910 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u853 (
    .a(\u2_Display/n3874 ),
    .b(\u2_Display/n3893 [16]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3909 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u854 (
    .a(\u2_Display/n3873 ),
    .b(\u2_Display/n3893 [17]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3908 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u855 (
    .a(\u2_Display/n3872 ),
    .b(\u2_Display/n3893 [18]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3907 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u856 (
    .a(\u2_Display/n3871 ),
    .b(\u2_Display/n3893 [19]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3906 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u857 (
    .a(\u2_Display/n3870 ),
    .b(\u2_Display/n3893 [20]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3905 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u858 (
    .a(\u2_Display/n3869 ),
    .b(\u2_Display/n3893 [21]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3904 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u859 (
    .a(\u2_Display/n3868 ),
    .b(\u2_Display/n3893 [22]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3903 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u860 (
    .a(\u2_Display/n3867 ),
    .b(\u2_Display/n3893 [23]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3902 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u861 (
    .a(\u2_Display/n3866 ),
    .b(\u2_Display/n3893 [24]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3901 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u862 (
    .a(\u2_Display/n3865 ),
    .b(\u2_Display/n3893 [25]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3900 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u863 (
    .a(\u2_Display/n3864 ),
    .b(\u2_Display/n3893 [26]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3899 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u864 (
    .a(\u2_Display/n3863 ),
    .b(\u2_Display/n3893 [27]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3898 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u865 (
    .a(\u2_Display/n3862 ),
    .b(\u2_Display/n3893 [28]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3897 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u866 (
    .a(\u2_Display/n3861 ),
    .b(\u2_Display/n3893 [29]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3896 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u867 (
    .a(\u2_Display/n3860 ),
    .b(\u2_Display/n3893 [30]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3895 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u868 (
    .a(\u2_Display/n3859 ),
    .b(\u2_Display/n3893 [31]),
    .c(\u2_Display/n3891 ),
    .o(\u2_Display/n3894 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u869 (
    .a(\u2_Display/n6171 ),
    .b(\u2_Display/n5016 [0]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6206 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u870 (
    .a(\u2_Display/n6170 ),
    .b(\u2_Display/n5016 [1]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6205 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u871 (
    .a(\u2_Display/n6169 ),
    .b(\u2_Display/n5016 [2]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6204 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u872 (
    .a(\u2_Display/n6168 ),
    .b(\u2_Display/n5016 [3]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6203 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u873 (
    .a(\u2_Display/n6167 ),
    .b(\u2_Display/n5016 [4]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6202 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u874 (
    .a(\u2_Display/n6166 ),
    .b(\u2_Display/n5016 [5]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6201 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u875 (
    .a(\u2_Display/n6165 ),
    .b(\u2_Display/n5016 [6]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6200 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u876 (
    .a(\u2_Display/n6164 ),
    .b(\u2_Display/n5016 [7]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6199 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u877 (
    .a(\u2_Display/n6163 ),
    .b(\u2_Display/n5016 [8]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6198 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u878 (
    .a(\u2_Display/n6162 ),
    .b(\u2_Display/n5016 [9]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6197 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u879 (
    .a(\u2_Display/n6161 ),
    .b(\u2_Display/n5016 [10]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6196 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u880 (
    .a(\u2_Display/n6160 ),
    .b(\u2_Display/n5016 [11]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6195 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u881 (
    .a(\u2_Display/n6159 ),
    .b(\u2_Display/n5016 [12]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6194 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u882 (
    .a(\u2_Display/n6158 ),
    .b(\u2_Display/n5016 [13]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6193 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u883 (
    .a(\u2_Display/n6157 ),
    .b(\u2_Display/n5016 [14]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6192 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u884 (
    .a(\u2_Display/n6156 ),
    .b(\u2_Display/n5016 [15]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6191 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u885 (
    .a(\u2_Display/n6155 ),
    .b(\u2_Display/n5016 [16]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6190 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u886 (
    .a(\u2_Display/n6154 ),
    .b(\u2_Display/n5016 [17]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6189 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u887 (
    .a(\u2_Display/n6153 ),
    .b(\u2_Display/n5016 [18]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6188 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u888 (
    .a(\u2_Display/n6152 ),
    .b(\u2_Display/n5016 [19]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6187 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u889 (
    .a(\u2_Display/n6151 ),
    .b(\u2_Display/n5016 [20]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6186 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u890 (
    .a(\u2_Display/n6150 ),
    .b(\u2_Display/n5016 [21]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6185 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u891 (
    .a(\u2_Display/n6149 ),
    .b(\u2_Display/n5016 [22]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6184 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u892 (
    .a(\u2_Display/n6148 ),
    .b(\u2_Display/n5016 [23]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6183 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u893 (
    .a(\u2_Display/n6147 ),
    .b(\u2_Display/n5016 [24]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6182 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u894 (
    .a(\u2_Display/n6146 ),
    .b(\u2_Display/n5016 [25]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6181 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u895 (
    .a(\u2_Display/n6145 ),
    .b(\u2_Display/n5016 [26]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6180 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u896 (
    .a(\u2_Display/n6144 ),
    .b(\u2_Display/n5016 [27]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6179 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u897 (
    .a(\u2_Display/n6143 ),
    .b(\u2_Display/n5016 [28]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6178 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u898 (
    .a(\u2_Display/n6142 ),
    .b(\u2_Display/n5016 [29]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6177 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u899 (
    .a(\u2_Display/n6141 ),
    .b(\u2_Display/n5016 [30]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6176 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u900 (
    .a(\u2_Display/n6140 ),
    .b(\u2_Display/n5016 [31]),
    .c(\u2_Display/n5014 ),
    .o(\u2_Display/n6175 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u901 (
    .a(\u2_Display/n521 ),
    .b(\u2_Display/n524 [0]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n556 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u902 (
    .a(\u2_Display/n520 ),
    .b(\u2_Display/n524 [1]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n555 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u903 (
    .a(\u2_Display/n519 ),
    .b(\u2_Display/n524 [2]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n554 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u904 (
    .a(\u2_Display/n518 ),
    .b(\u2_Display/n524 [3]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n553 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u905 (
    .a(\u2_Display/n517 ),
    .b(\u2_Display/n524 [4]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n552 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u906 (
    .a(\u2_Display/n516 ),
    .b(\u2_Display/n524 [5]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n551 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u907 (
    .a(\u2_Display/n515 ),
    .b(\u2_Display/n524 [6]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n550 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u908 (
    .a(\u2_Display/n514 ),
    .b(\u2_Display/n524 [7]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n549 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u909 (
    .a(\u2_Display/n513 ),
    .b(\u2_Display/n524 [8]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n548 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u910 (
    .a(\u2_Display/n512 ),
    .b(\u2_Display/n524 [9]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n547 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u911 (
    .a(\u2_Display/n511 ),
    .b(\u2_Display/n524 [10]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n546 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u912 (
    .a(\u2_Display/n510 ),
    .b(\u2_Display/n524 [11]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n545 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u913 (
    .a(\u2_Display/n509 ),
    .b(\u2_Display/n524 [12]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n544 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u914 (
    .a(\u2_Display/n508 ),
    .b(\u2_Display/n524 [13]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n543 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u915 (
    .a(\u2_Display/n507 ),
    .b(\u2_Display/n524 [14]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n542 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u916 (
    .a(\u2_Display/n506 ),
    .b(\u2_Display/n524 [15]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n541 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u917 (
    .a(\u2_Display/n505 ),
    .b(\u2_Display/n524 [16]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n540 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u918 (
    .a(\u2_Display/n504 ),
    .b(\u2_Display/n524 [17]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n539 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u919 (
    .a(\u2_Display/n503 ),
    .b(\u2_Display/n524 [18]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n538 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u920 (
    .a(\u2_Display/n502 ),
    .b(\u2_Display/n524 [19]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n537 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u921 (
    .a(\u2_Display/n501 ),
    .b(\u2_Display/n524 [20]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n536 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u922 (
    .a(\u2_Display/n500 ),
    .b(\u2_Display/n524 [21]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n535 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u923 (
    .a(\u2_Display/n499 ),
    .b(\u2_Display/n524 [22]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n534 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u924 (
    .a(\u2_Display/n498 ),
    .b(\u2_Display/n524 [23]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n533 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u925 (
    .a(\u2_Display/n497 ),
    .b(\u2_Display/n524 [24]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n532 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u926 (
    .a(\u2_Display/n496 ),
    .b(\u2_Display/n524 [25]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n531 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u927 (
    .a(\u2_Display/n495 ),
    .b(\u2_Display/n524 [26]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n530 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u928 (
    .a(\u2_Display/n494 ),
    .b(\u2_Display/n524 [27]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n529 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u929 (
    .a(\u2_Display/n493 ),
    .b(\u2_Display/n524 [28]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n528 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u930 (
    .a(\u2_Display/n492 ),
    .b(\u2_Display/n524 [29]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n527 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u931 (
    .a(\u2_Display/n491 ),
    .b(\u2_Display/n524 [30]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n526 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u932 (
    .a(\u2_Display/n490 ),
    .b(\u2_Display/n524 [31]),
    .c(\u2_Display/n522 ),
    .o(\u2_Display/n525 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u933 (
    .a(\u2_Display/n1644 ),
    .b(\u2_Display/n1647 [0]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1679 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u934 (
    .a(\u2_Display/n1643 ),
    .b(\u2_Display/n1647 [1]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1678 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u935 (
    .a(\u2_Display/n1642 ),
    .b(\u2_Display/n1647 [2]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1677 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u936 (
    .a(\u2_Display/n1641 ),
    .b(\u2_Display/n1647 [3]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1676 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u937 (
    .a(\u2_Display/n1640 ),
    .b(\u2_Display/n1647 [4]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1675 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u938 (
    .a(\u2_Display/n1639 ),
    .b(\u2_Display/n1647 [5]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1674 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u939 (
    .a(\u2_Display/n1638 ),
    .b(\u2_Display/n1647 [6]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1673 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u940 (
    .a(\u2_Display/n1637 ),
    .b(\u2_Display/n1647 [7]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1672 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u941 (
    .a(\u2_Display/n1636 ),
    .b(\u2_Display/n1647 [8]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1671 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u942 (
    .a(\u2_Display/n1635 ),
    .b(\u2_Display/n1647 [9]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1670 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u943 (
    .a(\u2_Display/n1634 ),
    .b(\u2_Display/n1647 [10]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1669 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u944 (
    .a(\u2_Display/n1633 ),
    .b(\u2_Display/n1647 [11]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1668 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u945 (
    .a(\u2_Display/n1632 ),
    .b(\u2_Display/n1647 [12]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1667 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u946 (
    .a(\u2_Display/n1631 ),
    .b(\u2_Display/n1647 [13]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1666 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u947 (
    .a(\u2_Display/n1630 ),
    .b(\u2_Display/n1647 [14]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1665 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u948 (
    .a(\u2_Display/n1629 ),
    .b(\u2_Display/n1647 [15]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1664 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u949 (
    .a(\u2_Display/n1628 ),
    .b(\u2_Display/n1647 [16]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1663 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u950 (
    .a(\u2_Display/n1627 ),
    .b(\u2_Display/n1647 [17]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1662 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u951 (
    .a(\u2_Display/n1626 ),
    .b(\u2_Display/n1647 [18]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1661 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u952 (
    .a(\u2_Display/n1625 ),
    .b(\u2_Display/n1647 [19]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1660 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u953 (
    .a(\u2_Display/n1624 ),
    .b(\u2_Display/n1647 [20]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1659 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u954 (
    .a(\u2_Display/n1623 ),
    .b(\u2_Display/n1647 [21]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1658 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u955 (
    .a(\u2_Display/n1622 ),
    .b(\u2_Display/n1647 [22]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1657 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u956 (
    .a(\u2_Display/n1621 ),
    .b(\u2_Display/n1647 [23]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1656 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u957 (
    .a(\u2_Display/n1620 ),
    .b(\u2_Display/n1647 [24]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1655 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u958 (
    .a(\u2_Display/n1619 ),
    .b(\u2_Display/n1647 [25]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1654 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u959 (
    .a(\u2_Display/n1618 ),
    .b(\u2_Display/n1647 [26]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1653 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u960 (
    .a(\u2_Display/n1617 ),
    .b(\u2_Display/n1647 [27]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1652 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u961 (
    .a(\u2_Display/n1616 ),
    .b(\u2_Display/n1647 [28]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1651 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u962 (
    .a(\u2_Display/n1615 ),
    .b(\u2_Display/n1647 [29]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1650 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u963 (
    .a(\u2_Display/n1614 ),
    .b(\u2_Display/n1647 [30]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1649 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u964 (
    .a(\u2_Display/n1613 ),
    .b(\u2_Display/n1647 [31]),
    .c(\u2_Display/n1645 ),
    .o(\u2_Display/n1648 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u965 (
    .a(\u2_Display/n2767 ),
    .b(\u2_Display/n2770 [0]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2802 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u966 (
    .a(\u2_Display/n2766 ),
    .b(\u2_Display/n2770 [1]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2801 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u967 (
    .a(\u2_Display/n2765 ),
    .b(\u2_Display/n2770 [2]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2800 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u968 (
    .a(\u2_Display/n2764 ),
    .b(\u2_Display/n2770 [3]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2799 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u969 (
    .a(\u2_Display/n2763 ),
    .b(\u2_Display/n2770 [4]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2798 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u970 (
    .a(\u2_Display/n2762 ),
    .b(\u2_Display/n2770 [5]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2797 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u971 (
    .a(\u2_Display/n2761 ),
    .b(\u2_Display/n2770 [6]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2796 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u972 (
    .a(\u2_Display/n2760 ),
    .b(\u2_Display/n2770 [7]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2795 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u973 (
    .a(\u2_Display/n2759 ),
    .b(\u2_Display/n2770 [8]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2794 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u974 (
    .a(\u2_Display/n2758 ),
    .b(\u2_Display/n2770 [9]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2793 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u975 (
    .a(\u2_Display/n2757 ),
    .b(\u2_Display/n2770 [10]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2792 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u976 (
    .a(\u2_Display/n2756 ),
    .b(\u2_Display/n2770 [11]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2791 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u977 (
    .a(\u2_Display/n2755 ),
    .b(\u2_Display/n2770 [12]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2790 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u978 (
    .a(\u2_Display/n2754 ),
    .b(\u2_Display/n2770 [13]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2789 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u979 (
    .a(\u2_Display/n2753 ),
    .b(\u2_Display/n2770 [14]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2788 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u980 (
    .a(\u2_Display/n2752 ),
    .b(\u2_Display/n2770 [15]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2787 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u981 (
    .a(\u2_Display/n2751 ),
    .b(\u2_Display/n2770 [16]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2786 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u982 (
    .a(\u2_Display/n2750 ),
    .b(\u2_Display/n2770 [17]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2785 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u983 (
    .a(\u2_Display/n2749 ),
    .b(\u2_Display/n2770 [18]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2784 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u984 (
    .a(\u2_Display/n2748 ),
    .b(\u2_Display/n2770 [19]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2783 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u985 (
    .a(\u2_Display/n2747 ),
    .b(\u2_Display/n2770 [20]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2782 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u986 (
    .a(\u2_Display/n2746 ),
    .b(\u2_Display/n2770 [21]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2781 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u987 (
    .a(\u2_Display/n2745 ),
    .b(\u2_Display/n2770 [22]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2780 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u988 (
    .a(\u2_Display/n2744 ),
    .b(\u2_Display/n2770 [23]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2779 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u989 (
    .a(\u2_Display/n2743 ),
    .b(\u2_Display/n2770 [24]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2778 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u990 (
    .a(\u2_Display/n2742 ),
    .b(\u2_Display/n2770 [25]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2777 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u991 (
    .a(\u2_Display/n2741 ),
    .b(\u2_Display/n2770 [26]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2776 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u992 (
    .a(\u2_Display/n2740 ),
    .b(\u2_Display/n2770 [27]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2775 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u993 (
    .a(\u2_Display/n2739 ),
    .b(\u2_Display/n2770 [28]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2774 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u994 (
    .a(\u2_Display/n2738 ),
    .b(\u2_Display/n2770 [29]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2773 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u995 (
    .a(\u2_Display/n2737 ),
    .b(\u2_Display/n2770 [30]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2772 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u996 (
    .a(\u2_Display/n2736 ),
    .b(\u2_Display/n2770 [31]),
    .c(\u2_Display/n2768 ),
    .o(\u2_Display/n2771 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u997 (
    .a(\u1_Driver/hcnt [0]),
    .b(\u1_Driver/hcnt [1]),
    .c(\u1_Driver/hcnt [10]),
    .d(\u1_Driver/hcnt [11]),
    .o(_al_u997_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    _al_u998 (
    .a(_al_u997_o),
    .b(\u1_Driver/hcnt [2]),
    .c(\u1_Driver/hcnt [3]),
    .d(\u1_Driver/hcnt [4]),
    .e(\u1_Driver/hcnt [5]),
    .o(_al_u998_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*A)"),
    .INIT(32'h00200000))
    _al_u999 (
    .a(_al_u998_o),
    .b(\u1_Driver/hcnt [6]),
    .c(\u1_Driver/hcnt [7]),
    .d(\u1_Driver/hcnt [8]),
    .e(\u1_Driver/hcnt [9]),
    .o(\u1_Driver/n5 ));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  EG_PHY_GCLK \u0_PLL/uut/bufg_feedback  (
    .clki(\u0_PLL/uut/clk0_buf ),
    .clko(clk_vga));  // al_ip/PLL.v(34)
  EG_PHY_PLL #(
    .CLKC0_CPHASE(8),
    .CLKC0_DIV(9),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(1),
    .CLKC1_DIV(1),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_ENABLE("DISABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(1),
    .CLKC2_DIV(1),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("DISABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(1),
    .CLKC3_DIV(1),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("DISABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(9),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("24.000"),
    .FREQ_LOCK_ACCURACY(2),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .REFCLK_DIV(2),
    .REFCLK_SEL("INTERNAL"),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \u0_PLL/uut/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dwe(1'b0),
    .fbclk(clk_vga),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(clk_24m_pad),
    .reset(\u0_PLL/n0 ),
    .stdby(1'b0),
    .clkc({open_n697,open_n698,open_n699,open_n700,\u0_PLL/uut/clk0_buf }));  // al_ip/PLL.v(57)
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add0/ucin_al_u5013"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add0/u11_al_u5016  (
    .a({open_n711,\u1_Driver/hcnt [11]}),
    .c(2'b00),
    .d({open_n716,1'b0}),
    .fci(\u1_Driver/add0/c11 ),
    .f({open_n733,\u1_Driver/n2 [11]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add0/ucin_al_u5013"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add0/u3_al_u5014  (
    .a({\u1_Driver/hcnt [5],\u1_Driver/hcnt [3]}),
    .b({\u1_Driver/hcnt [6],\u1_Driver/hcnt [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u1_Driver/add0/c3 ),
    .f({\u1_Driver/n2 [5],\u1_Driver/n2 [3]}),
    .fco(\u1_Driver/add0/c7 ),
    .fx({\u1_Driver/n2 [6],\u1_Driver/n2 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add0/ucin_al_u5013"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add0/u7_al_u5015  (
    .a({\u1_Driver/hcnt [9],\u1_Driver/hcnt [7]}),
    .b({\u1_Driver/hcnt [10],\u1_Driver/hcnt [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u1_Driver/add0/c7 ),
    .f({\u1_Driver/n2 [9],\u1_Driver/n2 [7]}),
    .fco(\u1_Driver/add0/c11 ),
    .fx({\u1_Driver/n2 [10],\u1_Driver/n2 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add0/ucin_al_u5013"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add0/ucin_al_u5013  (
    .a({\u1_Driver/hcnt [1],1'b0}),
    .b({\u1_Driver/hcnt [2],\u1_Driver/hcnt [0]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .f({\u1_Driver/n2 [1],open_n792}),
    .fco(\u1_Driver/add0/c3 ),
    .fx({\u1_Driver/n2 [2],\u1_Driver/n2 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add1/ucin_al_u5017"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add1/u11_al_u5020  (
    .a({open_n795,\u1_Driver/vcnt [11]}),
    .c(2'b00),
    .d({open_n800,1'b0}),
    .fci(\u1_Driver/add1/c11 ),
    .f({open_n817,\u1_Driver/n7 [11]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add1/ucin_al_u5017"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add1/u3_al_u5018  (
    .a({\u1_Driver/vcnt [5],\u1_Driver/vcnt [3]}),
    .b({\u1_Driver/vcnt [6],\u1_Driver/vcnt [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u1_Driver/add1/c3 ),
    .f({\u1_Driver/n7 [5],\u1_Driver/n7 [3]}),
    .fco(\u1_Driver/add1/c7 ),
    .fx({\u1_Driver/n7 [6],\u1_Driver/n7 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add1/ucin_al_u5017"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add1/u7_al_u5019  (
    .a({\u1_Driver/vcnt [9],\u1_Driver/vcnt [7]}),
    .b({\u1_Driver/vcnt [10],\u1_Driver/vcnt [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u1_Driver/add1/c7 ),
    .f({\u1_Driver/n7 [9],\u1_Driver/n7 [7]}),
    .fco(\u1_Driver/add1/c11 ),
    .fx({\u1_Driver/n7 [10],\u1_Driver/n7 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/add1/ucin_al_u5017"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/add1/ucin_al_u5017  (
    .a({\u1_Driver/vcnt [1],1'b0}),
    .b({\u1_Driver/vcnt [2],\u1_Driver/vcnt [0]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .f({\u1_Driver/n7 [1],open_n876}),
    .fco(\u1_Driver/add1/c3 ),
    .fx({\u1_Driver/n7 [2],\u1_Driver/n7 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_0|u1_Driver/lt0_cin  (
    .a({\u1_Driver/hcnt [0],1'b0}),
    .b({1'b1,open_n879}),
    .fco(\u1_Driver/lt0_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_10|u1_Driver/lt0_9  (
    .a(\u1_Driver/hcnt [10:9]),
    .b(2'b11),
    .fci(\u1_Driver/lt0_c9 ),
    .fco(\u1_Driver/lt0_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_2|u1_Driver/lt0_1  (
    .a(\u1_Driver/hcnt [2:1]),
    .b(2'b11),
    .fci(\u1_Driver/lt0_c1 ),
    .fco(\u1_Driver/lt0_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_4|u1_Driver/lt0_3  (
    .a(\u1_Driver/hcnt [4:3]),
    .b(2'b10),
    .fci(\u1_Driver/lt0_c3 ),
    .fco(\u1_Driver/lt0_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_6|u1_Driver/lt0_5  (
    .a(\u1_Driver/hcnt [6:5]),
    .b(2'b00),
    .fci(\u1_Driver/lt0_c5 ),
    .fco(\u1_Driver/lt0_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_8|u1_Driver/lt0_7  (
    .a(\u1_Driver/hcnt [8:7]),
    .b(2'b01),
    .fci(\u1_Driver/lt0_c7 ),
    .fco(\u1_Driver/lt0_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt0_0|u1_Driver/lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt0_cout|u1_Driver/lt0_11  (
    .a({1'b0,\u1_Driver/hcnt [11]}),
    .b(2'b10),
    .fci(\u1_Driver/lt0_c11 ),
    .f({\u1_Driver/n1 ,open_n1043}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_0|u1_Driver/lt1_cin  (
    .a({\u1_Driver/hcnt [0],1'b1}),
    .b({1'b1,open_n1049}),
    .fco(\u1_Driver/lt1_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_10|u1_Driver/lt1_9  (
    .a(\u1_Driver/hcnt [10:9]),
    .b(2'b00),
    .fci(\u1_Driver/lt1_c9 ),
    .fco(\u1_Driver/lt1_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_2|u1_Driver/lt1_1  (
    .a(\u1_Driver/hcnt [2:1]),
    .b(2'b11),
    .fci(\u1_Driver/lt1_c1 ),
    .fco(\u1_Driver/lt1_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_4|u1_Driver/lt1_3  (
    .a(\u1_Driver/hcnt [4:3]),
    .b(2'b01),
    .fci(\u1_Driver/lt1_c3 ),
    .fco(\u1_Driver/lt1_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_6|u1_Driver/lt1_5  (
    .a(\u1_Driver/hcnt [6:5]),
    .b(2'b11),
    .fci(\u1_Driver/lt1_c5 ),
    .fco(\u1_Driver/lt1_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_8|u1_Driver/lt1_7  (
    .a(\u1_Driver/hcnt [8:7]),
    .b(2'b00),
    .fci(\u1_Driver/lt1_c7 ),
    .fco(\u1_Driver/lt1_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt1_0|u1_Driver/lt1_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt1_cout|u1_Driver/lt1_11  (
    .a({1'b0,\u1_Driver/hcnt [11]}),
    .b(2'b10),
    .fci(\u1_Driver/lt1_c11 ),
    .f({\u1_Driver/n4 ,open_n1213}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_0|u1_Driver/lt2_cin  (
    .a({\u1_Driver/vcnt [0],1'b1}),
    .b({1'b0,open_n1219}),
    .fco(\u1_Driver/lt2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_10|u1_Driver/lt2_9  (
    .a(\u1_Driver/vcnt [10:9]),
    .b(2'b00),
    .fci(\u1_Driver/lt2_c9 ),
    .fco(\u1_Driver/lt2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_2|u1_Driver/lt2_1  (
    .a(\u1_Driver/vcnt [2:1]),
    .b(2'b01),
    .fci(\u1_Driver/lt2_c1 ),
    .fco(\u1_Driver/lt2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_4|u1_Driver/lt2_3  (
    .a(\u1_Driver/vcnt [4:3]),
    .b(2'b00),
    .fci(\u1_Driver/lt2_c3 ),
    .fco(\u1_Driver/lt2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_6|u1_Driver/lt2_5  (
    .a(\u1_Driver/vcnt [6:5]),
    .b(2'b00),
    .fci(\u1_Driver/lt2_c5 ),
    .fco(\u1_Driver/lt2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_8|u1_Driver/lt2_7  (
    .a(\u1_Driver/vcnt [8:7]),
    .b(2'b00),
    .fci(\u1_Driver/lt2_c7 ),
    .fco(\u1_Driver/lt2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt2_0|u1_Driver/lt2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt2_cout|u1_Driver/lt2_11  (
    .a({1'b0,\u1_Driver/vcnt [11]}),
    .b(2'b10),
    .fci(\u1_Driver/lt2_c11 ),
    .f({\u1_Driver/n10 ,open_n1383}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_0|u1_Driver/lt3_cin  (
    .a(2'b01),
    .b({\u1_Driver/hcnt [0],open_n1389}),
    .fco(\u1_Driver/lt3_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_10|u1_Driver/lt3_9  (
    .a(2'b00),
    .b(\u1_Driver/hcnt [10:9]),
    .fci(\u1_Driver/lt3_c9 ),
    .fco(\u1_Driver/lt3_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_2|u1_Driver/lt3_1  (
    .a(2'b00),
    .b(\u1_Driver/hcnt [2:1]),
    .fci(\u1_Driver/lt3_c1 ),
    .fco(\u1_Driver/lt3_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_4|u1_Driver/lt3_3  (
    .a(2'b01),
    .b(\u1_Driver/hcnt [4:3]),
    .fci(\u1_Driver/lt3_c3 ),
    .fco(\u1_Driver/lt3_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_6|u1_Driver/lt3_5  (
    .a(2'b11),
    .b(\u1_Driver/hcnt [6:5]),
    .fci(\u1_Driver/lt3_c5 ),
    .fco(\u1_Driver/lt3_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_8|u1_Driver/lt3_7  (
    .a(2'b10),
    .b(\u1_Driver/hcnt [8:7]),
    .fci(\u1_Driver/lt3_c7 ),
    .fco(\u1_Driver/lt3_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt3_0|u1_Driver/lt3_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt3_cout|u1_Driver/lt3_11  (
    .a(2'b00),
    .b({1'b1,\u1_Driver/hcnt [11]}),
    .fci(\u1_Driver/lt3_c11 ),
    .f({\u1_Driver/n11 ,open_n1553}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_0|u1_Driver/lt4_cin  (
    .a({\u1_Driver/hcnt [0],1'b0}),
    .b({1'b0,open_n1559}),
    .fco(\u1_Driver/lt4_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_10|u1_Driver/lt4_9  (
    .a(\u1_Driver/hcnt [10:9]),
    .b(2'b11),
    .fci(\u1_Driver/lt4_c9 ),
    .fco(\u1_Driver/lt4_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_2|u1_Driver/lt4_1  (
    .a(\u1_Driver/hcnt [2:1]),
    .b(2'b00),
    .fci(\u1_Driver/lt4_c1 ),
    .fco(\u1_Driver/lt4_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_4|u1_Driver/lt4_3  (
    .a(\u1_Driver/hcnt [4:3]),
    .b(2'b01),
    .fci(\u1_Driver/lt4_c3 ),
    .fco(\u1_Driver/lt4_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_6|u1_Driver/lt4_5  (
    .a(\u1_Driver/hcnt [6:5]),
    .b(2'b11),
    .fci(\u1_Driver/lt4_c5 ),
    .fco(\u1_Driver/lt4_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_8|u1_Driver/lt4_7  (
    .a(\u1_Driver/hcnt [8:7]),
    .b(2'b00),
    .fci(\u1_Driver/lt4_c7 ),
    .fco(\u1_Driver/lt4_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt4_0|u1_Driver/lt4_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt4_cout|u1_Driver/lt4_11  (
    .a({1'b0,\u1_Driver/hcnt [11]}),
    .b(2'b10),
    .fci(\u1_Driver/lt4_c11 ),
    .f({\u1_Driver/n12 ,open_n1723}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_0|u1_Driver/lt5_cin  (
    .a(2'b11),
    .b({\u1_Driver/vcnt [0],open_n1729}),
    .fco(\u1_Driver/lt5_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_10|u1_Driver/lt5_9  (
    .a(2'b00),
    .b(\u1_Driver/vcnt [10:9]),
    .fci(\u1_Driver/lt5_c9 ),
    .fco(\u1_Driver/lt5_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_2|u1_Driver/lt5_1  (
    .a(2'b00),
    .b(\u1_Driver/vcnt [2:1]),
    .fci(\u1_Driver/lt5_c1 ),
    .fco(\u1_Driver/lt5_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_4|u1_Driver/lt5_3  (
    .a(2'b01),
    .b(\u1_Driver/vcnt [4:3]),
    .fci(\u1_Driver/lt5_c3 ),
    .fco(\u1_Driver/lt5_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_6|u1_Driver/lt5_5  (
    .a(2'b01),
    .b(\u1_Driver/vcnt [6:5]),
    .fci(\u1_Driver/lt5_c5 ),
    .fco(\u1_Driver/lt5_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_8|u1_Driver/lt5_7  (
    .a(2'b00),
    .b(\u1_Driver/vcnt [8:7]),
    .fci(\u1_Driver/lt5_c7 ),
    .fco(\u1_Driver/lt5_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt5_0|u1_Driver/lt5_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt5_cout|u1_Driver/lt5_11  (
    .a(2'b00),
    .b({1'b1,\u1_Driver/vcnt [11]}),
    .fci(\u1_Driver/lt5_c11 ),
    .f({\u1_Driver/n14 ,open_n1893}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_0|u1_Driver/lt6_cin  (
    .a({\u1_Driver/vcnt [0],1'b0}),
    .b({1'b1,open_n1899}),
    .fco(\u1_Driver/lt6_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_10|u1_Driver/lt6_9  (
    .a(\u1_Driver/vcnt [10:9]),
    .b(2'b10),
    .fci(\u1_Driver/lt6_c9 ),
    .fco(\u1_Driver/lt6_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_2|u1_Driver/lt6_1  (
    .a(\u1_Driver/vcnt [2:1]),
    .b(2'b00),
    .fci(\u1_Driver/lt6_c1 ),
    .fco(\u1_Driver/lt6_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_4|u1_Driver/lt6_3  (
    .a(\u1_Driver/vcnt [4:3]),
    .b(2'b01),
    .fci(\u1_Driver/lt6_c3 ),
    .fco(\u1_Driver/lt6_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_6|u1_Driver/lt6_5  (
    .a(\u1_Driver/vcnt [6:5]),
    .b(2'b01),
    .fci(\u1_Driver/lt6_c5 ),
    .fco(\u1_Driver/lt6_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_8|u1_Driver/lt6_7  (
    .a(\u1_Driver/vcnt [8:7]),
    .b(2'b00),
    .fci(\u1_Driver/lt6_c7 ),
    .fco(\u1_Driver/lt6_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt6_0|u1_Driver/lt6_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt6_cout|u1_Driver/lt6_11  (
    .a({1'b0,\u1_Driver/vcnt [11]}),
    .b(2'b10),
    .fci(\u1_Driver/lt6_c11 ),
    .f({\u1_Driver/n15 ,open_n2063}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_0|u1_Driver/lt7_cin  (
    .a(2'b11),
    .b({\u1_Driver/hcnt [0],open_n2069}),
    .fco(\u1_Driver/lt7_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_10|u1_Driver/lt7_9  (
    .a(2'b00),
    .b(\u1_Driver/hcnt [10:9]),
    .fci(\u1_Driver/lt7_c9 ),
    .fco(\u1_Driver/lt7_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_2|u1_Driver/lt7_1  (
    .a(2'b11),
    .b(\u1_Driver/hcnt [2:1]),
    .fci(\u1_Driver/lt7_c1 ),
    .fco(\u1_Driver/lt7_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_4|u1_Driver/lt7_3  (
    .a(2'b00),
    .b(\u1_Driver/hcnt [4:3]),
    .fci(\u1_Driver/lt7_c3 ),
    .fco(\u1_Driver/lt7_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_6|u1_Driver/lt7_5  (
    .a(2'b11),
    .b(\u1_Driver/hcnt [6:5]),
    .fci(\u1_Driver/lt7_c5 ),
    .fco(\u1_Driver/lt7_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_8|u1_Driver/lt7_7  (
    .a(2'b10),
    .b(\u1_Driver/hcnt [8:7]),
    .fci(\u1_Driver/lt7_c7 ),
    .fco(\u1_Driver/lt7_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt7_0|u1_Driver/lt7_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt7_cout|u1_Driver/lt7_11  (
    .a(2'b00),
    .b({1'b1,\u1_Driver/hcnt [11]}),
    .fci(\u1_Driver/lt7_c11 ),
    .f({\u1_Driver/n17 ,open_n2233}));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_0|u1_Driver/lt8_cin  (
    .a({\u1_Driver/hcnt [0],1'b0}),
    .b({1'b1,open_n2239}),
    .fco(\u1_Driver/lt8_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_10|u1_Driver/lt8_9  (
    .a(\u1_Driver/hcnt [10:9]),
    .b(2'b11),
    .fci(\u1_Driver/lt8_c9 ),
    .fco(\u1_Driver/lt8_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_2|u1_Driver/lt8_1  (
    .a(\u1_Driver/hcnt [2:1]),
    .b(2'b11),
    .fci(\u1_Driver/lt8_c1 ),
    .fco(\u1_Driver/lt8_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_4|u1_Driver/lt8_3  (
    .a(\u1_Driver/hcnt [4:3]),
    .b(2'b00),
    .fci(\u1_Driver/lt8_c3 ),
    .fco(\u1_Driver/lt8_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_6|u1_Driver/lt8_5  (
    .a(\u1_Driver/hcnt [6:5]),
    .b(2'b11),
    .fci(\u1_Driver/lt8_c5 ),
    .fco(\u1_Driver/lt8_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_8|u1_Driver/lt8_7  (
    .a(\u1_Driver/hcnt [8:7]),
    .b(2'b00),
    .fci(\u1_Driver/lt8_c7 ),
    .fco(\u1_Driver/lt8_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1_Driver/lt8_0|u1_Driver/lt8_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u1_Driver/lt8_cout|u1_Driver/lt8_11  (
    .a({1'b0,\u1_Driver/hcnt [11]}),
    .b(2'b10),
    .fci(\u1_Driver/lt8_c11 ),
    .f({\u1_Driver/n18 ,open_n2403}));
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b0  (
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d(\u1_Driver/n8 [0]),
    .sr(rst_n_pad),
    .q(\u1_Driver/vcnt [0]));  // source/rtl/Driver.v(78)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b1  (
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d(\u1_Driver/n8 [1]),
    .sr(rst_n_pad),
    .q(\u1_Driver/vcnt [1]));  // source/rtl/Driver.v(78)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b10  (
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d(\u1_Driver/n8 [10]),
    .sr(rst_n_pad),
    .q(\u1_Driver/vcnt [10]));  // source/rtl/Driver.v(78)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b11  (
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d(\u1_Driver/n8 [11]),
    .sr(rst_n_pad),
    .q(\u1_Driver/vcnt [11]));  // source/rtl/Driver.v(78)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b2  (
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d(\u1_Driver/n8 [2]),
    .sr(rst_n_pad),
    .q(\u1_Driver/vcnt [2]));  // source/rtl/Driver.v(78)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b3  (
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d(\u1_Driver/n8 [3]),
    .sr(rst_n_pad),
    .q(\u1_Driver/vcnt [3]));  // source/rtl/Driver.v(78)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b4  (
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d(\u1_Driver/n8 [4]),
    .sr(rst_n_pad),
    .q(\u1_Driver/vcnt [4]));  // source/rtl/Driver.v(78)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b5  (
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d(\u1_Driver/n8 [5]),
    .sr(rst_n_pad),
    .q(\u1_Driver/vcnt [5]));  // source/rtl/Driver.v(78)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b6  (
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d(\u1_Driver/n8 [6]),
    .sr(rst_n_pad),
    .q(\u1_Driver/vcnt [6]));  // source/rtl/Driver.v(78)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b7  (
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d(\u1_Driver/n8 [7]),
    .sr(rst_n_pad),
    .q(\u1_Driver/vcnt [7]));  // source/rtl/Driver.v(78)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b8  (
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d(\u1_Driver/n8 [8]),
    .sr(rst_n_pad),
    .q(\u1_Driver/vcnt [8]));  // source/rtl/Driver.v(78)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg0_b9  (
    .ce(\u1_Driver/n5 ),
    .clk(clk_vga),
    .d(\u1_Driver/n8 [9]),
    .sr(rst_n_pad),
    .q(\u1_Driver/vcnt [9]));  // source/rtl/Driver.v(78)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b0  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [0]),
    .sr(rst_n_pad),
    .q(\u1_Driver/hcnt [0]));  // source/rtl/Driver.v(62)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b1  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [1]),
    .sr(rst_n_pad),
    .q(\u1_Driver/hcnt [1]));  // source/rtl/Driver.v(62)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b10  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [10]),
    .sr(rst_n_pad),
    .q(\u1_Driver/hcnt [10]));  // source/rtl/Driver.v(62)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b11  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [11]),
    .sr(rst_n_pad),
    .q(\u1_Driver/hcnt [11]));  // source/rtl/Driver.v(62)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b2  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [2]),
    .sr(rst_n_pad),
    .q(\u1_Driver/hcnt [2]));  // source/rtl/Driver.v(62)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b3  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [3]),
    .sr(rst_n_pad),
    .q(\u1_Driver/hcnt [3]));  // source/rtl/Driver.v(62)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b4  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [4]),
    .sr(rst_n_pad),
    .q(\u1_Driver/hcnt [4]));  // source/rtl/Driver.v(62)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b5  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [5]),
    .sr(rst_n_pad),
    .q(\u1_Driver/hcnt [5]));  // source/rtl/Driver.v(62)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b6  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [6]),
    .sr(rst_n_pad),
    .q(\u1_Driver/hcnt [6]));  // source/rtl/Driver.v(62)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b7  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [7]),
    .sr(rst_n_pad),
    .q(\u1_Driver/hcnt [7]));  // source/rtl/Driver.v(62)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b8  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [8]),
    .sr(rst_n_pad),
    .q(\u1_Driver/hcnt [8]));  // source/rtl/Driver.v(62)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1_Driver/reg1_b9  (
    .clk(clk_vga),
    .d(\u1_Driver/n3 [9]),
    .sr(rst_n_pad),
    .q(\u1_Driver/hcnt [9]));  // source/rtl/Driver.v(62)
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub0/ucin_al_u5021"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub0/u11_al_u5024  (
    .a({open_n2421,\u1_Driver/hcnt [11]}),
    .c(2'b11),
    .d({open_n2426,1'b0}),
    .fci(\u1_Driver/sub0/c11 ),
    .f({open_n2443,\u1_Driver/n20 [11]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub0/ucin_al_u5021"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub0/u3_al_u5022  (
    .a({\u1_Driver/hcnt [5],\u1_Driver/hcnt [3]}),
    .b({\u1_Driver/hcnt [6],\u1_Driver/hcnt [4]}),
    .c(2'b11),
    .d(2'b10),
    .e(2'b10),
    .fci(\u1_Driver/sub0/c3 ),
    .f({\u1_Driver/n20 [5],\u1_Driver/n20 [3]}),
    .fco(\u1_Driver/sub0/c7 ),
    .fx({\u1_Driver/n20 [6],\u1_Driver/n20 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub0/ucin_al_u5021"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub0/u7_al_u5023  (
    .a({\u1_Driver/hcnt [9],\u1_Driver/hcnt [7]}),
    .b({\u1_Driver/hcnt [10],\u1_Driver/hcnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b01),
    .fci(\u1_Driver/sub0/c7 ),
    .f({\u1_Driver/n20 [9],\u1_Driver/n20 [7]}),
    .fco(\u1_Driver/sub0/c11 ),
    .fx({\u1_Driver/n20 [10],\u1_Driver/n20 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub0/ucin_al_u5021"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub0/ucin_al_u5021  (
    .a({\u1_Driver/hcnt [1],1'b0}),
    .b({\u1_Driver/hcnt [2],\u1_Driver/hcnt [0]}),
    .c(2'b11),
    .d(2'b11),
    .e(2'b11),
    .f({\u1_Driver/n20 [1],open_n2502}),
    .fco(\u1_Driver/sub0/c3 ),
    .fx({\u1_Driver/n20 [2],\u1_Driver/n20 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub1/ucin_al_u5025"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub1/u11_al_u5028  (
    .a({open_n2505,\u1_Driver/vcnt [11]}),
    .c(2'b11),
    .d({open_n2510,1'b0}),
    .fci(\u1_Driver/sub1/c11 ),
    .f({open_n2527,\u1_Driver/n21 [11]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub1/ucin_al_u5025"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub1/u3_al_u5026  (
    .a({\u1_Driver/vcnt [5],\u1_Driver/vcnt [3]}),
    .b({\u1_Driver/vcnt [6],\u1_Driver/vcnt [4]}),
    .c(2'b11),
    .d(2'b11),
    .e(2'b00),
    .fci(\u1_Driver/sub1/c3 ),
    .f({\u1_Driver/n21 [5],\u1_Driver/n21 [3]}),
    .fco(\u1_Driver/sub1/c7 ),
    .fx({\u1_Driver/n21 [6],\u1_Driver/n21 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub1/ucin_al_u5025"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub1/u7_al_u5027  (
    .a({\u1_Driver/vcnt [9],\u1_Driver/vcnt [7]}),
    .b({\u1_Driver/vcnt [10],\u1_Driver/vcnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\u1_Driver/sub1/c7 ),
    .f({\u1_Driver/n21 [9],\u1_Driver/n21 [7]}),
    .fco(\u1_Driver/sub1/c11 ),
    .fx({\u1_Driver/n21 [10],\u1_Driver/n21 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1_Driver/sub1/ucin_al_u5025"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1_Driver/sub1/ucin_al_u5025  (
    .a({\u1_Driver/vcnt [1],1'b0}),
    .b({\u1_Driver/vcnt [2],\u1_Driver/vcnt [0]}),
    .c(2'b11),
    .d(2'b01),
    .e(2'b01),
    .f({\u1_Driver/n21 [1],open_n2586}),
    .fco(\u1_Driver/sub1/c3 ),
    .fx({\u1_Driver/n21 [2],\u1_Driver/n21 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u11_al_u5008  (
    .a({\u2_Display/n [13],\u2_Display/n [11]}),
    .b({\u2_Display/n [14],\u2_Display/n [12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c11 ),
    .f({\u2_Display/n37 [13],\u2_Display/n37 [11]}),
    .fco(\u2_Display/add0/c15 ),
    .fx({\u2_Display/n37 [14],\u2_Display/n37 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u15_al_u5009  (
    .a({\u2_Display/n [17],\u2_Display/n [15]}),
    .b({\u2_Display/n [18],\u2_Display/n [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c15 ),
    .f({\u2_Display/n37 [17],\u2_Display/n37 [15]}),
    .fco(\u2_Display/add0/c19 ),
    .fx({\u2_Display/n37 [18],\u2_Display/n37 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u19_al_u5010  (
    .a({\u2_Display/n [21],\u2_Display/n [19]}),
    .b({\u2_Display/n [22],\u2_Display/n [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c19 ),
    .f({\u2_Display/n37 [21],\u2_Display/n37 [19]}),
    .fco(\u2_Display/add0/c23 ),
    .fx({\u2_Display/n37 [22],\u2_Display/n37 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u23_al_u5011  (
    .a({\u2_Display/n [25],\u2_Display/n [23]}),
    .b({\u2_Display/n [26],\u2_Display/n [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c23 ),
    .f({\u2_Display/n37 [25],\u2_Display/n37 [23]}),
    .fco(\u2_Display/add0/c27 ),
    .fx({\u2_Display/n37 [26],\u2_Display/n37 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u27_al_u5012  (
    .a({\u2_Display/n [29],\u2_Display/n [27]}),
    .b({\u2_Display/n [30],\u2_Display/n [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c27 ),
    .f({\u2_Display/n37 [29],\u2_Display/n37 [27]}),
    .fx({\u2_Display/n37 [30],\u2_Display/n37 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u3_al_u5006  (
    .a({\u2_Display/n [5],\u2_Display/n [3]}),
    .b({\u2_Display/n [6],\u2_Display/n [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c3 ),
    .f({\u2_Display/n37 [5],\u2_Display/n37 [3]}),
    .fco(\u2_Display/add0/c7 ),
    .fx({\u2_Display/n37 [6],\u2_Display/n37 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/u7_al_u5007  (
    .a({\u2_Display/n [9],\u2_Display/n [7]}),
    .b({\u2_Display/n [10],\u2_Display/n [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add0/c7 ),
    .f({\u2_Display/n37 [9],\u2_Display/n37 [7]}),
    .fco(\u2_Display/add0/c11 ),
    .fx({\u2_Display/n37 [10],\u2_Display/n37 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add0/ucin_al_u5005"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add0/ucin_al_u5005  (
    .a({\u2_Display/n [1],1'b0}),
    .b({\u2_Display/n [2],\u2_Display/n [0]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .f({\u2_Display/n37 [1],open_n2733}),
    .fco(\u2_Display/add0/c3 ),
    .fx({\u2_Display/n37 [2],\u2_Display/n37 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u11_al_u4009  (
    .a({\u2_Display/counta [13],\u2_Display/counta [11]}),
    .b({\u2_Display/counta [14],\u2_Display/counta [12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c11 ),
    .f({\u2_Display/n41 [13],\u2_Display/n41 [11]}),
    .fco(\u2_Display/add1/c15 ),
    .fx({\u2_Display/n41 [14],\u2_Display/n41 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u15_al_u4010  (
    .a({\u2_Display/counta [17],\u2_Display/counta [15]}),
    .b({\u2_Display/counta [18],\u2_Display/counta [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c15 ),
    .f({\u2_Display/n41 [17],\u2_Display/n41 [15]}),
    .fco(\u2_Display/add1/c19 ),
    .fx({\u2_Display/n41 [18],\u2_Display/n41 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u19_al_u4011  (
    .a({\u2_Display/counta [21],\u2_Display/counta [19]}),
    .b({\u2_Display/counta [22],\u2_Display/counta [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c19 ),
    .f({\u2_Display/n41 [21],\u2_Display/n41 [19]}),
    .fco(\u2_Display/add1/c23 ),
    .fx({\u2_Display/n41 [22],\u2_Display/n41 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u23_al_u4012  (
    .a({\u2_Display/counta [25],\u2_Display/counta [23]}),
    .b({\u2_Display/counta [26],\u2_Display/counta [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c23 ),
    .f({\u2_Display/n41 [25],\u2_Display/n41 [23]}),
    .fco(\u2_Display/add1/c27 ),
    .fx({\u2_Display/n41 [26],\u2_Display/n41 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u27_al_u4013  (
    .a({\u2_Display/counta [29],\u2_Display/counta [27]}),
    .b({\u2_Display/counta [30],\u2_Display/counta [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c27 ),
    .f({\u2_Display/n41 [29],\u2_Display/n41 [27]}),
    .fco(\u2_Display/add1/c31 ),
    .fx({\u2_Display/n41 [30],\u2_Display/n41 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u31_al_u4014  (
    .a({open_n2826,\u2_Display/counta [31]}),
    .c(2'b00),
    .d({open_n2831,1'b0}),
    .fci(\u2_Display/add1/c31 ),
    .f({open_n2848,\u2_Display/n41 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u3_al_u4007  (
    .a({\u2_Display/counta [5],\u2_Display/counta [3]}),
    .b({\u2_Display/counta [6],\u2_Display/counta [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c3 ),
    .f({\u2_Display/n41 [5],\u2_Display/n41 [3]}),
    .fco(\u2_Display/add1/c7 ),
    .fx({\u2_Display/n41 [6],\u2_Display/n41 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/u7_al_u4008  (
    .a({\u2_Display/counta [9],\u2_Display/counta [7]}),
    .b({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add1/c7 ),
    .f({\u2_Display/n41 [9],\u2_Display/n41 [7]}),
    .fco(\u2_Display/add1/c11 ),
    .fx({\u2_Display/n41 [10],\u2_Display/n41 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add1/ucin_al_u4006"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add1/ucin_al_u4006  (
    .a({\u2_Display/counta [1],1'b0}),
    .b({\u2_Display/counta [2],\u2_Display/counta [0]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .f({\u2_Display/n41 [1],open_n2907}),
    .fco(\u2_Display/add1/c3 ),
    .fx({\u2_Display/n41 [2],\u2_Display/n41 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u11_al_u4018  (
    .a({\u2_Display/n3209 ,\u2_Display/n3211 }),
    .b({\u2_Display/n3208 ,\u2_Display/n3210 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add100/c11 ),
    .f({\u2_Display/n3225 [13],\u2_Display/n3225 [11]}),
    .fco(\u2_Display/add100/c15 ),
    .fx({\u2_Display/n3225 [14],\u2_Display/n3225 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u15_al_u4019  (
    .a({\u2_Display/n3205 ,\u2_Display/n3207 }),
    .b({\u2_Display/n3204 ,\u2_Display/n3206 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add100/c15 ),
    .f({\u2_Display/n3225 [17],\u2_Display/n3225 [15]}),
    .fco(\u2_Display/add100/c19 ),
    .fx({\u2_Display/n3225 [18],\u2_Display/n3225 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u19_al_u4020  (
    .a({\u2_Display/n3201 ,\u2_Display/n3203 }),
    .b({\u2_Display/n3200 ,\u2_Display/n3202 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add100/c19 ),
    .f({\u2_Display/n3225 [21],\u2_Display/n3225 [19]}),
    .fco(\u2_Display/add100/c23 ),
    .fx({\u2_Display/n3225 [22],\u2_Display/n3225 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u23_al_u4021  (
    .a({\u2_Display/n3197 ,\u2_Display/n3199 }),
    .b({\u2_Display/n3196 ,\u2_Display/n3198 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add100/c23 ),
    .f({\u2_Display/n3225 [25],\u2_Display/n3225 [23]}),
    .fco(\u2_Display/add100/c27 ),
    .fx({\u2_Display/n3225 [26],\u2_Display/n3225 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u27_al_u4022  (
    .a({\u2_Display/n3193 ,\u2_Display/n3195 }),
    .b({\u2_Display/n3192 ,\u2_Display/n3194 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add100/c27 ),
    .f({\u2_Display/n3225 [29],\u2_Display/n3225 [27]}),
    .fco(\u2_Display/add100/c31 ),
    .fx({\u2_Display/n3225 [30],\u2_Display/n3225 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u31_al_u4023  (
    .a({open_n3000,\u2_Display/n3191 }),
    .c(2'b00),
    .d({open_n3005,1'b1}),
    .fci(\u2_Display/add100/c31 ),
    .f({open_n3022,\u2_Display/n3225 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u3_al_u4016  (
    .a({\u2_Display/n3217 ,\u2_Display/n3219 }),
    .b({\u2_Display/n3216 ,\u2_Display/n3218 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add100/c3 ),
    .f({\u2_Display/n3225 [5],\u2_Display/n3225 [3]}),
    .fco(\u2_Display/add100/c7 ),
    .fx({\u2_Display/n3225 [6],\u2_Display/n3225 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/u7_al_u4017  (
    .a({\u2_Display/n3213 ,\u2_Display/n3215 }),
    .b({\u2_Display/n3212 ,\u2_Display/n3214 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add100/c7 ),
    .f({\u2_Display/n3225 [9],\u2_Display/n3225 [7]}),
    .fco(\u2_Display/add100/c11 ),
    .fx({\u2_Display/n3225 [10],\u2_Display/n3225 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add100/ucin_al_u4015"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add100/ucin_al_u4015  (
    .a({\u2_Display/n3221 ,1'b1}),
    .b({\u2_Display/n3220 ,\u2_Display/n3222 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3225 [1],open_n3081}),
    .fco(\u2_Display/add100/c3 ),
    .fx({\u2_Display/n3225 [2],\u2_Display/n3225 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u11_al_u4027  (
    .a({\u2_Display/n3244 ,\u2_Display/n3246 }),
    .b({\u2_Display/n3243 ,\u2_Display/n3245 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add101/c11 ),
    .f({\u2_Display/n3260 [13],\u2_Display/n3260 [11]}),
    .fco(\u2_Display/add101/c15 ),
    .fx({\u2_Display/n3260 [14],\u2_Display/n3260 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u15_al_u4028  (
    .a({\u2_Display/n3240 ,\u2_Display/n3242 }),
    .b({\u2_Display/n3239 ,\u2_Display/n3241 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add101/c15 ),
    .f({\u2_Display/n3260 [17],\u2_Display/n3260 [15]}),
    .fco(\u2_Display/add101/c19 ),
    .fx({\u2_Display/n3260 [18],\u2_Display/n3260 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u19_al_u4029  (
    .a({\u2_Display/n3236 ,\u2_Display/n3238 }),
    .b({\u2_Display/n3235 ,\u2_Display/n3237 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add101/c19 ),
    .f({\u2_Display/n3260 [21],\u2_Display/n3260 [19]}),
    .fco(\u2_Display/add101/c23 ),
    .fx({\u2_Display/n3260 [22],\u2_Display/n3260 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u23_al_u4030  (
    .a({\u2_Display/n3232 ,\u2_Display/n3234 }),
    .b({\u2_Display/n3231 ,\u2_Display/n3233 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add101/c23 ),
    .f({\u2_Display/n3260 [25],\u2_Display/n3260 [23]}),
    .fco(\u2_Display/add101/c27 ),
    .fx({\u2_Display/n3260 [26],\u2_Display/n3260 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u27_al_u4031  (
    .a({\u2_Display/n3228 ,\u2_Display/n3230 }),
    .b({\u2_Display/n3227 ,\u2_Display/n3229 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add101/c27 ),
    .f({\u2_Display/n3260 [29],\u2_Display/n3260 [27]}),
    .fco(\u2_Display/add101/c31 ),
    .fx({\u2_Display/n3260 [30],\u2_Display/n3260 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u31_al_u4032  (
    .a({open_n3174,\u2_Display/n3226 }),
    .c(2'b00),
    .d({open_n3179,1'b1}),
    .fci(\u2_Display/add101/c31 ),
    .f({open_n3196,\u2_Display/n3260 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u3_al_u4025  (
    .a({\u2_Display/n3252 ,\u2_Display/n3254 }),
    .b({\u2_Display/n3251 ,\u2_Display/n3253 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add101/c3 ),
    .f({\u2_Display/n3260 [5],\u2_Display/n3260 [3]}),
    .fco(\u2_Display/add101/c7 ),
    .fx({\u2_Display/n3260 [6],\u2_Display/n3260 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/u7_al_u4026  (
    .a({\u2_Display/n3248 ,\u2_Display/n3250 }),
    .b({\u2_Display/n3247 ,\u2_Display/n3249 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add101/c7 ),
    .f({\u2_Display/n3260 [9],\u2_Display/n3260 [7]}),
    .fco(\u2_Display/add101/c11 ),
    .fx({\u2_Display/n3260 [10],\u2_Display/n3260 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add101/ucin_al_u4024"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add101/ucin_al_u4024  (
    .a({\u2_Display/n3256 ,1'b1}),
    .b({\u2_Display/n3255 ,\u2_Display/n3257 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3260 [1],open_n3255}),
    .fco(\u2_Display/add101/c3 ),
    .fx({\u2_Display/n3260 [2],\u2_Display/n3260 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u11_al_u4036  (
    .a({\u2_Display/n3279 ,\u2_Display/n3281 }),
    .b({\u2_Display/n3278 ,\u2_Display/n3280 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add102/c11 ),
    .f({\u2_Display/n3295 [13],\u2_Display/n3295 [11]}),
    .fco(\u2_Display/add102/c15 ),
    .fx({\u2_Display/n3295 [14],\u2_Display/n3295 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u15_al_u4037  (
    .a({\u2_Display/n3275 ,\u2_Display/n3277 }),
    .b({\u2_Display/n3274 ,\u2_Display/n3276 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add102/c15 ),
    .f({\u2_Display/n3295 [17],\u2_Display/n3295 [15]}),
    .fco(\u2_Display/add102/c19 ),
    .fx({\u2_Display/n3295 [18],\u2_Display/n3295 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u19_al_u4038  (
    .a({\u2_Display/n3271 ,\u2_Display/n3273 }),
    .b({\u2_Display/n3270 ,\u2_Display/n3272 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add102/c19 ),
    .f({\u2_Display/n3295 [21],\u2_Display/n3295 [19]}),
    .fco(\u2_Display/add102/c23 ),
    .fx({\u2_Display/n3295 [22],\u2_Display/n3295 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u23_al_u4039  (
    .a({\u2_Display/n3267 ,\u2_Display/n3269 }),
    .b({\u2_Display/n3266 ,\u2_Display/n3268 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add102/c23 ),
    .f({\u2_Display/n3295 [25],\u2_Display/n3295 [23]}),
    .fco(\u2_Display/add102/c27 ),
    .fx({\u2_Display/n3295 [26],\u2_Display/n3295 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u27_al_u4040  (
    .a({\u2_Display/n3263 ,\u2_Display/n3265 }),
    .b({\u2_Display/n3262 ,\u2_Display/n3264 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add102/c27 ),
    .f({\u2_Display/n3295 [29],\u2_Display/n3295 [27]}),
    .fco(\u2_Display/add102/c31 ),
    .fx({\u2_Display/n3295 [30],\u2_Display/n3295 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u31_al_u4041  (
    .a({open_n3348,\u2_Display/n3261 }),
    .c(2'b00),
    .d({open_n3353,1'b1}),
    .fci(\u2_Display/add102/c31 ),
    .f({open_n3370,\u2_Display/n3295 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u3_al_u4034  (
    .a({\u2_Display/n3287 ,\u2_Display/n3289 }),
    .b({\u2_Display/n3286 ,\u2_Display/n3288 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add102/c3 ),
    .f({\u2_Display/n3295 [5],\u2_Display/n3295 [3]}),
    .fco(\u2_Display/add102/c7 ),
    .fx({\u2_Display/n3295 [6],\u2_Display/n3295 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/u7_al_u4035  (
    .a({\u2_Display/n3283 ,\u2_Display/n3285 }),
    .b({\u2_Display/n3282 ,\u2_Display/n3284 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b00),
    .fci(\u2_Display/add102/c7 ),
    .f({\u2_Display/n3295 [9],\u2_Display/n3295 [7]}),
    .fco(\u2_Display/add102/c11 ),
    .fx({\u2_Display/n3295 [10],\u2_Display/n3295 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add102/ucin_al_u4033"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add102/ucin_al_u4033  (
    .a({\u2_Display/n3291 ,1'b1}),
    .b({\u2_Display/n3290 ,\u2_Display/n3292 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3295 [1],open_n3429}),
    .fco(\u2_Display/add102/c3 ),
    .fx({\u2_Display/n3295 [2],\u2_Display/n3295 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u11_al_u4045  (
    .a({\u2_Display/n3314 ,\u2_Display/n3316 }),
    .b({\u2_Display/n3313 ,\u2_Display/n3315 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add103/c11 ),
    .f({\u2_Display/n3330 [13],\u2_Display/n3330 [11]}),
    .fco(\u2_Display/add103/c15 ),
    .fx({\u2_Display/n3330 [14],\u2_Display/n3330 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u15_al_u4046  (
    .a({\u2_Display/n3310 ,\u2_Display/n3312 }),
    .b({\u2_Display/n3309 ,\u2_Display/n3311 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add103/c15 ),
    .f({\u2_Display/n3330 [17],\u2_Display/n3330 [15]}),
    .fco(\u2_Display/add103/c19 ),
    .fx({\u2_Display/n3330 [18],\u2_Display/n3330 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u19_al_u4047  (
    .a({\u2_Display/n3306 ,\u2_Display/n3308 }),
    .b({\u2_Display/n3305 ,\u2_Display/n3307 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add103/c19 ),
    .f({\u2_Display/n3330 [21],\u2_Display/n3330 [19]}),
    .fco(\u2_Display/add103/c23 ),
    .fx({\u2_Display/n3330 [22],\u2_Display/n3330 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u23_al_u4048  (
    .a({\u2_Display/n3302 ,\u2_Display/n3304 }),
    .b({\u2_Display/n3301 ,\u2_Display/n3303 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add103/c23 ),
    .f({\u2_Display/n3330 [25],\u2_Display/n3330 [23]}),
    .fco(\u2_Display/add103/c27 ),
    .fx({\u2_Display/n3330 [26],\u2_Display/n3330 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u27_al_u4049  (
    .a({\u2_Display/n3298 ,\u2_Display/n3300 }),
    .b({\u2_Display/n3297 ,\u2_Display/n3299 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add103/c27 ),
    .f({\u2_Display/n3330 [29],\u2_Display/n3330 [27]}),
    .fco(\u2_Display/add103/c31 ),
    .fx({\u2_Display/n3330 [30],\u2_Display/n3330 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u31_al_u4050  (
    .a({open_n3522,\u2_Display/n3296 }),
    .c(2'b00),
    .d({open_n3527,1'b1}),
    .fci(\u2_Display/add103/c31 ),
    .f({open_n3544,\u2_Display/n3330 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u3_al_u4043  (
    .a({\u2_Display/n3322 ,\u2_Display/n3324 }),
    .b({\u2_Display/n3321 ,\u2_Display/n3323 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add103/c3 ),
    .f({\u2_Display/n3330 [5],\u2_Display/n3330 [3]}),
    .fco(\u2_Display/add103/c7 ),
    .fx({\u2_Display/n3330 [6],\u2_Display/n3330 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/u7_al_u4044  (
    .a({\u2_Display/n3318 ,\u2_Display/n3320 }),
    .b({\u2_Display/n3317 ,\u2_Display/n3319 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add103/c7 ),
    .f({\u2_Display/n3330 [9],\u2_Display/n3330 [7]}),
    .fco(\u2_Display/add103/c11 ),
    .fx({\u2_Display/n3330 [10],\u2_Display/n3330 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add103/ucin_al_u4042"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add103/ucin_al_u4042  (
    .a({\u2_Display/n3326 ,1'b1}),
    .b({\u2_Display/n3325 ,\u2_Display/n3327 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3330 [1],open_n3603}),
    .fco(\u2_Display/add103/c3 ),
    .fx({\u2_Display/n3330 [2],\u2_Display/n3330 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u11_al_u4054  (
    .a({\u2_Display/n3349 ,\u2_Display/n3351 }),
    .b({\u2_Display/n3348 ,\u2_Display/n3350 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add104/c11 ),
    .f({\u2_Display/n3365 [13],\u2_Display/n3365 [11]}),
    .fco(\u2_Display/add104/c15 ),
    .fx({\u2_Display/n3365 [14],\u2_Display/n3365 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u15_al_u4055  (
    .a({\u2_Display/n3345 ,\u2_Display/n3347 }),
    .b({\u2_Display/n3344 ,\u2_Display/n3346 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add104/c15 ),
    .f({\u2_Display/n3365 [17],\u2_Display/n3365 [15]}),
    .fco(\u2_Display/add104/c19 ),
    .fx({\u2_Display/n3365 [18],\u2_Display/n3365 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u19_al_u4056  (
    .a({\u2_Display/n3341 ,\u2_Display/n3343 }),
    .b({\u2_Display/n3340 ,\u2_Display/n3342 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add104/c19 ),
    .f({\u2_Display/n3365 [21],\u2_Display/n3365 [19]}),
    .fco(\u2_Display/add104/c23 ),
    .fx({\u2_Display/n3365 [22],\u2_Display/n3365 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u23_al_u4057  (
    .a({\u2_Display/n3337 ,\u2_Display/n3339 }),
    .b({\u2_Display/n3336 ,\u2_Display/n3338 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add104/c23 ),
    .f({\u2_Display/n3365 [25],\u2_Display/n3365 [23]}),
    .fco(\u2_Display/add104/c27 ),
    .fx({\u2_Display/n3365 [26],\u2_Display/n3365 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u27_al_u4058  (
    .a({\u2_Display/n3333 ,\u2_Display/n3335 }),
    .b({\u2_Display/n3332 ,\u2_Display/n3334 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add104/c27 ),
    .f({\u2_Display/n3365 [29],\u2_Display/n3365 [27]}),
    .fco(\u2_Display/add104/c31 ),
    .fx({\u2_Display/n3365 [30],\u2_Display/n3365 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u31_al_u4059  (
    .a({open_n3696,\u2_Display/n3331 }),
    .c(2'b00),
    .d({open_n3701,1'b1}),
    .fci(\u2_Display/add104/c31 ),
    .f({open_n3718,\u2_Display/n3365 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u3_al_u4052  (
    .a({\u2_Display/n3357 ,\u2_Display/n3359 }),
    .b({\u2_Display/n3356 ,\u2_Display/n3358 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add104/c3 ),
    .f({\u2_Display/n3365 [5],\u2_Display/n3365 [3]}),
    .fco(\u2_Display/add104/c7 ),
    .fx({\u2_Display/n3365 [6],\u2_Display/n3365 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/u7_al_u4053  (
    .a({\u2_Display/n3353 ,\u2_Display/n3355 }),
    .b({\u2_Display/n3352 ,\u2_Display/n3354 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add104/c7 ),
    .f({\u2_Display/n3365 [9],\u2_Display/n3365 [7]}),
    .fco(\u2_Display/add104/c11 ),
    .fx({\u2_Display/n3365 [10],\u2_Display/n3365 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add104/ucin_al_u4051"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add104/ucin_al_u4051  (
    .a({\u2_Display/n3361 ,1'b1}),
    .b({\u2_Display/n3360 ,\u2_Display/n3362 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3365 [1],open_n3777}),
    .fco(\u2_Display/add104/c3 ),
    .fx({\u2_Display/n3365 [2],\u2_Display/n3365 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u11_al_u4063  (
    .a({\u2_Display/n3384 ,\u2_Display/n3386 }),
    .b({\u2_Display/n3383 ,\u2_Display/n3385 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add105/c11 ),
    .f({\u2_Display/n3400 [13],\u2_Display/n3400 [11]}),
    .fco(\u2_Display/add105/c15 ),
    .fx({\u2_Display/n3400 [14],\u2_Display/n3400 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u15_al_u4064  (
    .a({\u2_Display/n3380 ,\u2_Display/n3382 }),
    .b({\u2_Display/n3379 ,\u2_Display/n3381 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add105/c15 ),
    .f({\u2_Display/n3400 [17],\u2_Display/n3400 [15]}),
    .fco(\u2_Display/add105/c19 ),
    .fx({\u2_Display/n3400 [18],\u2_Display/n3400 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u19_al_u4065  (
    .a({\u2_Display/n3376 ,\u2_Display/n3378 }),
    .b({\u2_Display/n3375 ,\u2_Display/n3377 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add105/c19 ),
    .f({\u2_Display/n3400 [21],\u2_Display/n3400 [19]}),
    .fco(\u2_Display/add105/c23 ),
    .fx({\u2_Display/n3400 [22],\u2_Display/n3400 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u23_al_u4066  (
    .a({\u2_Display/n3372 ,\u2_Display/n3374 }),
    .b({\u2_Display/n3371 ,\u2_Display/n3373 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add105/c23 ),
    .f({\u2_Display/n3400 [25],\u2_Display/n3400 [23]}),
    .fco(\u2_Display/add105/c27 ),
    .fx({\u2_Display/n3400 [26],\u2_Display/n3400 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u27_al_u4067  (
    .a({\u2_Display/n3368 ,\u2_Display/n3370 }),
    .b({\u2_Display/n3367 ,\u2_Display/n3369 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add105/c27 ),
    .f({\u2_Display/n3400 [29],\u2_Display/n3400 [27]}),
    .fco(\u2_Display/add105/c31 ),
    .fx({\u2_Display/n3400 [30],\u2_Display/n3400 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u31_al_u4068  (
    .a({open_n3870,\u2_Display/n3366 }),
    .c(2'b00),
    .d({open_n3875,1'b1}),
    .fci(\u2_Display/add105/c31 ),
    .f({open_n3892,\u2_Display/n3400 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u3_al_u4061  (
    .a({\u2_Display/n3392 ,\u2_Display/n3394 }),
    .b({\u2_Display/n3391 ,\u2_Display/n3393 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add105/c3 ),
    .f({\u2_Display/n3400 [5],\u2_Display/n3400 [3]}),
    .fco(\u2_Display/add105/c7 ),
    .fx({\u2_Display/n3400 [6],\u2_Display/n3400 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/u7_al_u4062  (
    .a({\u2_Display/n3388 ,\u2_Display/n3390 }),
    .b({\u2_Display/n3387 ,\u2_Display/n3389 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add105/c7 ),
    .f({\u2_Display/n3400 [9],\u2_Display/n3400 [7]}),
    .fco(\u2_Display/add105/c11 ),
    .fx({\u2_Display/n3400 [10],\u2_Display/n3400 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add105/ucin_al_u4060"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add105/ucin_al_u4060  (
    .a({\u2_Display/n3396 ,1'b1}),
    .b({\u2_Display/n3395 ,\u2_Display/n3397 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3400 [1],open_n3951}),
    .fco(\u2_Display/add105/c3 ),
    .fx({\u2_Display/n3400 [2],\u2_Display/n3400 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add106/ucin_al_u5043"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add106/u3_al_u5044  (
    .a({\u2_Display/n3427 ,\u2_Display/n3429 }),
    .b({\u2_Display/n3426 ,\u2_Display/n3428 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b00),
    .fci(\u2_Display/add106/c3 ),
    .f({\u2_Display/n3435 [5],\u2_Display/n3435 [3]}),
    .fco(\u2_Display/add106/c7 ),
    .fx({\u2_Display/n3435 [6],\u2_Display/n3435 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add106/ucin_al_u5043"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add106/u7_al_u5045  (
    .a({\u2_Display/n3423 ,\u2_Display/n3425 }),
    .b({open_n3972,\u2_Display/n3424 }),
    .c(2'b00),
    .d(2'b01),
    .e({open_n3975,1'b1}),
    .fci(\u2_Display/add106/c7 ),
    .f({\u2_Display/n3435 [9],\u2_Display/n3435 [7]}),
    .fx({open_n3991,\u2_Display/n3435 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add106/ucin_al_u5043"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add106/ucin_al_u5043  (
    .a({\u2_Display/n3431 ,1'b1}),
    .b({\u2_Display/n3430 ,\u2_Display/n3432 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3435 [1],open_n4011}),
    .fco(\u2_Display/add106/c3 ),
    .fx({\u2_Display/n3435 [2],\u2_Display/n3435 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u11_al_u4072  (
    .a({\u2_Display/counta [13],\u2_Display/counta [11]}),
    .b({\u2_Display/counta [14],\u2_Display/counta [12]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add117/c11 ),
    .f({\u2_Display/n3788 [13],\u2_Display/n3788 [11]}),
    .fco(\u2_Display/add117/c15 ),
    .fx({\u2_Display/n3788 [14],\u2_Display/n3788 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u15_al_u4073  (
    .a({\u2_Display/counta [17],\u2_Display/counta [15]}),
    .b({\u2_Display/counta [18],\u2_Display/counta [16]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add117/c15 ),
    .f({\u2_Display/n3788 [17],\u2_Display/n3788 [15]}),
    .fco(\u2_Display/add117/c19 ),
    .fx({\u2_Display/n3788 [18],\u2_Display/n3788 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u19_al_u4074  (
    .a({\u2_Display/counta [21],\u2_Display/counta [19]}),
    .b({\u2_Display/counta [22],\u2_Display/counta [20]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add117/c19 ),
    .f({\u2_Display/n3788 [21],\u2_Display/n3788 [19]}),
    .fco(\u2_Display/add117/c23 ),
    .fx({\u2_Display/n3788 [22],\u2_Display/n3788 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u23_al_u4075  (
    .a({\u2_Display/counta [25],\u2_Display/counta [23]}),
    .b({\u2_Display/counta [26],\u2_Display/counta [24]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add117/c23 ),
    .f({\u2_Display/n3788 [25],\u2_Display/n3788 [23]}),
    .fco(\u2_Display/add117/c27 ),
    .fx({\u2_Display/n3788 [26],\u2_Display/n3788 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u27_al_u4076  (
    .a({\u2_Display/counta [29],\u2_Display/counta [27]}),
    .b({\u2_Display/counta [30],\u2_Display/counta [28]}),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add117/c27 ),
    .f({\u2_Display/n3788 [29],\u2_Display/n3788 [27]}),
    .fco(\u2_Display/add117/c31 ),
    .fx({\u2_Display/n3788 [30],\u2_Display/n3788 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u31_al_u4077  (
    .a({open_n4104,\u2_Display/counta [31]}),
    .c(2'b00),
    .d({open_n4109,1'b0}),
    .fci(\u2_Display/add117/c31 ),
    .f({open_n4126,\u2_Display/n3788 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u3_al_u4070  (
    .a({\u2_Display/counta [5],\u2_Display/counta [3]}),
    .b({\u2_Display/counta [6],\u2_Display/counta [4]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add117/c3 ),
    .f({\u2_Display/n3788 [5],\u2_Display/n3788 [3]}),
    .fco(\u2_Display/add117/c7 ),
    .fx({\u2_Display/n3788 [6],\u2_Display/n3788 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/u7_al_u4071  (
    .a({\u2_Display/counta [9],\u2_Display/counta [7]}),
    .b({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add117/c7 ),
    .f({\u2_Display/n3788 [9],\u2_Display/n3788 [7]}),
    .fco(\u2_Display/add117/c11 ),
    .fx({\u2_Display/n3788 [10],\u2_Display/n3788 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add117/ucin_al_u4069"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add117/ucin_al_u4069  (
    .a({\u2_Display/counta [1],1'b1}),
    .b({\u2_Display/counta [2],\u2_Display/counta [0]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3788 [1],open_n4185}),
    .fco(\u2_Display/add117/c3 ),
    .fx({\u2_Display/n3788 [2],\u2_Display/n3788 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u11_al_u4081  (
    .a({\u2_Display/n3807 ,\u2_Display/n3809 }),
    .b({\u2_Display/n3806 ,\u2_Display/n3808 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add118/c11 ),
    .f({\u2_Display/n3823 [13],\u2_Display/n3823 [11]}),
    .fco(\u2_Display/add118/c15 ),
    .fx({\u2_Display/n3823 [14],\u2_Display/n3823 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u15_al_u4082  (
    .a({\u2_Display/n3803 ,\u2_Display/n3805 }),
    .b({\u2_Display/n3802 ,\u2_Display/n3804 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add118/c15 ),
    .f({\u2_Display/n3823 [17],\u2_Display/n3823 [15]}),
    .fco(\u2_Display/add118/c19 ),
    .fx({\u2_Display/n3823 [18],\u2_Display/n3823 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u19_al_u4083  (
    .a({\u2_Display/n3799 ,\u2_Display/n3801 }),
    .b({\u2_Display/n3798 ,\u2_Display/n3800 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add118/c19 ),
    .f({\u2_Display/n3823 [21],\u2_Display/n3823 [19]}),
    .fco(\u2_Display/add118/c23 ),
    .fx({\u2_Display/n3823 [22],\u2_Display/n3823 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u23_al_u4084  (
    .a({\u2_Display/n3795 ,\u2_Display/n3797 }),
    .b({\u2_Display/n3794 ,\u2_Display/n3796 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add118/c23 ),
    .f({\u2_Display/n3823 [25],\u2_Display/n3823 [23]}),
    .fco(\u2_Display/add118/c27 ),
    .fx({\u2_Display/n3823 [26],\u2_Display/n3823 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u27_al_u4085  (
    .a({\u2_Display/n3791 ,\u2_Display/n3793 }),
    .b({\u2_Display/n3790 ,\u2_Display/n3792 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add118/c27 ),
    .f({\u2_Display/n3823 [29],\u2_Display/n3823 [27]}),
    .fco(\u2_Display/add118/c31 ),
    .fx({\u2_Display/n3823 [30],\u2_Display/n3823 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u31_al_u4086  (
    .a({open_n4278,\u2_Display/n3789 }),
    .c(2'b00),
    .d({open_n4283,1'b1}),
    .fci(\u2_Display/add118/c31 ),
    .f({open_n4300,\u2_Display/n3823 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u3_al_u4079  (
    .a({\u2_Display/n3815 ,\u2_Display/n3817 }),
    .b({\u2_Display/n3814 ,\u2_Display/n3816 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add118/c3 ),
    .f({\u2_Display/n3823 [5],\u2_Display/n3823 [3]}),
    .fco(\u2_Display/add118/c7 ),
    .fx({\u2_Display/n3823 [6],\u2_Display/n3823 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/u7_al_u4080  (
    .a({\u2_Display/n3811 ,\u2_Display/n3813 }),
    .b({\u2_Display/n3810 ,\u2_Display/n3812 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add118/c7 ),
    .f({\u2_Display/n3823 [9],\u2_Display/n3823 [7]}),
    .fco(\u2_Display/add118/c11 ),
    .fx({\u2_Display/n3823 [10],\u2_Display/n3823 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add118/ucin_al_u4078"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add118/ucin_al_u4078  (
    .a({\u2_Display/n3819 ,1'b1}),
    .b({\u2_Display/n3818 ,\u2_Display/n3820 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3823 [1],open_n4359}),
    .fco(\u2_Display/add118/c3 ),
    .fx({\u2_Display/n3823 [2],\u2_Display/n3823 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u11_al_u4090  (
    .a({\u2_Display/n3842 ,\u2_Display/n3844 }),
    .b({\u2_Display/n3841 ,\u2_Display/n3843 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add119/c11 ),
    .f({\u2_Display/n3858 [13],\u2_Display/n3858 [11]}),
    .fco(\u2_Display/add119/c15 ),
    .fx({\u2_Display/n3858 [14],\u2_Display/n3858 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u15_al_u4091  (
    .a({\u2_Display/n3838 ,\u2_Display/n3840 }),
    .b({\u2_Display/n3837 ,\u2_Display/n3839 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add119/c15 ),
    .f({\u2_Display/n3858 [17],\u2_Display/n3858 [15]}),
    .fco(\u2_Display/add119/c19 ),
    .fx({\u2_Display/n3858 [18],\u2_Display/n3858 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u19_al_u4092  (
    .a({\u2_Display/n3834 ,\u2_Display/n3836 }),
    .b({\u2_Display/n3833 ,\u2_Display/n3835 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add119/c19 ),
    .f({\u2_Display/n3858 [21],\u2_Display/n3858 [19]}),
    .fco(\u2_Display/add119/c23 ),
    .fx({\u2_Display/n3858 [22],\u2_Display/n3858 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u23_al_u4093  (
    .a({\u2_Display/n3830 ,\u2_Display/n3832 }),
    .b({\u2_Display/n3829 ,\u2_Display/n3831 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add119/c23 ),
    .f({\u2_Display/n3858 [25],\u2_Display/n3858 [23]}),
    .fco(\u2_Display/add119/c27 ),
    .fx({\u2_Display/n3858 [26],\u2_Display/n3858 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u27_al_u4094  (
    .a({\u2_Display/n3826 ,\u2_Display/n3828 }),
    .b({\u2_Display/n3825 ,\u2_Display/n3827 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add119/c27 ),
    .f({\u2_Display/n3858 [29],\u2_Display/n3858 [27]}),
    .fco(\u2_Display/add119/c31 ),
    .fx({\u2_Display/n3858 [30],\u2_Display/n3858 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u31_al_u4095  (
    .a({open_n4452,\u2_Display/n3824 }),
    .c(2'b00),
    .d({open_n4457,1'b1}),
    .fci(\u2_Display/add119/c31 ),
    .f({open_n4474,\u2_Display/n3858 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u3_al_u4088  (
    .a({\u2_Display/n3850 ,\u2_Display/n3852 }),
    .b({\u2_Display/n3849 ,\u2_Display/n3851 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add119/c3 ),
    .f({\u2_Display/n3858 [5],\u2_Display/n3858 [3]}),
    .fco(\u2_Display/add119/c7 ),
    .fx({\u2_Display/n3858 [6],\u2_Display/n3858 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/u7_al_u4089  (
    .a({\u2_Display/n3846 ,\u2_Display/n3848 }),
    .b({\u2_Display/n3845 ,\u2_Display/n3847 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add119/c7 ),
    .f({\u2_Display/n3858 [9],\u2_Display/n3858 [7]}),
    .fco(\u2_Display/add119/c11 ),
    .fx({\u2_Display/n3858 [10],\u2_Display/n3858 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add119/ucin_al_u4087"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add119/ucin_al_u4087  (
    .a({\u2_Display/n3854 ,1'b1}),
    .b({\u2_Display/n3853 ,\u2_Display/n3855 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3858 [1],open_n4533}),
    .fco(\u2_Display/add119/c3 ),
    .fx({\u2_Display/n3858 [2],\u2_Display/n3858 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u11_al_u4099  (
    .a({\u2_Display/n3877 ,\u2_Display/n3879 }),
    .b({\u2_Display/n3876 ,\u2_Display/n3878 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add120/c11 ),
    .f({\u2_Display/n3893 [13],\u2_Display/n3893 [11]}),
    .fco(\u2_Display/add120/c15 ),
    .fx({\u2_Display/n3893 [14],\u2_Display/n3893 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u15_al_u4100  (
    .a({\u2_Display/n3873 ,\u2_Display/n3875 }),
    .b({\u2_Display/n3872 ,\u2_Display/n3874 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add120/c15 ),
    .f({\u2_Display/n3893 [17],\u2_Display/n3893 [15]}),
    .fco(\u2_Display/add120/c19 ),
    .fx({\u2_Display/n3893 [18],\u2_Display/n3893 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u19_al_u4101  (
    .a({\u2_Display/n3869 ,\u2_Display/n3871 }),
    .b({\u2_Display/n3868 ,\u2_Display/n3870 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add120/c19 ),
    .f({\u2_Display/n3893 [21],\u2_Display/n3893 [19]}),
    .fco(\u2_Display/add120/c23 ),
    .fx({\u2_Display/n3893 [22],\u2_Display/n3893 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u23_al_u4102  (
    .a({\u2_Display/n3865 ,\u2_Display/n3867 }),
    .b({\u2_Display/n3864 ,\u2_Display/n3866 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add120/c23 ),
    .f({\u2_Display/n3893 [25],\u2_Display/n3893 [23]}),
    .fco(\u2_Display/add120/c27 ),
    .fx({\u2_Display/n3893 [26],\u2_Display/n3893 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u27_al_u4103  (
    .a({\u2_Display/n3861 ,\u2_Display/n3863 }),
    .b({\u2_Display/n3860 ,\u2_Display/n3862 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add120/c27 ),
    .f({\u2_Display/n3893 [29],\u2_Display/n3893 [27]}),
    .fco(\u2_Display/add120/c31 ),
    .fx({\u2_Display/n3893 [30],\u2_Display/n3893 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u31_al_u4104  (
    .a({open_n4626,\u2_Display/n3859 }),
    .c(2'b00),
    .d({open_n4631,1'b1}),
    .fci(\u2_Display/add120/c31 ),
    .f({open_n4648,\u2_Display/n3893 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u3_al_u4097  (
    .a({\u2_Display/n3885 ,\u2_Display/n3887 }),
    .b({\u2_Display/n3884 ,\u2_Display/n3886 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add120/c3 ),
    .f({\u2_Display/n3893 [5],\u2_Display/n3893 [3]}),
    .fco(\u2_Display/add120/c7 ),
    .fx({\u2_Display/n3893 [6],\u2_Display/n3893 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/u7_al_u4098  (
    .a({\u2_Display/n3881 ,\u2_Display/n3883 }),
    .b({\u2_Display/n3880 ,\u2_Display/n3882 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add120/c7 ),
    .f({\u2_Display/n3893 [9],\u2_Display/n3893 [7]}),
    .fco(\u2_Display/add120/c11 ),
    .fx({\u2_Display/n3893 [10],\u2_Display/n3893 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add120/ucin_al_u4096"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add120/ucin_al_u4096  (
    .a({\u2_Display/n3889 ,1'b1}),
    .b({\u2_Display/n3888 ,\u2_Display/n3890 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3893 [1],open_n4707}),
    .fco(\u2_Display/add120/c3 ),
    .fx({\u2_Display/n3893 [2],\u2_Display/n3893 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u11_al_u4108  (
    .a({\u2_Display/n3912 ,\u2_Display/n3914 }),
    .b({\u2_Display/n3911 ,\u2_Display/n3913 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add121/c11 ),
    .f({\u2_Display/n3928 [13],\u2_Display/n3928 [11]}),
    .fco(\u2_Display/add121/c15 ),
    .fx({\u2_Display/n3928 [14],\u2_Display/n3928 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u15_al_u4109  (
    .a({\u2_Display/n3908 ,\u2_Display/n3910 }),
    .b({\u2_Display/n3907 ,\u2_Display/n3909 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add121/c15 ),
    .f({\u2_Display/n3928 [17],\u2_Display/n3928 [15]}),
    .fco(\u2_Display/add121/c19 ),
    .fx({\u2_Display/n3928 [18],\u2_Display/n3928 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u19_al_u4110  (
    .a({\u2_Display/n3904 ,\u2_Display/n3906 }),
    .b({\u2_Display/n3903 ,\u2_Display/n3905 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add121/c19 ),
    .f({\u2_Display/n3928 [21],\u2_Display/n3928 [19]}),
    .fco(\u2_Display/add121/c23 ),
    .fx({\u2_Display/n3928 [22],\u2_Display/n3928 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u23_al_u4111  (
    .a({\u2_Display/n3900 ,\u2_Display/n3902 }),
    .b({\u2_Display/n3899 ,\u2_Display/n3901 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add121/c23 ),
    .f({\u2_Display/n3928 [25],\u2_Display/n3928 [23]}),
    .fco(\u2_Display/add121/c27 ),
    .fx({\u2_Display/n3928 [26],\u2_Display/n3928 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u27_al_u4112  (
    .a({\u2_Display/n3896 ,\u2_Display/n3898 }),
    .b({\u2_Display/n3895 ,\u2_Display/n3897 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add121/c27 ),
    .f({\u2_Display/n3928 [29],\u2_Display/n3928 [27]}),
    .fco(\u2_Display/add121/c31 ),
    .fx({\u2_Display/n3928 [30],\u2_Display/n3928 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u31_al_u4113  (
    .a({open_n4800,\u2_Display/n3894 }),
    .c(2'b00),
    .d({open_n4805,1'b1}),
    .fci(\u2_Display/add121/c31 ),
    .f({open_n4822,\u2_Display/n3928 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u3_al_u4106  (
    .a({\u2_Display/n3920 ,\u2_Display/n3922 }),
    .b({\u2_Display/n3919 ,\u2_Display/n3921 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add121/c3 ),
    .f({\u2_Display/n3928 [5],\u2_Display/n3928 [3]}),
    .fco(\u2_Display/add121/c7 ),
    .fx({\u2_Display/n3928 [6],\u2_Display/n3928 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/u7_al_u4107  (
    .a({\u2_Display/n3916 ,\u2_Display/n3918 }),
    .b({\u2_Display/n3915 ,\u2_Display/n3917 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add121/c7 ),
    .f({\u2_Display/n3928 [9],\u2_Display/n3928 [7]}),
    .fco(\u2_Display/add121/c11 ),
    .fx({\u2_Display/n3928 [10],\u2_Display/n3928 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add121/ucin_al_u4105"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add121/ucin_al_u4105  (
    .a({\u2_Display/n3924 ,1'b1}),
    .b({\u2_Display/n3923 ,\u2_Display/n3925 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3928 [1],open_n4881}),
    .fco(\u2_Display/add121/c3 ),
    .fx({\u2_Display/n3928 [2],\u2_Display/n3928 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u11_al_u4117  (
    .a({\u2_Display/n3947 ,\u2_Display/n3949 }),
    .b({\u2_Display/n3946 ,\u2_Display/n3948 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add122/c11 ),
    .f({\u2_Display/n3963 [13],\u2_Display/n3963 [11]}),
    .fco(\u2_Display/add122/c15 ),
    .fx({\u2_Display/n3963 [14],\u2_Display/n3963 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u15_al_u4118  (
    .a({\u2_Display/n3943 ,\u2_Display/n3945 }),
    .b({\u2_Display/n3942 ,\u2_Display/n3944 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add122/c15 ),
    .f({\u2_Display/n3963 [17],\u2_Display/n3963 [15]}),
    .fco(\u2_Display/add122/c19 ),
    .fx({\u2_Display/n3963 [18],\u2_Display/n3963 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u19_al_u4119  (
    .a({\u2_Display/n3939 ,\u2_Display/n3941 }),
    .b({\u2_Display/n3938 ,\u2_Display/n3940 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add122/c19 ),
    .f({\u2_Display/n3963 [21],\u2_Display/n3963 [19]}),
    .fco(\u2_Display/add122/c23 ),
    .fx({\u2_Display/n3963 [22],\u2_Display/n3963 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u23_al_u4120  (
    .a({\u2_Display/n3935 ,\u2_Display/n3937 }),
    .b({\u2_Display/n3934 ,\u2_Display/n3936 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add122/c23 ),
    .f({\u2_Display/n3963 [25],\u2_Display/n3963 [23]}),
    .fco(\u2_Display/add122/c27 ),
    .fx({\u2_Display/n3963 [26],\u2_Display/n3963 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u27_al_u4121  (
    .a({\u2_Display/n3931 ,\u2_Display/n3933 }),
    .b({\u2_Display/n3930 ,\u2_Display/n3932 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add122/c27 ),
    .f({\u2_Display/n3963 [29],\u2_Display/n3963 [27]}),
    .fco(\u2_Display/add122/c31 ),
    .fx({\u2_Display/n3963 [30],\u2_Display/n3963 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u31_al_u4122  (
    .a({open_n4974,\u2_Display/n3929 }),
    .c(2'b00),
    .d({open_n4979,1'b1}),
    .fci(\u2_Display/add122/c31 ),
    .f({open_n4996,\u2_Display/n3963 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u3_al_u4115  (
    .a({\u2_Display/n3955 ,\u2_Display/n3957 }),
    .b({\u2_Display/n3954 ,\u2_Display/n3956 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add122/c3 ),
    .f({\u2_Display/n3963 [5],\u2_Display/n3963 [3]}),
    .fco(\u2_Display/add122/c7 ),
    .fx({\u2_Display/n3963 [6],\u2_Display/n3963 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/u7_al_u4116  (
    .a({\u2_Display/n3951 ,\u2_Display/n3953 }),
    .b({\u2_Display/n3950 ,\u2_Display/n3952 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add122/c7 ),
    .f({\u2_Display/n3963 [9],\u2_Display/n3963 [7]}),
    .fco(\u2_Display/add122/c11 ),
    .fx({\u2_Display/n3963 [10],\u2_Display/n3963 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add122/ucin_al_u4114"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add122/ucin_al_u4114  (
    .a({\u2_Display/n3959 ,1'b1}),
    .b({\u2_Display/n3958 ,\u2_Display/n3960 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3963 [1],open_n5055}),
    .fco(\u2_Display/add122/c3 ),
    .fx({\u2_Display/n3963 [2],\u2_Display/n3963 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u11_al_u4126  (
    .a({\u2_Display/n3982 ,\u2_Display/n3984 }),
    .b({\u2_Display/n3981 ,\u2_Display/n3983 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add123/c11 ),
    .f({\u2_Display/n3998 [13],\u2_Display/n3998 [11]}),
    .fco(\u2_Display/add123/c15 ),
    .fx({\u2_Display/n3998 [14],\u2_Display/n3998 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u15_al_u4127  (
    .a({\u2_Display/n3978 ,\u2_Display/n3980 }),
    .b({\u2_Display/n3977 ,\u2_Display/n3979 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add123/c15 ),
    .f({\u2_Display/n3998 [17],\u2_Display/n3998 [15]}),
    .fco(\u2_Display/add123/c19 ),
    .fx({\u2_Display/n3998 [18],\u2_Display/n3998 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u19_al_u4128  (
    .a({\u2_Display/n3974 ,\u2_Display/n3976 }),
    .b({\u2_Display/n3973 ,\u2_Display/n3975 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add123/c19 ),
    .f({\u2_Display/n3998 [21],\u2_Display/n3998 [19]}),
    .fco(\u2_Display/add123/c23 ),
    .fx({\u2_Display/n3998 [22],\u2_Display/n3998 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u23_al_u4129  (
    .a({\u2_Display/n3970 ,\u2_Display/n3972 }),
    .b({\u2_Display/n3969 ,\u2_Display/n3971 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add123/c23 ),
    .f({\u2_Display/n3998 [25],\u2_Display/n3998 [23]}),
    .fco(\u2_Display/add123/c27 ),
    .fx({\u2_Display/n3998 [26],\u2_Display/n3998 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u27_al_u4130  (
    .a({\u2_Display/n3966 ,\u2_Display/n3968 }),
    .b({\u2_Display/n3965 ,\u2_Display/n3967 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add123/c27 ),
    .f({\u2_Display/n3998 [29],\u2_Display/n3998 [27]}),
    .fco(\u2_Display/add123/c31 ),
    .fx({\u2_Display/n3998 [30],\u2_Display/n3998 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u31_al_u4131  (
    .a({open_n5148,\u2_Display/n3964 }),
    .c(2'b00),
    .d({open_n5153,1'b1}),
    .fci(\u2_Display/add123/c31 ),
    .f({open_n5170,\u2_Display/n3998 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u3_al_u4124  (
    .a({\u2_Display/n3990 ,\u2_Display/n3992 }),
    .b({\u2_Display/n3989 ,\u2_Display/n3991 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add123/c3 ),
    .f({\u2_Display/n3998 [5],\u2_Display/n3998 [3]}),
    .fco(\u2_Display/add123/c7 ),
    .fx({\u2_Display/n3998 [6],\u2_Display/n3998 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/u7_al_u4125  (
    .a({\u2_Display/n3986 ,\u2_Display/n3988 }),
    .b({\u2_Display/n3985 ,\u2_Display/n3987 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add123/c7 ),
    .f({\u2_Display/n3998 [9],\u2_Display/n3998 [7]}),
    .fco(\u2_Display/add123/c11 ),
    .fx({\u2_Display/n3998 [10],\u2_Display/n3998 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add123/ucin_al_u4123"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add123/ucin_al_u4123  (
    .a({\u2_Display/n3994 ,1'b1}),
    .b({\u2_Display/n3993 ,\u2_Display/n3995 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3998 [1],open_n5229}),
    .fco(\u2_Display/add123/c3 ),
    .fx({\u2_Display/n3998 [2],\u2_Display/n3998 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u11_al_u4135  (
    .a({\u2_Display/n4017 ,\u2_Display/n4019 }),
    .b({\u2_Display/n4016 ,\u2_Display/n4018 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add124/c11 ),
    .f({\u2_Display/n4033 [13],\u2_Display/n4033 [11]}),
    .fco(\u2_Display/add124/c15 ),
    .fx({\u2_Display/n4033 [14],\u2_Display/n4033 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u15_al_u4136  (
    .a({\u2_Display/n4013 ,\u2_Display/n4015 }),
    .b({\u2_Display/n4012 ,\u2_Display/n4014 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add124/c15 ),
    .f({\u2_Display/n4033 [17],\u2_Display/n4033 [15]}),
    .fco(\u2_Display/add124/c19 ),
    .fx({\u2_Display/n4033 [18],\u2_Display/n4033 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u19_al_u4137  (
    .a({\u2_Display/n4009 ,\u2_Display/n4011 }),
    .b({\u2_Display/n4008 ,\u2_Display/n4010 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add124/c19 ),
    .f({\u2_Display/n4033 [21],\u2_Display/n4033 [19]}),
    .fco(\u2_Display/add124/c23 ),
    .fx({\u2_Display/n4033 [22],\u2_Display/n4033 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u23_al_u4138  (
    .a({\u2_Display/n4005 ,\u2_Display/n4007 }),
    .b({\u2_Display/n4004 ,\u2_Display/n4006 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add124/c23 ),
    .f({\u2_Display/n4033 [25],\u2_Display/n4033 [23]}),
    .fco(\u2_Display/add124/c27 ),
    .fx({\u2_Display/n4033 [26],\u2_Display/n4033 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u27_al_u4139  (
    .a({\u2_Display/n4001 ,\u2_Display/n4003 }),
    .b({\u2_Display/n4000 ,\u2_Display/n4002 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add124/c27 ),
    .f({\u2_Display/n4033 [29],\u2_Display/n4033 [27]}),
    .fco(\u2_Display/add124/c31 ),
    .fx({\u2_Display/n4033 [30],\u2_Display/n4033 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u31_al_u4140  (
    .a({open_n5322,\u2_Display/n3999 }),
    .c(2'b00),
    .d({open_n5327,1'b1}),
    .fci(\u2_Display/add124/c31 ),
    .f({open_n5344,\u2_Display/n4033 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u3_al_u4133  (
    .a({\u2_Display/n4025 ,\u2_Display/n4027 }),
    .b({\u2_Display/n4024 ,\u2_Display/n4026 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add124/c3 ),
    .f({\u2_Display/n4033 [5],\u2_Display/n4033 [3]}),
    .fco(\u2_Display/add124/c7 ),
    .fx({\u2_Display/n4033 [6],\u2_Display/n4033 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/u7_al_u4134  (
    .a({\u2_Display/n4021 ,\u2_Display/n4023 }),
    .b({\u2_Display/n4020 ,\u2_Display/n4022 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add124/c7 ),
    .f({\u2_Display/n4033 [9],\u2_Display/n4033 [7]}),
    .fco(\u2_Display/add124/c11 ),
    .fx({\u2_Display/n4033 [10],\u2_Display/n4033 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add124/ucin_al_u4132"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add124/ucin_al_u4132  (
    .a({\u2_Display/n4029 ,1'b1}),
    .b({\u2_Display/n4028 ,\u2_Display/n4030 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4033 [1],open_n5403}),
    .fco(\u2_Display/add124/c3 ),
    .fx({\u2_Display/n4033 [2],\u2_Display/n4033 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u11_al_u4144  (
    .a({\u2_Display/n4052 ,\u2_Display/n4054 }),
    .b({\u2_Display/n4051 ,\u2_Display/n4053 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add125/c11 ),
    .f({\u2_Display/n4068 [13],\u2_Display/n4068 [11]}),
    .fco(\u2_Display/add125/c15 ),
    .fx({\u2_Display/n4068 [14],\u2_Display/n4068 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u15_al_u4145  (
    .a({\u2_Display/n4048 ,\u2_Display/n4050 }),
    .b({\u2_Display/n4047 ,\u2_Display/n4049 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add125/c15 ),
    .f({\u2_Display/n4068 [17],\u2_Display/n4068 [15]}),
    .fco(\u2_Display/add125/c19 ),
    .fx({\u2_Display/n4068 [18],\u2_Display/n4068 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u19_al_u4146  (
    .a({\u2_Display/n4044 ,\u2_Display/n4046 }),
    .b({\u2_Display/n4043 ,\u2_Display/n4045 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add125/c19 ),
    .f({\u2_Display/n4068 [21],\u2_Display/n4068 [19]}),
    .fco(\u2_Display/add125/c23 ),
    .fx({\u2_Display/n4068 [22],\u2_Display/n4068 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u23_al_u4147  (
    .a({\u2_Display/n4040 ,\u2_Display/n4042 }),
    .b({\u2_Display/n4039 ,\u2_Display/n4041 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add125/c23 ),
    .f({\u2_Display/n4068 [25],\u2_Display/n4068 [23]}),
    .fco(\u2_Display/add125/c27 ),
    .fx({\u2_Display/n4068 [26],\u2_Display/n4068 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u27_al_u4148  (
    .a({\u2_Display/n4036 ,\u2_Display/n4038 }),
    .b({\u2_Display/n4035 ,\u2_Display/n4037 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add125/c27 ),
    .f({\u2_Display/n4068 [29],\u2_Display/n4068 [27]}),
    .fco(\u2_Display/add125/c31 ),
    .fx({\u2_Display/n4068 [30],\u2_Display/n4068 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u31_al_u4149  (
    .a({open_n5496,\u2_Display/n4034 }),
    .c(2'b00),
    .d({open_n5501,1'b1}),
    .fci(\u2_Display/add125/c31 ),
    .f({open_n5518,\u2_Display/n4068 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u3_al_u4142  (
    .a({\u2_Display/n4060 ,\u2_Display/n4062 }),
    .b({\u2_Display/n4059 ,\u2_Display/n4061 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add125/c3 ),
    .f({\u2_Display/n4068 [5],\u2_Display/n4068 [3]}),
    .fco(\u2_Display/add125/c7 ),
    .fx({\u2_Display/n4068 [6],\u2_Display/n4068 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/u7_al_u4143  (
    .a({\u2_Display/n4056 ,\u2_Display/n4058 }),
    .b({\u2_Display/n4055 ,\u2_Display/n4057 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add125/c7 ),
    .f({\u2_Display/n4068 [9],\u2_Display/n4068 [7]}),
    .fco(\u2_Display/add125/c11 ),
    .fx({\u2_Display/n4068 [10],\u2_Display/n4068 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add125/ucin_al_u4141"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add125/ucin_al_u4141  (
    .a({\u2_Display/n4064 ,1'b1}),
    .b({\u2_Display/n4063 ,\u2_Display/n4065 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4068 [1],open_n5577}),
    .fco(\u2_Display/add125/c3 ),
    .fx({\u2_Display/n4068 [2],\u2_Display/n4068 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u11_al_u4153  (
    .a({\u2_Display/n4087 ,\u2_Display/n4089 }),
    .b({\u2_Display/n4086 ,\u2_Display/n4088 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add126/c11 ),
    .f({\u2_Display/n4103 [13],\u2_Display/n4103 [11]}),
    .fco(\u2_Display/add126/c15 ),
    .fx({\u2_Display/n4103 [14],\u2_Display/n4103 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u15_al_u4154  (
    .a({\u2_Display/n4083 ,\u2_Display/n4085 }),
    .b({\u2_Display/n4082 ,\u2_Display/n4084 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add126/c15 ),
    .f({\u2_Display/n4103 [17],\u2_Display/n4103 [15]}),
    .fco(\u2_Display/add126/c19 ),
    .fx({\u2_Display/n4103 [18],\u2_Display/n4103 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u19_al_u4155  (
    .a({\u2_Display/n4079 ,\u2_Display/n4081 }),
    .b({\u2_Display/n4078 ,\u2_Display/n4080 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add126/c19 ),
    .f({\u2_Display/n4103 [21],\u2_Display/n4103 [19]}),
    .fco(\u2_Display/add126/c23 ),
    .fx({\u2_Display/n4103 [22],\u2_Display/n4103 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u23_al_u4156  (
    .a({\u2_Display/n4075 ,\u2_Display/n4077 }),
    .b({\u2_Display/n4074 ,\u2_Display/n4076 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add126/c23 ),
    .f({\u2_Display/n4103 [25],\u2_Display/n4103 [23]}),
    .fco(\u2_Display/add126/c27 ),
    .fx({\u2_Display/n4103 [26],\u2_Display/n4103 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u27_al_u4157  (
    .a({\u2_Display/n4071 ,\u2_Display/n4073 }),
    .b({\u2_Display/n4070 ,\u2_Display/n4072 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add126/c27 ),
    .f({\u2_Display/n4103 [29],\u2_Display/n4103 [27]}),
    .fco(\u2_Display/add126/c31 ),
    .fx({\u2_Display/n4103 [30],\u2_Display/n4103 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u31_al_u4158  (
    .a({open_n5670,\u2_Display/n4069 }),
    .c(2'b00),
    .d({open_n5675,1'b1}),
    .fci(\u2_Display/add126/c31 ),
    .f({open_n5692,\u2_Display/n4103 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u3_al_u4151  (
    .a({\u2_Display/n4095 ,\u2_Display/n4097 }),
    .b({\u2_Display/n4094 ,\u2_Display/n4096 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add126/c3 ),
    .f({\u2_Display/n4103 [5],\u2_Display/n4103 [3]}),
    .fco(\u2_Display/add126/c7 ),
    .fx({\u2_Display/n4103 [6],\u2_Display/n4103 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/u7_al_u4152  (
    .a({\u2_Display/n4091 ,\u2_Display/n4093 }),
    .b({\u2_Display/n4090 ,\u2_Display/n4092 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add126/c7 ),
    .f({\u2_Display/n4103 [9],\u2_Display/n4103 [7]}),
    .fco(\u2_Display/add126/c11 ),
    .fx({\u2_Display/n4103 [10],\u2_Display/n4103 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add126/ucin_al_u4150"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add126/ucin_al_u4150  (
    .a({\u2_Display/n4099 ,1'b1}),
    .b({\u2_Display/n4098 ,\u2_Display/n4100 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4103 [1],open_n5751}),
    .fco(\u2_Display/add126/c3 ),
    .fx({\u2_Display/n4103 [2],\u2_Display/n4103 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u11_al_u4162  (
    .a({\u2_Display/n4122 ,\u2_Display/n4124 }),
    .b({\u2_Display/n4121 ,\u2_Display/n4123 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add127/c11 ),
    .f({\u2_Display/n4138 [13],\u2_Display/n4138 [11]}),
    .fco(\u2_Display/add127/c15 ),
    .fx({\u2_Display/n4138 [14],\u2_Display/n4138 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u15_al_u4163  (
    .a({\u2_Display/n4118 ,\u2_Display/n4120 }),
    .b({\u2_Display/n4117 ,\u2_Display/n4119 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add127/c15 ),
    .f({\u2_Display/n4138 [17],\u2_Display/n4138 [15]}),
    .fco(\u2_Display/add127/c19 ),
    .fx({\u2_Display/n4138 [18],\u2_Display/n4138 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u19_al_u4164  (
    .a({\u2_Display/n4114 ,\u2_Display/n4116 }),
    .b({\u2_Display/n4113 ,\u2_Display/n4115 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add127/c19 ),
    .f({\u2_Display/n4138 [21],\u2_Display/n4138 [19]}),
    .fco(\u2_Display/add127/c23 ),
    .fx({\u2_Display/n4138 [22],\u2_Display/n4138 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u23_al_u4165  (
    .a({\u2_Display/n4110 ,\u2_Display/n4112 }),
    .b({\u2_Display/n4109 ,\u2_Display/n4111 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add127/c23 ),
    .f({\u2_Display/n4138 [25],\u2_Display/n4138 [23]}),
    .fco(\u2_Display/add127/c27 ),
    .fx({\u2_Display/n4138 [26],\u2_Display/n4138 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u27_al_u4166  (
    .a({\u2_Display/n4106 ,\u2_Display/n4108 }),
    .b({\u2_Display/n4105 ,\u2_Display/n4107 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add127/c27 ),
    .f({\u2_Display/n4138 [29],\u2_Display/n4138 [27]}),
    .fco(\u2_Display/add127/c31 ),
    .fx({\u2_Display/n4138 [30],\u2_Display/n4138 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u31_al_u4167  (
    .a({open_n5844,\u2_Display/n4104 }),
    .c(2'b00),
    .d({open_n5849,1'b1}),
    .fci(\u2_Display/add127/c31 ),
    .f({open_n5866,\u2_Display/n4138 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u3_al_u4160  (
    .a({\u2_Display/n4130 ,\u2_Display/n4132 }),
    .b({\u2_Display/n4129 ,\u2_Display/n4131 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add127/c3 ),
    .f({\u2_Display/n4138 [5],\u2_Display/n4138 [3]}),
    .fco(\u2_Display/add127/c7 ),
    .fx({\u2_Display/n4138 [6],\u2_Display/n4138 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/u7_al_u4161  (
    .a({\u2_Display/n4126 ,\u2_Display/n4128 }),
    .b({\u2_Display/n4125 ,\u2_Display/n4127 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add127/c7 ),
    .f({\u2_Display/n4138 [9],\u2_Display/n4138 [7]}),
    .fco(\u2_Display/add127/c11 ),
    .fx({\u2_Display/n4138 [10],\u2_Display/n4138 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add127/ucin_al_u4159"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add127/ucin_al_u4159  (
    .a({\u2_Display/n4134 ,1'b1}),
    .b({\u2_Display/n4133 ,\u2_Display/n4135 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4138 [1],open_n5925}),
    .fco(\u2_Display/add127/c3 ),
    .fx({\u2_Display/n4138 [2],\u2_Display/n4138 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u11_al_u4171  (
    .a({\u2_Display/n4157 ,\u2_Display/n4159 }),
    .b({\u2_Display/n4156 ,\u2_Display/n4158 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add128/c11 ),
    .f({\u2_Display/n4173 [13],\u2_Display/n4173 [11]}),
    .fco(\u2_Display/add128/c15 ),
    .fx({\u2_Display/n4173 [14],\u2_Display/n4173 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u15_al_u4172  (
    .a({\u2_Display/n4153 ,\u2_Display/n4155 }),
    .b({\u2_Display/n4152 ,\u2_Display/n4154 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add128/c15 ),
    .f({\u2_Display/n4173 [17],\u2_Display/n4173 [15]}),
    .fco(\u2_Display/add128/c19 ),
    .fx({\u2_Display/n4173 [18],\u2_Display/n4173 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u19_al_u4173  (
    .a({\u2_Display/n4149 ,\u2_Display/n4151 }),
    .b({\u2_Display/n4148 ,\u2_Display/n4150 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add128/c19 ),
    .f({\u2_Display/n4173 [21],\u2_Display/n4173 [19]}),
    .fco(\u2_Display/add128/c23 ),
    .fx({\u2_Display/n4173 [22],\u2_Display/n4173 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u23_al_u4174  (
    .a({\u2_Display/n4145 ,\u2_Display/n4147 }),
    .b({\u2_Display/n4144 ,\u2_Display/n4146 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add128/c23 ),
    .f({\u2_Display/n4173 [25],\u2_Display/n4173 [23]}),
    .fco(\u2_Display/add128/c27 ),
    .fx({\u2_Display/n4173 [26],\u2_Display/n4173 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u27_al_u4175  (
    .a({\u2_Display/n4141 ,\u2_Display/n4143 }),
    .b({\u2_Display/n4140 ,\u2_Display/n4142 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add128/c27 ),
    .f({\u2_Display/n4173 [29],\u2_Display/n4173 [27]}),
    .fco(\u2_Display/add128/c31 ),
    .fx({\u2_Display/n4173 [30],\u2_Display/n4173 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u31_al_u4176  (
    .a({open_n6018,\u2_Display/n4139 }),
    .c(2'b00),
    .d({open_n6023,1'b1}),
    .fci(\u2_Display/add128/c31 ),
    .f({open_n6040,\u2_Display/n4173 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u3_al_u4169  (
    .a({\u2_Display/n4165 ,\u2_Display/n4167 }),
    .b({\u2_Display/n4164 ,\u2_Display/n4166 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add128/c3 ),
    .f({\u2_Display/n4173 [5],\u2_Display/n4173 [3]}),
    .fco(\u2_Display/add128/c7 ),
    .fx({\u2_Display/n4173 [6],\u2_Display/n4173 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/u7_al_u4170  (
    .a({\u2_Display/n4161 ,\u2_Display/n4163 }),
    .b({\u2_Display/n4160 ,\u2_Display/n4162 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add128/c7 ),
    .f({\u2_Display/n4173 [9],\u2_Display/n4173 [7]}),
    .fco(\u2_Display/add128/c11 ),
    .fx({\u2_Display/n4173 [10],\u2_Display/n4173 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add128/ucin_al_u4168"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add128/ucin_al_u4168  (
    .a({\u2_Display/n4169 ,1'b1}),
    .b({\u2_Display/n4168 ,\u2_Display/n4170 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4173 [1],open_n6099}),
    .fco(\u2_Display/add128/c3 ),
    .fx({\u2_Display/n4173 [2],\u2_Display/n4173 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u11_al_u4180  (
    .a({\u2_Display/n4192 ,\u2_Display/n4194 }),
    .b({\u2_Display/n4191 ,\u2_Display/n4193 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add129/c11 ),
    .f({\u2_Display/n4208 [13],\u2_Display/n4208 [11]}),
    .fco(\u2_Display/add129/c15 ),
    .fx({\u2_Display/n4208 [14],\u2_Display/n4208 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u15_al_u4181  (
    .a({\u2_Display/n4188 ,\u2_Display/n4190 }),
    .b({\u2_Display/n4187 ,\u2_Display/n4189 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add129/c15 ),
    .f({\u2_Display/n4208 [17],\u2_Display/n4208 [15]}),
    .fco(\u2_Display/add129/c19 ),
    .fx({\u2_Display/n4208 [18],\u2_Display/n4208 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u19_al_u4182  (
    .a({\u2_Display/n4184 ,\u2_Display/n4186 }),
    .b({\u2_Display/n4183 ,\u2_Display/n4185 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add129/c19 ),
    .f({\u2_Display/n4208 [21],\u2_Display/n4208 [19]}),
    .fco(\u2_Display/add129/c23 ),
    .fx({\u2_Display/n4208 [22],\u2_Display/n4208 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u23_al_u4183  (
    .a({\u2_Display/n4180 ,\u2_Display/n4182 }),
    .b({\u2_Display/n4179 ,\u2_Display/n4181 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add129/c23 ),
    .f({\u2_Display/n4208 [25],\u2_Display/n4208 [23]}),
    .fco(\u2_Display/add129/c27 ),
    .fx({\u2_Display/n4208 [26],\u2_Display/n4208 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u27_al_u4184  (
    .a({\u2_Display/n4176 ,\u2_Display/n4178 }),
    .b({\u2_Display/n4175 ,\u2_Display/n4177 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add129/c27 ),
    .f({\u2_Display/n4208 [29],\u2_Display/n4208 [27]}),
    .fco(\u2_Display/add129/c31 ),
    .fx({\u2_Display/n4208 [30],\u2_Display/n4208 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u31_al_u4185  (
    .a({open_n6192,\u2_Display/n4174 }),
    .c(2'b00),
    .d({open_n6197,1'b1}),
    .fci(\u2_Display/add129/c31 ),
    .f({open_n6214,\u2_Display/n4208 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u3_al_u4178  (
    .a({\u2_Display/n4200 ,\u2_Display/n4202 }),
    .b({\u2_Display/n4199 ,\u2_Display/n4201 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add129/c3 ),
    .f({\u2_Display/n4208 [5],\u2_Display/n4208 [3]}),
    .fco(\u2_Display/add129/c7 ),
    .fx({\u2_Display/n4208 [6],\u2_Display/n4208 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/u7_al_u4179  (
    .a({\u2_Display/n4196 ,\u2_Display/n4198 }),
    .b({\u2_Display/n4195 ,\u2_Display/n4197 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add129/c7 ),
    .f({\u2_Display/n4208 [9],\u2_Display/n4208 [7]}),
    .fco(\u2_Display/add129/c11 ),
    .fx({\u2_Display/n4208 [10],\u2_Display/n4208 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add129/ucin_al_u4177"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add129/ucin_al_u4177  (
    .a({\u2_Display/n4204 ,1'b1}),
    .b({\u2_Display/n4203 ,\u2_Display/n4205 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4208 [1],open_n6273}),
    .fco(\u2_Display/add129/c3 ),
    .fx({\u2_Display/n4208 [2],\u2_Display/n4208 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u11_al_u4189  (
    .a({\u2_Display/n4227 ,\u2_Display/n4229 }),
    .b({\u2_Display/n4226 ,\u2_Display/n4228 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add130/c11 ),
    .f({\u2_Display/n4243 [13],\u2_Display/n4243 [11]}),
    .fco(\u2_Display/add130/c15 ),
    .fx({\u2_Display/n4243 [14],\u2_Display/n4243 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u15_al_u4190  (
    .a({\u2_Display/n4223 ,\u2_Display/n4225 }),
    .b({\u2_Display/n4222 ,\u2_Display/n4224 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add130/c15 ),
    .f({\u2_Display/n4243 [17],\u2_Display/n4243 [15]}),
    .fco(\u2_Display/add130/c19 ),
    .fx({\u2_Display/n4243 [18],\u2_Display/n4243 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u19_al_u4191  (
    .a({\u2_Display/n4219 ,\u2_Display/n4221 }),
    .b({\u2_Display/n4218 ,\u2_Display/n4220 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add130/c19 ),
    .f({\u2_Display/n4243 [21],\u2_Display/n4243 [19]}),
    .fco(\u2_Display/add130/c23 ),
    .fx({\u2_Display/n4243 [22],\u2_Display/n4243 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u23_al_u4192  (
    .a({\u2_Display/n4215 ,\u2_Display/n4217 }),
    .b({\u2_Display/n4214 ,\u2_Display/n4216 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add130/c23 ),
    .f({\u2_Display/n4243 [25],\u2_Display/n4243 [23]}),
    .fco(\u2_Display/add130/c27 ),
    .fx({\u2_Display/n4243 [26],\u2_Display/n4243 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u27_al_u4193  (
    .a({\u2_Display/n4211 ,\u2_Display/n4213 }),
    .b({\u2_Display/n4210 ,\u2_Display/n4212 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add130/c27 ),
    .f({\u2_Display/n4243 [29],\u2_Display/n4243 [27]}),
    .fco(\u2_Display/add130/c31 ),
    .fx({\u2_Display/n4243 [30],\u2_Display/n4243 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u31_al_u4194  (
    .a({open_n6366,\u2_Display/n4209 }),
    .c(2'b00),
    .d({open_n6371,1'b1}),
    .fci(\u2_Display/add130/c31 ),
    .f({open_n6388,\u2_Display/n4243 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u3_al_u4187  (
    .a({\u2_Display/n4235 ,\u2_Display/n4237 }),
    .b({\u2_Display/n4234 ,\u2_Display/n4236 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add130/c3 ),
    .f({\u2_Display/n4243 [5],\u2_Display/n4243 [3]}),
    .fco(\u2_Display/add130/c7 ),
    .fx({\u2_Display/n4243 [6],\u2_Display/n4243 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/u7_al_u4188  (
    .a({\u2_Display/n4231 ,\u2_Display/n4233 }),
    .b({\u2_Display/n4230 ,\u2_Display/n4232 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add130/c7 ),
    .f({\u2_Display/n4243 [9],\u2_Display/n4243 [7]}),
    .fco(\u2_Display/add130/c11 ),
    .fx({\u2_Display/n4243 [10],\u2_Display/n4243 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add130/ucin_al_u4186"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add130/ucin_al_u4186  (
    .a({\u2_Display/n4239 ,1'b1}),
    .b({\u2_Display/n4238 ,\u2_Display/n4240 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4243 [1],open_n6447}),
    .fco(\u2_Display/add130/c3 ),
    .fx({\u2_Display/n4243 [2],\u2_Display/n4243 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u11_al_u4198  (
    .a({\u2_Display/n4262 ,\u2_Display/n4264 }),
    .b({\u2_Display/n4261 ,\u2_Display/n4263 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add131/c11 ),
    .f({\u2_Display/n4278 [13],\u2_Display/n4278 [11]}),
    .fco(\u2_Display/add131/c15 ),
    .fx({\u2_Display/n4278 [14],\u2_Display/n4278 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u15_al_u4199  (
    .a({\u2_Display/n4258 ,\u2_Display/n4260 }),
    .b({\u2_Display/n4257 ,\u2_Display/n4259 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add131/c15 ),
    .f({\u2_Display/n4278 [17],\u2_Display/n4278 [15]}),
    .fco(\u2_Display/add131/c19 ),
    .fx({\u2_Display/n4278 [18],\u2_Display/n4278 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u19_al_u4200  (
    .a({\u2_Display/n4254 ,\u2_Display/n4256 }),
    .b({\u2_Display/n4253 ,\u2_Display/n4255 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add131/c19 ),
    .f({\u2_Display/n4278 [21],\u2_Display/n4278 [19]}),
    .fco(\u2_Display/add131/c23 ),
    .fx({\u2_Display/n4278 [22],\u2_Display/n4278 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u23_al_u4201  (
    .a({\u2_Display/n4250 ,\u2_Display/n4252 }),
    .b({\u2_Display/n4249 ,\u2_Display/n4251 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add131/c23 ),
    .f({\u2_Display/n4278 [25],\u2_Display/n4278 [23]}),
    .fco(\u2_Display/add131/c27 ),
    .fx({\u2_Display/n4278 [26],\u2_Display/n4278 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u27_al_u4202  (
    .a({\u2_Display/n4246 ,\u2_Display/n4248 }),
    .b({\u2_Display/n4245 ,\u2_Display/n4247 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add131/c27 ),
    .f({\u2_Display/n4278 [29],\u2_Display/n4278 [27]}),
    .fco(\u2_Display/add131/c31 ),
    .fx({\u2_Display/n4278 [30],\u2_Display/n4278 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u31_al_u4203  (
    .a({open_n6540,\u2_Display/n4244 }),
    .c(2'b00),
    .d({open_n6545,1'b1}),
    .fci(\u2_Display/add131/c31 ),
    .f({open_n6562,\u2_Display/n4278 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u3_al_u4196  (
    .a({\u2_Display/n4270 ,\u2_Display/n4272 }),
    .b({\u2_Display/n4269 ,\u2_Display/n4271 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add131/c3 ),
    .f({\u2_Display/n4278 [5],\u2_Display/n4278 [3]}),
    .fco(\u2_Display/add131/c7 ),
    .fx({\u2_Display/n4278 [6],\u2_Display/n4278 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/u7_al_u4197  (
    .a({\u2_Display/n4266 ,\u2_Display/n4268 }),
    .b({\u2_Display/n4265 ,\u2_Display/n4267 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add131/c7 ),
    .f({\u2_Display/n4278 [9],\u2_Display/n4278 [7]}),
    .fco(\u2_Display/add131/c11 ),
    .fx({\u2_Display/n4278 [10],\u2_Display/n4278 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add131/ucin_al_u4195"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add131/ucin_al_u4195  (
    .a({\u2_Display/n4274 ,1'b1}),
    .b({\u2_Display/n4273 ,\u2_Display/n4275 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4278 [1],open_n6621}),
    .fco(\u2_Display/add131/c3 ),
    .fx({\u2_Display/n4278 [2],\u2_Display/n4278 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u11_al_u4207  (
    .a({\u2_Display/n4297 ,\u2_Display/n4299 }),
    .b({\u2_Display/n4296 ,\u2_Display/n4298 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add132/c11 ),
    .f({\u2_Display/n4313 [13],\u2_Display/n4313 [11]}),
    .fco(\u2_Display/add132/c15 ),
    .fx({\u2_Display/n4313 [14],\u2_Display/n4313 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u15_al_u4208  (
    .a({\u2_Display/n4293 ,\u2_Display/n4295 }),
    .b({\u2_Display/n4292 ,\u2_Display/n4294 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add132/c15 ),
    .f({\u2_Display/n4313 [17],\u2_Display/n4313 [15]}),
    .fco(\u2_Display/add132/c19 ),
    .fx({\u2_Display/n4313 [18],\u2_Display/n4313 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u19_al_u4209  (
    .a({\u2_Display/n4289 ,\u2_Display/n4291 }),
    .b({\u2_Display/n4288 ,\u2_Display/n4290 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add132/c19 ),
    .f({\u2_Display/n4313 [21],\u2_Display/n4313 [19]}),
    .fco(\u2_Display/add132/c23 ),
    .fx({\u2_Display/n4313 [22],\u2_Display/n4313 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u23_al_u4210  (
    .a({\u2_Display/n4285 ,\u2_Display/n4287 }),
    .b({\u2_Display/n4284 ,\u2_Display/n4286 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add132/c23 ),
    .f({\u2_Display/n4313 [25],\u2_Display/n4313 [23]}),
    .fco(\u2_Display/add132/c27 ),
    .fx({\u2_Display/n4313 [26],\u2_Display/n4313 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u27_al_u4211  (
    .a({\u2_Display/n4281 ,\u2_Display/n4283 }),
    .b({\u2_Display/n4280 ,\u2_Display/n4282 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add132/c27 ),
    .f({\u2_Display/n4313 [29],\u2_Display/n4313 [27]}),
    .fco(\u2_Display/add132/c31 ),
    .fx({\u2_Display/n4313 [30],\u2_Display/n4313 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u31_al_u4212  (
    .a({open_n6714,\u2_Display/n4279 }),
    .c(2'b00),
    .d({open_n6719,1'b1}),
    .fci(\u2_Display/add132/c31 ),
    .f({open_n6736,\u2_Display/n4313 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u3_al_u4205  (
    .a({\u2_Display/n4305 ,\u2_Display/n4307 }),
    .b({\u2_Display/n4304 ,\u2_Display/n4306 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add132/c3 ),
    .f({\u2_Display/n4313 [5],\u2_Display/n4313 [3]}),
    .fco(\u2_Display/add132/c7 ),
    .fx({\u2_Display/n4313 [6],\u2_Display/n4313 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/u7_al_u4206  (
    .a({\u2_Display/n4301 ,\u2_Display/n4303 }),
    .b({\u2_Display/n4300 ,\u2_Display/n4302 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add132/c7 ),
    .f({\u2_Display/n4313 [9],\u2_Display/n4313 [7]}),
    .fco(\u2_Display/add132/c11 ),
    .fx({\u2_Display/n4313 [10],\u2_Display/n4313 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add132/ucin_al_u4204"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add132/ucin_al_u4204  (
    .a({\u2_Display/n4309 ,1'b1}),
    .b({\u2_Display/n4308 ,\u2_Display/n4310 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4313 [1],open_n6795}),
    .fco(\u2_Display/add132/c3 ),
    .fx({\u2_Display/n4313 [2],\u2_Display/n4313 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u11_al_u4216  (
    .a({\u2_Display/n4332 ,\u2_Display/n4334 }),
    .b({\u2_Display/n4331 ,\u2_Display/n4333 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add133/c11 ),
    .f({\u2_Display/n4348 [13],\u2_Display/n4348 [11]}),
    .fco(\u2_Display/add133/c15 ),
    .fx({\u2_Display/n4348 [14],\u2_Display/n4348 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u15_al_u4217  (
    .a({\u2_Display/n4328 ,\u2_Display/n4330 }),
    .b({\u2_Display/n4327 ,\u2_Display/n4329 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add133/c15 ),
    .f({\u2_Display/n4348 [17],\u2_Display/n4348 [15]}),
    .fco(\u2_Display/add133/c19 ),
    .fx({\u2_Display/n4348 [18],\u2_Display/n4348 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u19_al_u4218  (
    .a({\u2_Display/n4324 ,\u2_Display/n4326 }),
    .b({\u2_Display/n4323 ,\u2_Display/n4325 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add133/c19 ),
    .f({\u2_Display/n4348 [21],\u2_Display/n4348 [19]}),
    .fco(\u2_Display/add133/c23 ),
    .fx({\u2_Display/n4348 [22],\u2_Display/n4348 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u23_al_u4219  (
    .a({\u2_Display/n4320 ,\u2_Display/n4322 }),
    .b({\u2_Display/n4319 ,\u2_Display/n4321 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add133/c23 ),
    .f({\u2_Display/n4348 [25],\u2_Display/n4348 [23]}),
    .fco(\u2_Display/add133/c27 ),
    .fx({\u2_Display/n4348 [26],\u2_Display/n4348 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u27_al_u4220  (
    .a({\u2_Display/n4316 ,\u2_Display/n4318 }),
    .b({\u2_Display/n4315 ,\u2_Display/n4317 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add133/c27 ),
    .f({\u2_Display/n4348 [29],\u2_Display/n4348 [27]}),
    .fco(\u2_Display/add133/c31 ),
    .fx({\u2_Display/n4348 [30],\u2_Display/n4348 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u31_al_u4221  (
    .a({open_n6888,\u2_Display/n4314 }),
    .c(2'b00),
    .d({open_n6893,1'b1}),
    .fci(\u2_Display/add133/c31 ),
    .f({open_n6910,\u2_Display/n4348 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u3_al_u4214  (
    .a({\u2_Display/n4340 ,\u2_Display/n4342 }),
    .b({\u2_Display/n4339 ,\u2_Display/n4341 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add133/c3 ),
    .f({\u2_Display/n4348 [5],\u2_Display/n4348 [3]}),
    .fco(\u2_Display/add133/c7 ),
    .fx({\u2_Display/n4348 [6],\u2_Display/n4348 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/u7_al_u4215  (
    .a({\u2_Display/n4336 ,\u2_Display/n4338 }),
    .b({\u2_Display/n4335 ,\u2_Display/n4337 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add133/c7 ),
    .f({\u2_Display/n4348 [9],\u2_Display/n4348 [7]}),
    .fco(\u2_Display/add133/c11 ),
    .fx({\u2_Display/n4348 [10],\u2_Display/n4348 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add133/ucin_al_u4213"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add133/ucin_al_u4213  (
    .a({\u2_Display/n4344 ,1'b1}),
    .b({\u2_Display/n4343 ,\u2_Display/n4345 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4348 [1],open_n6969}),
    .fco(\u2_Display/add133/c3 ),
    .fx({\u2_Display/n4348 [2],\u2_Display/n4348 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u11_al_u4225  (
    .a({\u2_Display/n4367 ,\u2_Display/n4369 }),
    .b({\u2_Display/n4366 ,\u2_Display/n4368 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add134/c11 ),
    .f({\u2_Display/n4383 [13],\u2_Display/n4383 [11]}),
    .fco(\u2_Display/add134/c15 ),
    .fx({\u2_Display/n4383 [14],\u2_Display/n4383 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u15_al_u4226  (
    .a({\u2_Display/n4363 ,\u2_Display/n4365 }),
    .b({\u2_Display/n4362 ,\u2_Display/n4364 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add134/c15 ),
    .f({\u2_Display/n4383 [17],\u2_Display/n4383 [15]}),
    .fco(\u2_Display/add134/c19 ),
    .fx({\u2_Display/n4383 [18],\u2_Display/n4383 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u19_al_u4227  (
    .a({\u2_Display/n4359 ,\u2_Display/n4361 }),
    .b({\u2_Display/n4358 ,\u2_Display/n4360 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add134/c19 ),
    .f({\u2_Display/n4383 [21],\u2_Display/n4383 [19]}),
    .fco(\u2_Display/add134/c23 ),
    .fx({\u2_Display/n4383 [22],\u2_Display/n4383 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u23_al_u4228  (
    .a({\u2_Display/n4355 ,\u2_Display/n4357 }),
    .b({\u2_Display/n4354 ,\u2_Display/n4356 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add134/c23 ),
    .f({\u2_Display/n4383 [25],\u2_Display/n4383 [23]}),
    .fco(\u2_Display/add134/c27 ),
    .fx({\u2_Display/n4383 [26],\u2_Display/n4383 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u27_al_u4229  (
    .a({\u2_Display/n4351 ,\u2_Display/n4353 }),
    .b({\u2_Display/n4350 ,\u2_Display/n4352 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add134/c27 ),
    .f({\u2_Display/n4383 [29],\u2_Display/n4383 [27]}),
    .fco(\u2_Display/add134/c31 ),
    .fx({\u2_Display/n4383 [30],\u2_Display/n4383 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u31_al_u4230  (
    .a({open_n7062,\u2_Display/n4349 }),
    .c(2'b00),
    .d({open_n7067,1'b1}),
    .fci(\u2_Display/add134/c31 ),
    .f({open_n7084,\u2_Display/n4383 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u3_al_u4223  (
    .a({\u2_Display/n4375 ,\u2_Display/n4377 }),
    .b({\u2_Display/n4374 ,\u2_Display/n4376 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add134/c3 ),
    .f({\u2_Display/n4383 [5],\u2_Display/n4383 [3]}),
    .fco(\u2_Display/add134/c7 ),
    .fx({\u2_Display/n4383 [6],\u2_Display/n4383 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/u7_al_u4224  (
    .a({\u2_Display/n4371 ,\u2_Display/n4373 }),
    .b({\u2_Display/n4370 ,\u2_Display/n4372 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add134/c7 ),
    .f({\u2_Display/n4383 [9],\u2_Display/n4383 [7]}),
    .fco(\u2_Display/add134/c11 ),
    .fx({\u2_Display/n4383 [10],\u2_Display/n4383 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add134/ucin_al_u4222"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add134/ucin_al_u4222  (
    .a({\u2_Display/n4379 ,1'b1}),
    .b({\u2_Display/n4378 ,\u2_Display/n4380 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4383 [1],open_n7143}),
    .fco(\u2_Display/add134/c3 ),
    .fx({\u2_Display/n4383 [2],\u2_Display/n4383 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u11_al_u4234  (
    .a({\u2_Display/n4402 ,\u2_Display/n4404 }),
    .b({\u2_Display/n4401 ,\u2_Display/n4403 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add135/c11 ),
    .f({\u2_Display/n4418 [13],\u2_Display/n4418 [11]}),
    .fco(\u2_Display/add135/c15 ),
    .fx({\u2_Display/n4418 [14],\u2_Display/n4418 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u15_al_u4235  (
    .a({\u2_Display/n4398 ,\u2_Display/n4400 }),
    .b({\u2_Display/n4397 ,\u2_Display/n4399 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add135/c15 ),
    .f({\u2_Display/n4418 [17],\u2_Display/n4418 [15]}),
    .fco(\u2_Display/add135/c19 ),
    .fx({\u2_Display/n4418 [18],\u2_Display/n4418 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u19_al_u4236  (
    .a({\u2_Display/n4394 ,\u2_Display/n4396 }),
    .b({\u2_Display/n4393 ,\u2_Display/n4395 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add135/c19 ),
    .f({\u2_Display/n4418 [21],\u2_Display/n4418 [19]}),
    .fco(\u2_Display/add135/c23 ),
    .fx({\u2_Display/n4418 [22],\u2_Display/n4418 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u23_al_u4237  (
    .a({\u2_Display/n4390 ,\u2_Display/n4392 }),
    .b({\u2_Display/n4389 ,\u2_Display/n4391 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add135/c23 ),
    .f({\u2_Display/n4418 [25],\u2_Display/n4418 [23]}),
    .fco(\u2_Display/add135/c27 ),
    .fx({\u2_Display/n4418 [26],\u2_Display/n4418 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u27_al_u4238  (
    .a({\u2_Display/n4386 ,\u2_Display/n4388 }),
    .b({\u2_Display/n4385 ,\u2_Display/n4387 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add135/c27 ),
    .f({\u2_Display/n4418 [29],\u2_Display/n4418 [27]}),
    .fco(\u2_Display/add135/c31 ),
    .fx({\u2_Display/n4418 [30],\u2_Display/n4418 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u31_al_u4239  (
    .a({open_n7236,\u2_Display/n4384 }),
    .c(2'b00),
    .d({open_n7241,1'b1}),
    .fci(\u2_Display/add135/c31 ),
    .f({open_n7258,\u2_Display/n4418 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u3_al_u4232  (
    .a({\u2_Display/n4410 ,\u2_Display/n4412 }),
    .b({\u2_Display/n4409 ,\u2_Display/n4411 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add135/c3 ),
    .f({\u2_Display/n4418 [5],\u2_Display/n4418 [3]}),
    .fco(\u2_Display/add135/c7 ),
    .fx({\u2_Display/n4418 [6],\u2_Display/n4418 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/u7_al_u4233  (
    .a({\u2_Display/n4406 ,\u2_Display/n4408 }),
    .b({\u2_Display/n4405 ,\u2_Display/n4407 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add135/c7 ),
    .f({\u2_Display/n4418 [9],\u2_Display/n4418 [7]}),
    .fco(\u2_Display/add135/c11 ),
    .fx({\u2_Display/n4418 [10],\u2_Display/n4418 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add135/ucin_al_u4231"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add135/ucin_al_u4231  (
    .a({\u2_Display/n4414 ,1'b1}),
    .b({\u2_Display/n4413 ,\u2_Display/n4415 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4418 [1],open_n7317}),
    .fco(\u2_Display/add135/c3 ),
    .fx({\u2_Display/n4418 [2],\u2_Display/n4418 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u11_al_u4243  (
    .a({\u2_Display/n4437 ,\u2_Display/n4439 }),
    .b({\u2_Display/n4436 ,\u2_Display/n4438 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add136/c11 ),
    .f({\u2_Display/n4453 [13],\u2_Display/n4453 [11]}),
    .fco(\u2_Display/add136/c15 ),
    .fx({\u2_Display/n4453 [14],\u2_Display/n4453 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u15_al_u4244  (
    .a({\u2_Display/n4433 ,\u2_Display/n4435 }),
    .b({\u2_Display/n4432 ,\u2_Display/n4434 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add136/c15 ),
    .f({\u2_Display/n4453 [17],\u2_Display/n4453 [15]}),
    .fco(\u2_Display/add136/c19 ),
    .fx({\u2_Display/n4453 [18],\u2_Display/n4453 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u19_al_u4245  (
    .a({\u2_Display/n4429 ,\u2_Display/n4431 }),
    .b({\u2_Display/n4428 ,\u2_Display/n4430 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add136/c19 ),
    .f({\u2_Display/n4453 [21],\u2_Display/n4453 [19]}),
    .fco(\u2_Display/add136/c23 ),
    .fx({\u2_Display/n4453 [22],\u2_Display/n4453 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u23_al_u4246  (
    .a({\u2_Display/n4425 ,\u2_Display/n4427 }),
    .b({\u2_Display/n4424 ,\u2_Display/n4426 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add136/c23 ),
    .f({\u2_Display/n4453 [25],\u2_Display/n4453 [23]}),
    .fco(\u2_Display/add136/c27 ),
    .fx({\u2_Display/n4453 [26],\u2_Display/n4453 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u27_al_u4247  (
    .a({\u2_Display/n4421 ,\u2_Display/n4423 }),
    .b({\u2_Display/n4420 ,\u2_Display/n4422 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add136/c27 ),
    .f({\u2_Display/n4453 [29],\u2_Display/n4453 [27]}),
    .fco(\u2_Display/add136/c31 ),
    .fx({\u2_Display/n4453 [30],\u2_Display/n4453 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u31_al_u4248  (
    .a({open_n7410,\u2_Display/n4419 }),
    .c(2'b00),
    .d({open_n7415,1'b1}),
    .fci(\u2_Display/add136/c31 ),
    .f({open_n7432,\u2_Display/n4453 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u3_al_u4241  (
    .a({\u2_Display/n4445 ,\u2_Display/n4447 }),
    .b({\u2_Display/n4444 ,\u2_Display/n4446 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add136/c3 ),
    .f({\u2_Display/n4453 [5],\u2_Display/n4453 [3]}),
    .fco(\u2_Display/add136/c7 ),
    .fx({\u2_Display/n4453 [6],\u2_Display/n4453 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/u7_al_u4242  (
    .a({\u2_Display/n4441 ,\u2_Display/n4443 }),
    .b({\u2_Display/n4440 ,\u2_Display/n4442 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add136/c7 ),
    .f({\u2_Display/n4453 [9],\u2_Display/n4453 [7]}),
    .fco(\u2_Display/add136/c11 ),
    .fx({\u2_Display/n4453 [10],\u2_Display/n4453 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add136/ucin_al_u4240"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add136/ucin_al_u4240  (
    .a({\u2_Display/n4449 ,1'b1}),
    .b({\u2_Display/n4448 ,\u2_Display/n4450 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4453 [1],open_n7491}),
    .fco(\u2_Display/add136/c3 ),
    .fx({\u2_Display/n4453 [2],\u2_Display/n4453 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u11_al_u4252  (
    .a({\u2_Display/n4472 ,\u2_Display/n4474 }),
    .b({\u2_Display/n4471 ,\u2_Display/n4473 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add137/c11 ),
    .f({\u2_Display/n4488 [13],\u2_Display/n4488 [11]}),
    .fco(\u2_Display/add137/c15 ),
    .fx({\u2_Display/n4488 [14],\u2_Display/n4488 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u15_al_u4253  (
    .a({\u2_Display/n4468 ,\u2_Display/n4470 }),
    .b({\u2_Display/n4467 ,\u2_Display/n4469 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add137/c15 ),
    .f({\u2_Display/n4488 [17],\u2_Display/n4488 [15]}),
    .fco(\u2_Display/add137/c19 ),
    .fx({\u2_Display/n4488 [18],\u2_Display/n4488 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u19_al_u4254  (
    .a({\u2_Display/n4464 ,\u2_Display/n4466 }),
    .b({\u2_Display/n4463 ,\u2_Display/n4465 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add137/c19 ),
    .f({\u2_Display/n4488 [21],\u2_Display/n4488 [19]}),
    .fco(\u2_Display/add137/c23 ),
    .fx({\u2_Display/n4488 [22],\u2_Display/n4488 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u23_al_u4255  (
    .a({\u2_Display/n4460 ,\u2_Display/n4462 }),
    .b({\u2_Display/n4459 ,\u2_Display/n4461 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add137/c23 ),
    .f({\u2_Display/n4488 [25],\u2_Display/n4488 [23]}),
    .fco(\u2_Display/add137/c27 ),
    .fx({\u2_Display/n4488 [26],\u2_Display/n4488 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u27_al_u4256  (
    .a({\u2_Display/n4456 ,\u2_Display/n4458 }),
    .b({\u2_Display/n4455 ,\u2_Display/n4457 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add137/c27 ),
    .f({\u2_Display/n4488 [29],\u2_Display/n4488 [27]}),
    .fco(\u2_Display/add137/c31 ),
    .fx({\u2_Display/n4488 [30],\u2_Display/n4488 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u31_al_u4257  (
    .a({open_n7584,\u2_Display/n4454 }),
    .c(2'b00),
    .d({open_n7589,1'b1}),
    .fci(\u2_Display/add137/c31 ),
    .f({open_n7606,\u2_Display/n4488 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u3_al_u4250  (
    .a({\u2_Display/n4480 ,\u2_Display/n4482 }),
    .b({\u2_Display/n4479 ,\u2_Display/n4481 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add137/c3 ),
    .f({\u2_Display/n4488 [5],\u2_Display/n4488 [3]}),
    .fco(\u2_Display/add137/c7 ),
    .fx({\u2_Display/n4488 [6],\u2_Display/n4488 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/u7_al_u4251  (
    .a({\u2_Display/n4476 ,\u2_Display/n4478 }),
    .b({\u2_Display/n4475 ,\u2_Display/n4477 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add137/c7 ),
    .f({\u2_Display/n4488 [9],\u2_Display/n4488 [7]}),
    .fco(\u2_Display/add137/c11 ),
    .fx({\u2_Display/n4488 [10],\u2_Display/n4488 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add137/ucin_al_u4249"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add137/ucin_al_u4249  (
    .a({\u2_Display/n4484 ,1'b1}),
    .b({\u2_Display/n4483 ,\u2_Display/n4485 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4488 [1],open_n7665}),
    .fco(\u2_Display/add137/c3 ),
    .fx({\u2_Display/n4488 [2],\u2_Display/n4488 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u11_al_u4261  (
    .a({\u2_Display/n4507 ,\u2_Display/n4509 }),
    .b({\u2_Display/n4506 ,\u2_Display/n4508 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add138/c11 ),
    .f({\u2_Display/n4523 [13],\u2_Display/n4523 [11]}),
    .fco(\u2_Display/add138/c15 ),
    .fx({\u2_Display/n4523 [14],\u2_Display/n4523 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u15_al_u4262  (
    .a({\u2_Display/n4503 ,\u2_Display/n4505 }),
    .b({\u2_Display/n4502 ,\u2_Display/n4504 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add138/c15 ),
    .f({\u2_Display/n4523 [17],\u2_Display/n4523 [15]}),
    .fco(\u2_Display/add138/c19 ),
    .fx({\u2_Display/n4523 [18],\u2_Display/n4523 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u19_al_u4263  (
    .a({\u2_Display/n4499 ,\u2_Display/n4501 }),
    .b({\u2_Display/n4498 ,\u2_Display/n4500 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add138/c19 ),
    .f({\u2_Display/n4523 [21],\u2_Display/n4523 [19]}),
    .fco(\u2_Display/add138/c23 ),
    .fx({\u2_Display/n4523 [22],\u2_Display/n4523 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u23_al_u4264  (
    .a({\u2_Display/n4495 ,\u2_Display/n4497 }),
    .b({\u2_Display/n4494 ,\u2_Display/n4496 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add138/c23 ),
    .f({\u2_Display/n4523 [25],\u2_Display/n4523 [23]}),
    .fco(\u2_Display/add138/c27 ),
    .fx({\u2_Display/n4523 [26],\u2_Display/n4523 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u27_al_u4265  (
    .a({\u2_Display/n4491 ,\u2_Display/n4493 }),
    .b({\u2_Display/n4490 ,\u2_Display/n4492 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add138/c27 ),
    .f({\u2_Display/n4523 [29],\u2_Display/n4523 [27]}),
    .fco(\u2_Display/add138/c31 ),
    .fx({\u2_Display/n4523 [30],\u2_Display/n4523 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u31_al_u4266  (
    .a({open_n7758,\u2_Display/n4489 }),
    .c(2'b00),
    .d({open_n7763,1'b1}),
    .fci(\u2_Display/add138/c31 ),
    .f({open_n7780,\u2_Display/n4523 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u3_al_u4259  (
    .a({\u2_Display/n4515 ,\u2_Display/n4517 }),
    .b({\u2_Display/n4514 ,\u2_Display/n4516 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add138/c3 ),
    .f({\u2_Display/n4523 [5],\u2_Display/n4523 [3]}),
    .fco(\u2_Display/add138/c7 ),
    .fx({\u2_Display/n4523 [6],\u2_Display/n4523 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/u7_al_u4260  (
    .a({\u2_Display/n4511 ,\u2_Display/n4513 }),
    .b({\u2_Display/n4510 ,\u2_Display/n4512 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add138/c7 ),
    .f({\u2_Display/n4523 [9],\u2_Display/n4523 [7]}),
    .fco(\u2_Display/add138/c11 ),
    .fx({\u2_Display/n4523 [10],\u2_Display/n4523 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add138/ucin_al_u4258"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add138/ucin_al_u4258  (
    .a({\u2_Display/n4519 ,1'b1}),
    .b({\u2_Display/n4518 ,\u2_Display/n4520 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4523 [1],open_n7839}),
    .fco(\u2_Display/add138/c3 ),
    .fx({\u2_Display/n4523 [2],\u2_Display/n4523 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add139/ucin_al_u5046"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add139/u3_al_u5047  (
    .a({\u2_Display/n4550 ,\u2_Display/n4552 }),
    .b({\u2_Display/n4549 ,\u2_Display/n4551 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add139/c3 ),
    .f({\u2_Display/n4558 [5],\u2_Display/n4558 [3]}),
    .fco(\u2_Display/add139/c7 ),
    .fx({\u2_Display/n4558 [6],\u2_Display/n4558 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add139/ucin_al_u5046"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add139/u7_al_u5048  (
    .a({\u2_Display/n4546 ,\u2_Display/n4548 }),
    .b({open_n7860,\u2_Display/n4547 }),
    .c(2'b00),
    .d(2'b01),
    .e({open_n7863,1'b0}),
    .fci(\u2_Display/add139/c7 ),
    .f({\u2_Display/n4558 [9],\u2_Display/n4558 [7]}),
    .fx({open_n7879,\u2_Display/n4558 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add139/ucin_al_u5046"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add139/ucin_al_u5046  (
    .a({\u2_Display/n4554 ,1'b1}),
    .b({\u2_Display/n4553 ,\u2_Display/n4555 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4558 [1],open_n7899}),
    .fco(\u2_Display/add139/c3 ),
    .fx({\u2_Display/n4558 [2],\u2_Display/n4558 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u11_al_u4270  (
    .a({\u2_Display/counta [13],\u2_Display/counta [11]}),
    .b({\u2_Display/counta [14],\u2_Display/counta [12]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add14/c11 ),
    .f({\u2_Display/n4911 [13],\u2_Display/n4911 [11]}),
    .fco(\u2_Display/add14/c15 ),
    .fx({\u2_Display/n4911 [14],\u2_Display/n4911 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u15_al_u4271  (
    .a({\u2_Display/counta [17],\u2_Display/counta [15]}),
    .b({\u2_Display/counta [18],\u2_Display/counta [16]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add14/c15 ),
    .f({\u2_Display/n4911 [17],\u2_Display/n4911 [15]}),
    .fco(\u2_Display/add14/c19 ),
    .fx({\u2_Display/n4911 [18],\u2_Display/n4911 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u19_al_u4272  (
    .a({\u2_Display/counta [21],\u2_Display/counta [19]}),
    .b({\u2_Display/counta [22],\u2_Display/counta [20]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add14/c19 ),
    .f({\u2_Display/n4911 [21],\u2_Display/n4911 [19]}),
    .fco(\u2_Display/add14/c23 ),
    .fx({\u2_Display/n4911 [22],\u2_Display/n4911 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u23_al_u4273  (
    .a({\u2_Display/counta [25],\u2_Display/counta [23]}),
    .b({\u2_Display/counta [26],\u2_Display/counta [24]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add14/c23 ),
    .f({\u2_Display/n4911 [25],\u2_Display/n4911 [23]}),
    .fco(\u2_Display/add14/c27 ),
    .fx({\u2_Display/n4911 [26],\u2_Display/n4911 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u27_al_u4274  (
    .a({\u2_Display/counta [29],\u2_Display/counta [27]}),
    .b({\u2_Display/counta [30],\u2_Display/counta [28]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add14/c27 ),
    .f({\u2_Display/n4911 [29],\u2_Display/n4911 [27]}),
    .fco(\u2_Display/add14/c31 ),
    .fx({\u2_Display/n4911 [30],\u2_Display/n4911 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u31_al_u4275  (
    .a({open_n7992,\u2_Display/counta [31]}),
    .c(2'b00),
    .d({open_n7997,1'b0}),
    .fci(\u2_Display/add14/c31 ),
    .f({open_n8014,\u2_Display/n4911 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u3_al_u4268  (
    .a({\u2_Display/counta [5],\u2_Display/counta [3]}),
    .b({\u2_Display/counta [6],\u2_Display/counta [4]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add14/c3 ),
    .f({\u2_Display/n4911 [5],\u2_Display/n4911 [3]}),
    .fco(\u2_Display/add14/c7 ),
    .fx({\u2_Display/n4911 [6],\u2_Display/n4911 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/u7_al_u4269  (
    .a({\u2_Display/counta [9],\u2_Display/counta [7]}),
    .b({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add14/c7 ),
    .f({\u2_Display/n4911 [9],\u2_Display/n4911 [7]}),
    .fco(\u2_Display/add14/c11 ),
    .fx({\u2_Display/n4911 [10],\u2_Display/n4911 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add14/ucin_al_u4267"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add14/ucin_al_u4267  (
    .a({\u2_Display/counta [1],1'b1}),
    .b({\u2_Display/counta [2],\u2_Display/counta [0]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4911 [1],open_n8073}),
    .fco(\u2_Display/add14/c3 ),
    .fx({\u2_Display/n4911 [2],\u2_Display/n4911 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u11_al_u4279  (
    .a({\u2_Display/n6088 ,\u2_Display/n6090 }),
    .b({\u2_Display/n6087 ,\u2_Display/n6089 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add151/c11 ),
    .f({\u2_Display/n4946 [13],\u2_Display/n4946 [11]}),
    .fco(\u2_Display/add151/c15 ),
    .fx({\u2_Display/n4946 [14],\u2_Display/n4946 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u15_al_u4280  (
    .a({\u2_Display/n6084 ,\u2_Display/n6086 }),
    .b({\u2_Display/n6083 ,\u2_Display/n6085 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add151/c15 ),
    .f({\u2_Display/n4946 [17],\u2_Display/n4946 [15]}),
    .fco(\u2_Display/add151/c19 ),
    .fx({\u2_Display/n4946 [18],\u2_Display/n4946 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u19_al_u4281  (
    .a({\u2_Display/n6080 ,\u2_Display/n6082 }),
    .b({\u2_Display/n6079 ,\u2_Display/n6081 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add151/c19 ),
    .f({\u2_Display/n4946 [21],\u2_Display/n4946 [19]}),
    .fco(\u2_Display/add151/c23 ),
    .fx({\u2_Display/n4946 [22],\u2_Display/n4946 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u23_al_u4282  (
    .a({\u2_Display/n6076 ,\u2_Display/n6078 }),
    .b({\u2_Display/n6075 ,\u2_Display/n6077 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add151/c23 ),
    .f({\u2_Display/n4946 [25],\u2_Display/n4946 [23]}),
    .fco(\u2_Display/add151/c27 ),
    .fx({\u2_Display/n4946 [26],\u2_Display/n4946 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u27_al_u4283  (
    .a({\u2_Display/n6072 ,\u2_Display/n6074 }),
    .b({\u2_Display/n6071 ,\u2_Display/n6073 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add151/c27 ),
    .f({\u2_Display/n4946 [29],\u2_Display/n4946 [27]}),
    .fco(\u2_Display/add151/c31 ),
    .fx({\u2_Display/n4946 [30],\u2_Display/n4946 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u31_al_u4284  (
    .a({open_n8166,\u2_Display/n6070 }),
    .c(2'b00),
    .d({open_n8171,1'b1}),
    .fci(\u2_Display/add151/c31 ),
    .f({open_n8188,\u2_Display/n4946 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u3_al_u4277  (
    .a({\u2_Display/n6096 ,\u2_Display/n6098 }),
    .b({\u2_Display/n6095 ,\u2_Display/n6097 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add151/c3 ),
    .f({\u2_Display/n4946 [5],\u2_Display/n4946 [3]}),
    .fco(\u2_Display/add151/c7 ),
    .fx({\u2_Display/n4946 [6],\u2_Display/n4946 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/u7_al_u4278  (
    .a({\u2_Display/n6092 ,\u2_Display/n6094 }),
    .b({\u2_Display/n6091 ,\u2_Display/n6093 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add151/c7 ),
    .f({\u2_Display/n4946 [9],\u2_Display/n4946 [7]}),
    .fco(\u2_Display/add151/c11 ),
    .fx({\u2_Display/n4946 [10],\u2_Display/n4946 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add151/ucin_al_u4276"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add151/ucin_al_u4276  (
    .a({\u2_Display/n6100 ,1'b1}),
    .b({\u2_Display/n6099 ,\u2_Display/n6101 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4946 [1],open_n8247}),
    .fco(\u2_Display/add151/c3 ),
    .fx({\u2_Display/n4946 [2],\u2_Display/n4946 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u11_al_u4288  (
    .a({\u2_Display/n6123 ,\u2_Display/n6125 }),
    .b({\u2_Display/n6122 ,\u2_Display/n6124 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add152/c11 ),
    .f({\u2_Display/n4981 [13],\u2_Display/n4981 [11]}),
    .fco(\u2_Display/add152/c15 ),
    .fx({\u2_Display/n4981 [14],\u2_Display/n4981 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u15_al_u4289  (
    .a({\u2_Display/n6119 ,\u2_Display/n6121 }),
    .b({\u2_Display/n6118 ,\u2_Display/n6120 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add152/c15 ),
    .f({\u2_Display/n4981 [17],\u2_Display/n4981 [15]}),
    .fco(\u2_Display/add152/c19 ),
    .fx({\u2_Display/n4981 [18],\u2_Display/n4981 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u19_al_u4290  (
    .a({\u2_Display/n6115 ,\u2_Display/n6117 }),
    .b({\u2_Display/n6114 ,\u2_Display/n6116 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add152/c19 ),
    .f({\u2_Display/n4981 [21],\u2_Display/n4981 [19]}),
    .fco(\u2_Display/add152/c23 ),
    .fx({\u2_Display/n4981 [22],\u2_Display/n4981 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u23_al_u4291  (
    .a({\u2_Display/n6111 ,\u2_Display/n6113 }),
    .b({\u2_Display/n6110 ,\u2_Display/n6112 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add152/c23 ),
    .f({\u2_Display/n4981 [25],\u2_Display/n4981 [23]}),
    .fco(\u2_Display/add152/c27 ),
    .fx({\u2_Display/n4981 [26],\u2_Display/n4981 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u27_al_u4292  (
    .a({\u2_Display/n6107 ,\u2_Display/n6109 }),
    .b({\u2_Display/n6106 ,\u2_Display/n6108 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add152/c27 ),
    .f({\u2_Display/n4981 [29],\u2_Display/n4981 [27]}),
    .fco(\u2_Display/add152/c31 ),
    .fx({\u2_Display/n4981 [30],\u2_Display/n4981 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u31_al_u4293  (
    .a({open_n8340,\u2_Display/n6105 }),
    .c(2'b00),
    .d({open_n8345,1'b1}),
    .fci(\u2_Display/add152/c31 ),
    .f({open_n8362,\u2_Display/n4981 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u3_al_u4286  (
    .a({\u2_Display/n6131 ,\u2_Display/n6133 }),
    .b({\u2_Display/n6130 ,\u2_Display/n6132 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add152/c3 ),
    .f({\u2_Display/n4981 [5],\u2_Display/n4981 [3]}),
    .fco(\u2_Display/add152/c7 ),
    .fx({\u2_Display/n4981 [6],\u2_Display/n4981 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/u7_al_u4287  (
    .a({\u2_Display/n6127 ,\u2_Display/n6129 }),
    .b({\u2_Display/n6126 ,\u2_Display/n6128 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add152/c7 ),
    .f({\u2_Display/n4981 [9],\u2_Display/n4981 [7]}),
    .fco(\u2_Display/add152/c11 ),
    .fx({\u2_Display/n4981 [10],\u2_Display/n4981 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add152/ucin_al_u4285"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add152/ucin_al_u4285  (
    .a({\u2_Display/n6135 ,1'b1}),
    .b({\u2_Display/n6134 ,\u2_Display/n6136 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n4981 [1],open_n8421}),
    .fco(\u2_Display/add152/c3 ),
    .fx({\u2_Display/n4981 [2],\u2_Display/n4981 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u11_al_u4297  (
    .a({\u2_Display/n6158 ,\u2_Display/n6160 }),
    .b({\u2_Display/n6157 ,\u2_Display/n6159 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add153/c11 ),
    .f({\u2_Display/n5016 [13],\u2_Display/n5016 [11]}),
    .fco(\u2_Display/add153/c15 ),
    .fx({\u2_Display/n5016 [14],\u2_Display/n5016 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u15_al_u4298  (
    .a({\u2_Display/n6154 ,\u2_Display/n6156 }),
    .b({\u2_Display/n6153 ,\u2_Display/n6155 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add153/c15 ),
    .f({\u2_Display/n5016 [17],\u2_Display/n5016 [15]}),
    .fco(\u2_Display/add153/c19 ),
    .fx({\u2_Display/n5016 [18],\u2_Display/n5016 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u19_al_u4299  (
    .a({\u2_Display/n6150 ,\u2_Display/n6152 }),
    .b({\u2_Display/n6149 ,\u2_Display/n6151 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add153/c19 ),
    .f({\u2_Display/n5016 [21],\u2_Display/n5016 [19]}),
    .fco(\u2_Display/add153/c23 ),
    .fx({\u2_Display/n5016 [22],\u2_Display/n5016 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u23_al_u4300  (
    .a({\u2_Display/n6146 ,\u2_Display/n6148 }),
    .b({\u2_Display/n6145 ,\u2_Display/n6147 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add153/c23 ),
    .f({\u2_Display/n5016 [25],\u2_Display/n5016 [23]}),
    .fco(\u2_Display/add153/c27 ),
    .fx({\u2_Display/n5016 [26],\u2_Display/n5016 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u27_al_u4301  (
    .a({\u2_Display/n6142 ,\u2_Display/n6144 }),
    .b({\u2_Display/n6141 ,\u2_Display/n6143 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add153/c27 ),
    .f({\u2_Display/n5016 [29],\u2_Display/n5016 [27]}),
    .fco(\u2_Display/add153/c31 ),
    .fx({\u2_Display/n5016 [30],\u2_Display/n5016 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u31_al_u4302  (
    .a({open_n8514,\u2_Display/n6140 }),
    .c(2'b00),
    .d({open_n8519,1'b1}),
    .fci(\u2_Display/add153/c31 ),
    .f({open_n8536,\u2_Display/n5016 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u3_al_u4295  (
    .a({\u2_Display/n6166 ,\u2_Display/n6168 }),
    .b({\u2_Display/n6165 ,\u2_Display/n6167 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add153/c3 ),
    .f({\u2_Display/n5016 [5],\u2_Display/n5016 [3]}),
    .fco(\u2_Display/add153/c7 ),
    .fx({\u2_Display/n5016 [6],\u2_Display/n5016 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/u7_al_u4296  (
    .a({\u2_Display/n6162 ,\u2_Display/n6164 }),
    .b({\u2_Display/n6161 ,\u2_Display/n6163 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add153/c7 ),
    .f({\u2_Display/n5016 [9],\u2_Display/n5016 [7]}),
    .fco(\u2_Display/add153/c11 ),
    .fx({\u2_Display/n5016 [10],\u2_Display/n5016 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add153/ucin_al_u4294"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add153/ucin_al_u4294  (
    .a({\u2_Display/n6170 ,1'b1}),
    .b({\u2_Display/n6169 ,\u2_Display/n6171 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5016 [1],open_n8595}),
    .fco(\u2_Display/add153/c3 ),
    .fx({\u2_Display/n5016 [2],\u2_Display/n5016 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u11_al_u4306  (
    .a({\u2_Display/n6193 ,\u2_Display/n6195 }),
    .b({\u2_Display/n6192 ,\u2_Display/n6194 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add154/c11 ),
    .f({\u2_Display/n5051 [13],\u2_Display/n5051 [11]}),
    .fco(\u2_Display/add154/c15 ),
    .fx({\u2_Display/n5051 [14],\u2_Display/n5051 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u15_al_u4307  (
    .a({\u2_Display/n6189 ,\u2_Display/n6191 }),
    .b({\u2_Display/n6188 ,\u2_Display/n6190 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add154/c15 ),
    .f({\u2_Display/n5051 [17],\u2_Display/n5051 [15]}),
    .fco(\u2_Display/add154/c19 ),
    .fx({\u2_Display/n5051 [18],\u2_Display/n5051 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u19_al_u4308  (
    .a({\u2_Display/n6185 ,\u2_Display/n6187 }),
    .b({\u2_Display/n6184 ,\u2_Display/n6186 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add154/c19 ),
    .f({\u2_Display/n5051 [21],\u2_Display/n5051 [19]}),
    .fco(\u2_Display/add154/c23 ),
    .fx({\u2_Display/n5051 [22],\u2_Display/n5051 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u23_al_u4309  (
    .a({\u2_Display/n6181 ,\u2_Display/n6183 }),
    .b({\u2_Display/n6180 ,\u2_Display/n6182 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add154/c23 ),
    .f({\u2_Display/n5051 [25],\u2_Display/n5051 [23]}),
    .fco(\u2_Display/add154/c27 ),
    .fx({\u2_Display/n5051 [26],\u2_Display/n5051 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u27_al_u4310  (
    .a({\u2_Display/n6177 ,\u2_Display/n6179 }),
    .b({\u2_Display/n6176 ,\u2_Display/n6178 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add154/c27 ),
    .f({\u2_Display/n5051 [29],\u2_Display/n5051 [27]}),
    .fco(\u2_Display/add154/c31 ),
    .fx({\u2_Display/n5051 [30],\u2_Display/n5051 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u31_al_u4311  (
    .a({open_n8688,\u2_Display/n6175 }),
    .c(2'b00),
    .d({open_n8693,1'b1}),
    .fci(\u2_Display/add154/c31 ),
    .f({open_n8710,\u2_Display/n5051 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u3_al_u4304  (
    .a({\u2_Display/n6201 ,\u2_Display/n6203 }),
    .b({\u2_Display/n6200 ,\u2_Display/n6202 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add154/c3 ),
    .f({\u2_Display/n5051 [5],\u2_Display/n5051 [3]}),
    .fco(\u2_Display/add154/c7 ),
    .fx({\u2_Display/n5051 [6],\u2_Display/n5051 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/u7_al_u4305  (
    .a({\u2_Display/n6197 ,\u2_Display/n6199 }),
    .b({\u2_Display/n6196 ,\u2_Display/n6198 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add154/c7 ),
    .f({\u2_Display/n5051 [9],\u2_Display/n5051 [7]}),
    .fco(\u2_Display/add154/c11 ),
    .fx({\u2_Display/n5051 [10],\u2_Display/n5051 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add154/ucin_al_u4303"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add154/ucin_al_u4303  (
    .a({\u2_Display/n6205 ,1'b1}),
    .b({\u2_Display/n6204 ,\u2_Display/n6206 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5051 [1],open_n8769}),
    .fco(\u2_Display/add154/c3 ),
    .fx({\u2_Display/n5051 [2],\u2_Display/n5051 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u11_al_u4315  (
    .a({\u2_Display/n6228 ,\u2_Display/n6230 }),
    .b({\u2_Display/n6227 ,\u2_Display/n6229 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add155/c11 ),
    .f({\u2_Display/n5086 [13],\u2_Display/n5086 [11]}),
    .fco(\u2_Display/add155/c15 ),
    .fx({\u2_Display/n5086 [14],\u2_Display/n5086 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u15_al_u4316  (
    .a({\u2_Display/n6224 ,\u2_Display/n6226 }),
    .b({\u2_Display/n6223 ,\u2_Display/n6225 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add155/c15 ),
    .f({\u2_Display/n5086 [17],\u2_Display/n5086 [15]}),
    .fco(\u2_Display/add155/c19 ),
    .fx({\u2_Display/n5086 [18],\u2_Display/n5086 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u19_al_u4317  (
    .a({\u2_Display/n6220 ,\u2_Display/n6222 }),
    .b({\u2_Display/n6219 ,\u2_Display/n6221 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add155/c19 ),
    .f({\u2_Display/n5086 [21],\u2_Display/n5086 [19]}),
    .fco(\u2_Display/add155/c23 ),
    .fx({\u2_Display/n5086 [22],\u2_Display/n5086 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u23_al_u4318  (
    .a({\u2_Display/n6216 ,\u2_Display/n6218 }),
    .b({\u2_Display/n6215 ,\u2_Display/n6217 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add155/c23 ),
    .f({\u2_Display/n5086 [25],\u2_Display/n5086 [23]}),
    .fco(\u2_Display/add155/c27 ),
    .fx({\u2_Display/n5086 [26],\u2_Display/n5086 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u27_al_u4319  (
    .a({\u2_Display/n6212 ,\u2_Display/n6214 }),
    .b({\u2_Display/n6211 ,\u2_Display/n6213 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add155/c27 ),
    .f({\u2_Display/n5086 [29],\u2_Display/n5086 [27]}),
    .fco(\u2_Display/add155/c31 ),
    .fx({\u2_Display/n5086 [30],\u2_Display/n5086 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u31_al_u4320  (
    .a({open_n8862,\u2_Display/n6210 }),
    .c(2'b00),
    .d({open_n8867,1'b1}),
    .fci(\u2_Display/add155/c31 ),
    .f({open_n8884,\u2_Display/n5086 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u3_al_u4313  (
    .a({\u2_Display/n6236 ,\u2_Display/n6238 }),
    .b({\u2_Display/n6235 ,\u2_Display/n6237 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add155/c3 ),
    .f({\u2_Display/n5086 [5],\u2_Display/n5086 [3]}),
    .fco(\u2_Display/add155/c7 ),
    .fx({\u2_Display/n5086 [6],\u2_Display/n5086 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/u7_al_u4314  (
    .a({\u2_Display/n6232 ,\u2_Display/n6234 }),
    .b({\u2_Display/n6231 ,\u2_Display/n6233 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add155/c7 ),
    .f({\u2_Display/n5086 [9],\u2_Display/n5086 [7]}),
    .fco(\u2_Display/add155/c11 ),
    .fx({\u2_Display/n5086 [10],\u2_Display/n5086 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add155/ucin_al_u4312"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add155/ucin_al_u4312  (
    .a({\u2_Display/n6240 ,1'b1}),
    .b({\u2_Display/n6239 ,\u2_Display/n6241 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5086 [1],open_n8943}),
    .fco(\u2_Display/add155/c3 ),
    .fx({\u2_Display/n5086 [2],\u2_Display/n5086 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u11_al_u4324  (
    .a({\u2_Display/n6263 ,\u2_Display/n6265 }),
    .b({\u2_Display/n6262 ,\u2_Display/n6264 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add156/c11 ),
    .f({\u2_Display/n5121 [13],\u2_Display/n5121 [11]}),
    .fco(\u2_Display/add156/c15 ),
    .fx({\u2_Display/n5121 [14],\u2_Display/n5121 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u15_al_u4325  (
    .a({\u2_Display/n6259 ,\u2_Display/n6261 }),
    .b({\u2_Display/n6258 ,\u2_Display/n6260 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add156/c15 ),
    .f({\u2_Display/n5121 [17],\u2_Display/n5121 [15]}),
    .fco(\u2_Display/add156/c19 ),
    .fx({\u2_Display/n5121 [18],\u2_Display/n5121 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u19_al_u4326  (
    .a({\u2_Display/n6255 ,\u2_Display/n6257 }),
    .b({\u2_Display/n6254 ,\u2_Display/n6256 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add156/c19 ),
    .f({\u2_Display/n5121 [21],\u2_Display/n5121 [19]}),
    .fco(\u2_Display/add156/c23 ),
    .fx({\u2_Display/n5121 [22],\u2_Display/n5121 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u23_al_u4327  (
    .a({\u2_Display/n6251 ,\u2_Display/n6253 }),
    .b({\u2_Display/n6250 ,\u2_Display/n6252 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add156/c23 ),
    .f({\u2_Display/n5121 [25],\u2_Display/n5121 [23]}),
    .fco(\u2_Display/add156/c27 ),
    .fx({\u2_Display/n5121 [26],\u2_Display/n5121 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u27_al_u4328  (
    .a({\u2_Display/n6247 ,\u2_Display/n6249 }),
    .b({\u2_Display/n6246 ,\u2_Display/n6248 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add156/c27 ),
    .f({\u2_Display/n5121 [29],\u2_Display/n5121 [27]}),
    .fco(\u2_Display/add156/c31 ),
    .fx({\u2_Display/n5121 [30],\u2_Display/n5121 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u31_al_u4329  (
    .a({open_n9036,\u2_Display/n6245 }),
    .c(2'b00),
    .d({open_n9041,1'b1}),
    .fci(\u2_Display/add156/c31 ),
    .f({open_n9058,\u2_Display/n5121 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u3_al_u4322  (
    .a({\u2_Display/n6271 ,\u2_Display/n6273 }),
    .b({\u2_Display/n6270 ,\u2_Display/n6272 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add156/c3 ),
    .f({\u2_Display/n5121 [5],\u2_Display/n5121 [3]}),
    .fco(\u2_Display/add156/c7 ),
    .fx({\u2_Display/n5121 [6],\u2_Display/n5121 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/u7_al_u4323  (
    .a({\u2_Display/n6267 ,\u2_Display/n6269 }),
    .b({\u2_Display/n6266 ,\u2_Display/n6268 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add156/c7 ),
    .f({\u2_Display/n5121 [9],\u2_Display/n5121 [7]}),
    .fco(\u2_Display/add156/c11 ),
    .fx({\u2_Display/n5121 [10],\u2_Display/n5121 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add156/ucin_al_u4321"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add156/ucin_al_u4321  (
    .a({\u2_Display/n6275 ,1'b1}),
    .b({\u2_Display/n6274 ,\u2_Display/n6276 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5121 [1],open_n9117}),
    .fco(\u2_Display/add156/c3 ),
    .fx({\u2_Display/n5121 [2],\u2_Display/n5121 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u11_al_u4333  (
    .a({\u2_Display/n6298 ,\u2_Display/n6300 }),
    .b({\u2_Display/n6297 ,\u2_Display/n6299 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add157/c11 ),
    .f({\u2_Display/n5156 [13],\u2_Display/n5156 [11]}),
    .fco(\u2_Display/add157/c15 ),
    .fx({\u2_Display/n5156 [14],\u2_Display/n5156 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u15_al_u4334  (
    .a({\u2_Display/n6294 ,\u2_Display/n6296 }),
    .b({\u2_Display/n6293 ,\u2_Display/n6295 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add157/c15 ),
    .f({\u2_Display/n5156 [17],\u2_Display/n5156 [15]}),
    .fco(\u2_Display/add157/c19 ),
    .fx({\u2_Display/n5156 [18],\u2_Display/n5156 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u19_al_u4335  (
    .a({\u2_Display/n6290 ,\u2_Display/n6292 }),
    .b({\u2_Display/n6289 ,\u2_Display/n6291 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add157/c19 ),
    .f({\u2_Display/n5156 [21],\u2_Display/n5156 [19]}),
    .fco(\u2_Display/add157/c23 ),
    .fx({\u2_Display/n5156 [22],\u2_Display/n5156 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u23_al_u4336  (
    .a({\u2_Display/n6286 ,\u2_Display/n6288 }),
    .b({\u2_Display/n6285 ,\u2_Display/n6287 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add157/c23 ),
    .f({\u2_Display/n5156 [25],\u2_Display/n5156 [23]}),
    .fco(\u2_Display/add157/c27 ),
    .fx({\u2_Display/n5156 [26],\u2_Display/n5156 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u27_al_u4337  (
    .a({\u2_Display/n6282 ,\u2_Display/n6284 }),
    .b({\u2_Display/n6281 ,\u2_Display/n6283 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add157/c27 ),
    .f({\u2_Display/n5156 [29],\u2_Display/n5156 [27]}),
    .fco(\u2_Display/add157/c31 ),
    .fx({\u2_Display/n5156 [30],\u2_Display/n5156 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u31_al_u4338  (
    .a({open_n9210,\u2_Display/n6280 }),
    .c(2'b00),
    .d({open_n9215,1'b1}),
    .fci(\u2_Display/add157/c31 ),
    .f({open_n9232,\u2_Display/n5156 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u3_al_u4331  (
    .a({\u2_Display/n6306 ,\u2_Display/n6308 }),
    .b({\u2_Display/n6305 ,\u2_Display/n6307 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add157/c3 ),
    .f({\u2_Display/n5156 [5],\u2_Display/n5156 [3]}),
    .fco(\u2_Display/add157/c7 ),
    .fx({\u2_Display/n5156 [6],\u2_Display/n5156 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/u7_al_u4332  (
    .a({\u2_Display/n6302 ,\u2_Display/n6304 }),
    .b({\u2_Display/n6301 ,\u2_Display/n6303 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add157/c7 ),
    .f({\u2_Display/n5156 [9],\u2_Display/n5156 [7]}),
    .fco(\u2_Display/add157/c11 ),
    .fx({\u2_Display/n5156 [10],\u2_Display/n5156 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add157/ucin_al_u4330"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add157/ucin_al_u4330  (
    .a({\u2_Display/n6310 ,1'b1}),
    .b({\u2_Display/n6309 ,\u2_Display/n6311 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5156 [1],open_n9291}),
    .fco(\u2_Display/add157/c3 ),
    .fx({\u2_Display/n5156 [2],\u2_Display/n5156 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u11_al_u4342  (
    .a({\u2_Display/n6333 ,\u2_Display/n6335 }),
    .b({\u2_Display/n6332 ,\u2_Display/n6334 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add158/c11 ),
    .f({\u2_Display/n5191 [13],\u2_Display/n5191 [11]}),
    .fco(\u2_Display/add158/c15 ),
    .fx({\u2_Display/n5191 [14],\u2_Display/n5191 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u15_al_u4343  (
    .a({\u2_Display/n6329 ,\u2_Display/n6331 }),
    .b({\u2_Display/n6328 ,\u2_Display/n6330 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add158/c15 ),
    .f({\u2_Display/n5191 [17],\u2_Display/n5191 [15]}),
    .fco(\u2_Display/add158/c19 ),
    .fx({\u2_Display/n5191 [18],\u2_Display/n5191 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u19_al_u4344  (
    .a({\u2_Display/n6325 ,\u2_Display/n6327 }),
    .b({\u2_Display/n6324 ,\u2_Display/n6326 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add158/c19 ),
    .f({\u2_Display/n5191 [21],\u2_Display/n5191 [19]}),
    .fco(\u2_Display/add158/c23 ),
    .fx({\u2_Display/n5191 [22],\u2_Display/n5191 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u23_al_u4345  (
    .a({\u2_Display/n6321 ,\u2_Display/n6323 }),
    .b({\u2_Display/n6320 ,\u2_Display/n6322 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add158/c23 ),
    .f({\u2_Display/n5191 [25],\u2_Display/n5191 [23]}),
    .fco(\u2_Display/add158/c27 ),
    .fx({\u2_Display/n5191 [26],\u2_Display/n5191 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u27_al_u4346  (
    .a({\u2_Display/n6317 ,\u2_Display/n6319 }),
    .b({\u2_Display/n6316 ,\u2_Display/n6318 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add158/c27 ),
    .f({\u2_Display/n5191 [29],\u2_Display/n5191 [27]}),
    .fco(\u2_Display/add158/c31 ),
    .fx({\u2_Display/n5191 [30],\u2_Display/n5191 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u31_al_u4347  (
    .a({open_n9384,\u2_Display/n6315 }),
    .c(2'b00),
    .d({open_n9389,1'b1}),
    .fci(\u2_Display/add158/c31 ),
    .f({open_n9406,\u2_Display/n5191 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u3_al_u4340  (
    .a({\u2_Display/n6341 ,\u2_Display/n6343 }),
    .b({\u2_Display/n6340 ,\u2_Display/n6342 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add158/c3 ),
    .f({\u2_Display/n5191 [5],\u2_Display/n5191 [3]}),
    .fco(\u2_Display/add158/c7 ),
    .fx({\u2_Display/n5191 [6],\u2_Display/n5191 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/u7_al_u4341  (
    .a({\u2_Display/n6337 ,\u2_Display/n6339 }),
    .b({\u2_Display/n6336 ,\u2_Display/n6338 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add158/c7 ),
    .f({\u2_Display/n5191 [9],\u2_Display/n5191 [7]}),
    .fco(\u2_Display/add158/c11 ),
    .fx({\u2_Display/n5191 [10],\u2_Display/n5191 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add158/ucin_al_u4339"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add158/ucin_al_u4339  (
    .a({\u2_Display/n6345 ,1'b1}),
    .b({\u2_Display/n6344 ,\u2_Display/n6346 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5191 [1],open_n9465}),
    .fco(\u2_Display/add158/c3 ),
    .fx({\u2_Display/n5191 [2],\u2_Display/n5191 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u11_al_u4351  (
    .a({\u2_Display/n5210 ,\u2_Display/n5212 }),
    .b({\u2_Display/n5209 ,\u2_Display/n5211 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add159/c11 ),
    .f({\u2_Display/n5226 [13],\u2_Display/n5226 [11]}),
    .fco(\u2_Display/add159/c15 ),
    .fx({\u2_Display/n5226 [14],\u2_Display/n5226 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u15_al_u4352  (
    .a({\u2_Display/n5206 ,\u2_Display/n5208 }),
    .b({\u2_Display/n5205 ,\u2_Display/n5207 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add159/c15 ),
    .f({\u2_Display/n5226 [17],\u2_Display/n5226 [15]}),
    .fco(\u2_Display/add159/c19 ),
    .fx({\u2_Display/n5226 [18],\u2_Display/n5226 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u19_al_u4353  (
    .a({\u2_Display/n5202 ,\u2_Display/n5204 }),
    .b({\u2_Display/n5201 ,\u2_Display/n5203 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add159/c19 ),
    .f({\u2_Display/n5226 [21],\u2_Display/n5226 [19]}),
    .fco(\u2_Display/add159/c23 ),
    .fx({\u2_Display/n5226 [22],\u2_Display/n5226 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u23_al_u4354  (
    .a({\u2_Display/n5198 ,\u2_Display/n5200 }),
    .b({\u2_Display/n5197 ,\u2_Display/n5199 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add159/c23 ),
    .f({\u2_Display/n5226 [25],\u2_Display/n5226 [23]}),
    .fco(\u2_Display/add159/c27 ),
    .fx({\u2_Display/n5226 [26],\u2_Display/n5226 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u27_al_u4355  (
    .a({\u2_Display/n6352 ,\u2_Display/n5196 }),
    .b({\u2_Display/n6351 ,\u2_Display/n6353 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add159/c27 ),
    .f({\u2_Display/n5226 [29],\u2_Display/n5226 [27]}),
    .fco(\u2_Display/add159/c31 ),
    .fx({\u2_Display/n5226 [30],\u2_Display/n5226 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u31_al_u4356  (
    .a({open_n9558,\u2_Display/n6350 }),
    .c(2'b00),
    .d({open_n9563,1'b1}),
    .fci(\u2_Display/add159/c31 ),
    .f({open_n9580,\u2_Display/n5226 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u3_al_u4349  (
    .a({\u2_Display/n5218 ,\u2_Display/n5220 }),
    .b({\u2_Display/n5217 ,\u2_Display/n5219 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add159/c3 ),
    .f({\u2_Display/n5226 [5],\u2_Display/n5226 [3]}),
    .fco(\u2_Display/add159/c7 ),
    .fx({\u2_Display/n5226 [6],\u2_Display/n5226 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/u7_al_u4350  (
    .a({\u2_Display/n5214 ,\u2_Display/n5216 }),
    .b({\u2_Display/n5213 ,\u2_Display/n5215 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add159/c7 ),
    .f({\u2_Display/n5226 [9],\u2_Display/n5226 [7]}),
    .fco(\u2_Display/add159/c11 ),
    .fx({\u2_Display/n5226 [10],\u2_Display/n5226 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add159/ucin_al_u4348"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add159/ucin_al_u4348  (
    .a({\u2_Display/n5222 ,1'b1}),
    .b({\u2_Display/n5221 ,\u2_Display/n5223 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5226 [1],open_n9639}),
    .fco(\u2_Display/add159/c3 ),
    .fx({\u2_Display/n5226 [2],\u2_Display/n5226 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u11_al_u4360  (
    .a({\u2_Display/n5245 ,\u2_Display/n5247 }),
    .b({\u2_Display/n5244 ,\u2_Display/n5246 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add160/c11 ),
    .f({\u2_Display/n5261 [13],\u2_Display/n5261 [11]}),
    .fco(\u2_Display/add160/c15 ),
    .fx({\u2_Display/n5261 [14],\u2_Display/n5261 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u15_al_u4361  (
    .a({\u2_Display/n5241 ,\u2_Display/n5243 }),
    .b({\u2_Display/n5240 ,\u2_Display/n5242 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add160/c15 ),
    .f({\u2_Display/n5261 [17],\u2_Display/n5261 [15]}),
    .fco(\u2_Display/add160/c19 ),
    .fx({\u2_Display/n5261 [18],\u2_Display/n5261 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u19_al_u4362  (
    .a({\u2_Display/n5237 ,\u2_Display/n5239 }),
    .b({\u2_Display/n5236 ,\u2_Display/n5238 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add160/c19 ),
    .f({\u2_Display/n5261 [21],\u2_Display/n5261 [19]}),
    .fco(\u2_Display/add160/c23 ),
    .fx({\u2_Display/n5261 [22],\u2_Display/n5261 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u23_al_u4363  (
    .a({\u2_Display/n5233 ,\u2_Display/n5235 }),
    .b({\u2_Display/n5232 ,\u2_Display/n5234 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add160/c23 ),
    .f({\u2_Display/n5261 [25],\u2_Display/n5261 [23]}),
    .fco(\u2_Display/add160/c27 ),
    .fx({\u2_Display/n5261 [26],\u2_Display/n5261 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u27_al_u4364  (
    .a({\u2_Display/n5229 ,\u2_Display/n5231 }),
    .b({\u2_Display/n5228 ,\u2_Display/n5230 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add160/c27 ),
    .f({\u2_Display/n5261 [29],\u2_Display/n5261 [27]}),
    .fco(\u2_Display/add160/c31 ),
    .fx({\u2_Display/n5261 [30],\u2_Display/n5261 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u31_al_u4365  (
    .a({open_n9732,\u2_Display/n5227 }),
    .c(2'b00),
    .d({open_n9737,1'b1}),
    .fci(\u2_Display/add160/c31 ),
    .f({open_n9754,\u2_Display/n5261 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u3_al_u4358  (
    .a({\u2_Display/n5253 ,\u2_Display/n5255 }),
    .b({\u2_Display/n5252 ,\u2_Display/n5254 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add160/c3 ),
    .f({\u2_Display/n5261 [5],\u2_Display/n5261 [3]}),
    .fco(\u2_Display/add160/c7 ),
    .fx({\u2_Display/n5261 [6],\u2_Display/n5261 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/u7_al_u4359  (
    .a({\u2_Display/n5249 ,\u2_Display/n5251 }),
    .b({\u2_Display/n5248 ,\u2_Display/n5250 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add160/c7 ),
    .f({\u2_Display/n5261 [9],\u2_Display/n5261 [7]}),
    .fco(\u2_Display/add160/c11 ),
    .fx({\u2_Display/n5261 [10],\u2_Display/n5261 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add160/ucin_al_u4357"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add160/ucin_al_u4357  (
    .a({\u2_Display/n5257 ,1'b1}),
    .b({\u2_Display/n5256 ,\u2_Display/n5258 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5261 [1],open_n9813}),
    .fco(\u2_Display/add160/c3 ),
    .fx({\u2_Display/n5261 [2],\u2_Display/n5261 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u11_al_u4369  (
    .a({\u2_Display/n5280 ,\u2_Display/n5282 }),
    .b({\u2_Display/n5279 ,\u2_Display/n5281 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add161/c11 ),
    .f({\u2_Display/n5296 [13],\u2_Display/n5296 [11]}),
    .fco(\u2_Display/add161/c15 ),
    .fx({\u2_Display/n5296 [14],\u2_Display/n5296 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u15_al_u4370  (
    .a({\u2_Display/n5276 ,\u2_Display/n5278 }),
    .b({\u2_Display/n5275 ,\u2_Display/n5277 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add161/c15 ),
    .f({\u2_Display/n5296 [17],\u2_Display/n5296 [15]}),
    .fco(\u2_Display/add161/c19 ),
    .fx({\u2_Display/n5296 [18],\u2_Display/n5296 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u19_al_u4371  (
    .a({\u2_Display/n5272 ,\u2_Display/n5274 }),
    .b({\u2_Display/n5271 ,\u2_Display/n5273 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add161/c19 ),
    .f({\u2_Display/n5296 [21],\u2_Display/n5296 [19]}),
    .fco(\u2_Display/add161/c23 ),
    .fx({\u2_Display/n5296 [22],\u2_Display/n5296 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u23_al_u4372  (
    .a({\u2_Display/n5268 ,\u2_Display/n5270 }),
    .b({\u2_Display/n5267 ,\u2_Display/n5269 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add161/c23 ),
    .f({\u2_Display/n5296 [25],\u2_Display/n5296 [23]}),
    .fco(\u2_Display/add161/c27 ),
    .fx({\u2_Display/n5296 [26],\u2_Display/n5296 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u27_al_u4373  (
    .a({\u2_Display/n5264 ,\u2_Display/n5266 }),
    .b({\u2_Display/n5263 ,\u2_Display/n5265 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add161/c27 ),
    .f({\u2_Display/n5296 [29],\u2_Display/n5296 [27]}),
    .fco(\u2_Display/add161/c31 ),
    .fx({\u2_Display/n5296 [30],\u2_Display/n5296 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u31_al_u4374  (
    .a({open_n9906,\u2_Display/n5262 }),
    .c(2'b00),
    .d({open_n9911,1'b1}),
    .fci(\u2_Display/add161/c31 ),
    .f({open_n9928,\u2_Display/n5296 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u3_al_u4367  (
    .a({\u2_Display/n5288 ,\u2_Display/n5290 }),
    .b({\u2_Display/n5287 ,\u2_Display/n5289 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add161/c3 ),
    .f({\u2_Display/n5296 [5],\u2_Display/n5296 [3]}),
    .fco(\u2_Display/add161/c7 ),
    .fx({\u2_Display/n5296 [6],\u2_Display/n5296 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/u7_al_u4368  (
    .a({\u2_Display/n5284 ,\u2_Display/n5286 }),
    .b({\u2_Display/n5283 ,\u2_Display/n5285 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add161/c7 ),
    .f({\u2_Display/n5296 [9],\u2_Display/n5296 [7]}),
    .fco(\u2_Display/add161/c11 ),
    .fx({\u2_Display/n5296 [10],\u2_Display/n5296 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add161/ucin_al_u4366"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add161/ucin_al_u4366  (
    .a({\u2_Display/n5292 ,1'b1}),
    .b({\u2_Display/n5291 ,\u2_Display/n5293 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5296 [1],open_n9987}),
    .fco(\u2_Display/add161/c3 ),
    .fx({\u2_Display/n5296 [2],\u2_Display/n5296 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u11_al_u4378  (
    .a({\u2_Display/n5315 ,\u2_Display/n5317 }),
    .b({\u2_Display/n5314 ,\u2_Display/n5316 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add162/c11 ),
    .f({\u2_Display/n5331 [13],\u2_Display/n5331 [11]}),
    .fco(\u2_Display/add162/c15 ),
    .fx({\u2_Display/n5331 [14],\u2_Display/n5331 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u15_al_u4379  (
    .a({\u2_Display/n5311 ,\u2_Display/n5313 }),
    .b({\u2_Display/n5310 ,\u2_Display/n5312 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add162/c15 ),
    .f({\u2_Display/n5331 [17],\u2_Display/n5331 [15]}),
    .fco(\u2_Display/add162/c19 ),
    .fx({\u2_Display/n5331 [18],\u2_Display/n5331 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u19_al_u4380  (
    .a({\u2_Display/n5307 ,\u2_Display/n5309 }),
    .b({\u2_Display/n5306 ,\u2_Display/n5308 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add162/c19 ),
    .f({\u2_Display/n5331 [21],\u2_Display/n5331 [19]}),
    .fco(\u2_Display/add162/c23 ),
    .fx({\u2_Display/n5331 [22],\u2_Display/n5331 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u23_al_u4381  (
    .a({\u2_Display/n5303 ,\u2_Display/n5305 }),
    .b({\u2_Display/n5302 ,\u2_Display/n5304 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add162/c23 ),
    .f({\u2_Display/n5331 [25],\u2_Display/n5331 [23]}),
    .fco(\u2_Display/add162/c27 ),
    .fx({\u2_Display/n5331 [26],\u2_Display/n5331 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u27_al_u4382  (
    .a({\u2_Display/n5299 ,\u2_Display/n5301 }),
    .b({\u2_Display/n5298 ,\u2_Display/n5300 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add162/c27 ),
    .f({\u2_Display/n5331 [29],\u2_Display/n5331 [27]}),
    .fco(\u2_Display/add162/c31 ),
    .fx({\u2_Display/n5331 [30],\u2_Display/n5331 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u31_al_u4383  (
    .a({open_n10080,\u2_Display/n5297 }),
    .c(2'b00),
    .d({open_n10085,1'b1}),
    .fci(\u2_Display/add162/c31 ),
    .f({open_n10102,\u2_Display/n5331 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u3_al_u4376  (
    .a({\u2_Display/n5323 ,\u2_Display/n5325 }),
    .b({\u2_Display/n5322 ,\u2_Display/n5324 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add162/c3 ),
    .f({\u2_Display/n5331 [5],\u2_Display/n5331 [3]}),
    .fco(\u2_Display/add162/c7 ),
    .fx({\u2_Display/n5331 [6],\u2_Display/n5331 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/u7_al_u4377  (
    .a({\u2_Display/n5319 ,\u2_Display/n5321 }),
    .b({\u2_Display/n5318 ,\u2_Display/n5320 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add162/c7 ),
    .f({\u2_Display/n5331 [9],\u2_Display/n5331 [7]}),
    .fco(\u2_Display/add162/c11 ),
    .fx({\u2_Display/n5331 [10],\u2_Display/n5331 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add162/ucin_al_u4375"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add162/ucin_al_u4375  (
    .a({\u2_Display/n5327 ,1'b1}),
    .b({\u2_Display/n5326 ,\u2_Display/n5328 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5331 [1],open_n10161}),
    .fco(\u2_Display/add162/c3 ),
    .fx({\u2_Display/n5331 [2],\u2_Display/n5331 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u11_al_u4387  (
    .a({\u2_Display/n5350 ,\u2_Display/n5352 }),
    .b({\u2_Display/n5349 ,\u2_Display/n5351 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add163/c11 ),
    .f({\u2_Display/n5366 [13],\u2_Display/n5366 [11]}),
    .fco(\u2_Display/add163/c15 ),
    .fx({\u2_Display/n5366 [14],\u2_Display/n5366 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u15_al_u4388  (
    .a({\u2_Display/n5346 ,\u2_Display/n5348 }),
    .b({\u2_Display/n5345 ,\u2_Display/n5347 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add163/c15 ),
    .f({\u2_Display/n5366 [17],\u2_Display/n5366 [15]}),
    .fco(\u2_Display/add163/c19 ),
    .fx({\u2_Display/n5366 [18],\u2_Display/n5366 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u19_al_u4389  (
    .a({\u2_Display/n5342 ,\u2_Display/n5344 }),
    .b({\u2_Display/n5341 ,\u2_Display/n5343 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add163/c19 ),
    .f({\u2_Display/n5366 [21],\u2_Display/n5366 [19]}),
    .fco(\u2_Display/add163/c23 ),
    .fx({\u2_Display/n5366 [22],\u2_Display/n5366 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u23_al_u4390  (
    .a({\u2_Display/n5338 ,\u2_Display/n5340 }),
    .b({\u2_Display/n5337 ,\u2_Display/n5339 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add163/c23 ),
    .f({\u2_Display/n5366 [25],\u2_Display/n5366 [23]}),
    .fco(\u2_Display/add163/c27 ),
    .fx({\u2_Display/n5366 [26],\u2_Display/n5366 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u27_al_u4391  (
    .a({\u2_Display/n5334 ,\u2_Display/n5336 }),
    .b({\u2_Display/n5333 ,\u2_Display/n5335 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add163/c27 ),
    .f({\u2_Display/n5366 [29],\u2_Display/n5366 [27]}),
    .fco(\u2_Display/add163/c31 ),
    .fx({\u2_Display/n5366 [30],\u2_Display/n5366 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u31_al_u4392  (
    .a({open_n10254,\u2_Display/n5332 }),
    .c(2'b00),
    .d({open_n10259,1'b1}),
    .fci(\u2_Display/add163/c31 ),
    .f({open_n10276,\u2_Display/n5366 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u3_al_u4385  (
    .a({\u2_Display/n5358 ,\u2_Display/n5360 }),
    .b({\u2_Display/n5357 ,\u2_Display/n5359 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add163/c3 ),
    .f({\u2_Display/n5366 [5],\u2_Display/n5366 [3]}),
    .fco(\u2_Display/add163/c7 ),
    .fx({\u2_Display/n5366 [6],\u2_Display/n5366 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/u7_al_u4386  (
    .a({\u2_Display/n5354 ,\u2_Display/n5356 }),
    .b({\u2_Display/n5353 ,\u2_Display/n5355 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add163/c7 ),
    .f({\u2_Display/n5366 [9],\u2_Display/n5366 [7]}),
    .fco(\u2_Display/add163/c11 ),
    .fx({\u2_Display/n5366 [10],\u2_Display/n5366 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add163/ucin_al_u4384"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add163/ucin_al_u4384  (
    .a({\u2_Display/n5362 ,1'b1}),
    .b({\u2_Display/n5361 ,\u2_Display/n5363 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5366 [1],open_n10335}),
    .fco(\u2_Display/add163/c3 ),
    .fx({\u2_Display/n5366 [2],\u2_Display/n5366 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u11_al_u4396  (
    .a({\u2_Display/n5385 ,\u2_Display/n5387 }),
    .b({\u2_Display/n5384 ,\u2_Display/n5386 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add164/c11 ),
    .f({\u2_Display/n5401 [13],\u2_Display/n5401 [11]}),
    .fco(\u2_Display/add164/c15 ),
    .fx({\u2_Display/n5401 [14],\u2_Display/n5401 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u15_al_u4397  (
    .a({\u2_Display/n5381 ,\u2_Display/n5383 }),
    .b({\u2_Display/n5380 ,\u2_Display/n5382 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add164/c15 ),
    .f({\u2_Display/n5401 [17],\u2_Display/n5401 [15]}),
    .fco(\u2_Display/add164/c19 ),
    .fx({\u2_Display/n5401 [18],\u2_Display/n5401 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u19_al_u4398  (
    .a({\u2_Display/n5377 ,\u2_Display/n5379 }),
    .b({\u2_Display/n5376 ,\u2_Display/n5378 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add164/c19 ),
    .f({\u2_Display/n5401 [21],\u2_Display/n5401 [19]}),
    .fco(\u2_Display/add164/c23 ),
    .fx({\u2_Display/n5401 [22],\u2_Display/n5401 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u23_al_u4399  (
    .a({\u2_Display/n5373 ,\u2_Display/n5375 }),
    .b({\u2_Display/n5372 ,\u2_Display/n5374 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add164/c23 ),
    .f({\u2_Display/n5401 [25],\u2_Display/n5401 [23]}),
    .fco(\u2_Display/add164/c27 ),
    .fx({\u2_Display/n5401 [26],\u2_Display/n5401 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u27_al_u4400  (
    .a({\u2_Display/n5369 ,\u2_Display/n5371 }),
    .b({\u2_Display/n5368 ,\u2_Display/n5370 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add164/c27 ),
    .f({\u2_Display/n5401 [29],\u2_Display/n5401 [27]}),
    .fco(\u2_Display/add164/c31 ),
    .fx({\u2_Display/n5401 [30],\u2_Display/n5401 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u31_al_u4401  (
    .a({open_n10428,\u2_Display/n5367 }),
    .c(2'b00),
    .d({open_n10433,1'b1}),
    .fci(\u2_Display/add164/c31 ),
    .f({open_n10450,\u2_Display/n5401 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u3_al_u4394  (
    .a({\u2_Display/n5393 ,\u2_Display/n5395 }),
    .b({\u2_Display/n5392 ,\u2_Display/n5394 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add164/c3 ),
    .f({\u2_Display/n5401 [5],\u2_Display/n5401 [3]}),
    .fco(\u2_Display/add164/c7 ),
    .fx({\u2_Display/n5401 [6],\u2_Display/n5401 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/u7_al_u4395  (
    .a({\u2_Display/n5389 ,\u2_Display/n5391 }),
    .b({\u2_Display/n5388 ,\u2_Display/n5390 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add164/c7 ),
    .f({\u2_Display/n5401 [9],\u2_Display/n5401 [7]}),
    .fco(\u2_Display/add164/c11 ),
    .fx({\u2_Display/n5401 [10],\u2_Display/n5401 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add164/ucin_al_u4393"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add164/ucin_al_u4393  (
    .a({\u2_Display/n5397 ,1'b1}),
    .b({\u2_Display/n5396 ,\u2_Display/n5398 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5401 [1],open_n10509}),
    .fco(\u2_Display/add164/c3 ),
    .fx({\u2_Display/n5401 [2],\u2_Display/n5401 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u11_al_u4405  (
    .a({\u2_Display/n5420 ,\u2_Display/n5422 }),
    .b({\u2_Display/n5419 ,\u2_Display/n5421 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add165/c11 ),
    .f({\u2_Display/n5436 [13],\u2_Display/n5436 [11]}),
    .fco(\u2_Display/add165/c15 ),
    .fx({\u2_Display/n5436 [14],\u2_Display/n5436 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u15_al_u4406  (
    .a({\u2_Display/n5416 ,\u2_Display/n5418 }),
    .b({\u2_Display/n5415 ,\u2_Display/n5417 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add165/c15 ),
    .f({\u2_Display/n5436 [17],\u2_Display/n5436 [15]}),
    .fco(\u2_Display/add165/c19 ),
    .fx({\u2_Display/n5436 [18],\u2_Display/n5436 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u19_al_u4407  (
    .a({\u2_Display/n5412 ,\u2_Display/n5414 }),
    .b({\u2_Display/n5411 ,\u2_Display/n5413 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add165/c19 ),
    .f({\u2_Display/n5436 [21],\u2_Display/n5436 [19]}),
    .fco(\u2_Display/add165/c23 ),
    .fx({\u2_Display/n5436 [22],\u2_Display/n5436 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u23_al_u4408  (
    .a({\u2_Display/n5408 ,\u2_Display/n5410 }),
    .b({\u2_Display/n5407 ,\u2_Display/n5409 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add165/c23 ),
    .f({\u2_Display/n5436 [25],\u2_Display/n5436 [23]}),
    .fco(\u2_Display/add165/c27 ),
    .fx({\u2_Display/n5436 [26],\u2_Display/n5436 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u27_al_u4409  (
    .a({\u2_Display/n5404 ,\u2_Display/n5406 }),
    .b({\u2_Display/n5403 ,\u2_Display/n5405 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add165/c27 ),
    .f({\u2_Display/n5436 [29],\u2_Display/n5436 [27]}),
    .fco(\u2_Display/add165/c31 ),
    .fx({\u2_Display/n5436 [30],\u2_Display/n5436 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u31_al_u4410  (
    .a({open_n10602,\u2_Display/n5402 }),
    .c(2'b00),
    .d({open_n10607,1'b1}),
    .fci(\u2_Display/add165/c31 ),
    .f({open_n10624,\u2_Display/n5436 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u3_al_u4403  (
    .a({\u2_Display/n5428 ,\u2_Display/n5430 }),
    .b({\u2_Display/n5427 ,\u2_Display/n5429 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add165/c3 ),
    .f({\u2_Display/n5436 [5],\u2_Display/n5436 [3]}),
    .fco(\u2_Display/add165/c7 ),
    .fx({\u2_Display/n5436 [6],\u2_Display/n5436 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/u7_al_u4404  (
    .a({\u2_Display/n5424 ,\u2_Display/n5426 }),
    .b({\u2_Display/n5423 ,\u2_Display/n5425 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add165/c7 ),
    .f({\u2_Display/n5436 [9],\u2_Display/n5436 [7]}),
    .fco(\u2_Display/add165/c11 ),
    .fx({\u2_Display/n5436 [10],\u2_Display/n5436 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add165/ucin_al_u4402"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add165/ucin_al_u4402  (
    .a({\u2_Display/n5432 ,1'b1}),
    .b({\u2_Display/n5431 ,\u2_Display/n5433 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5436 [1],open_n10683}),
    .fco(\u2_Display/add165/c3 ),
    .fx({\u2_Display/n5436 [2],\u2_Display/n5436 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u11_al_u4414  (
    .a({\u2_Display/n5455 ,\u2_Display/n5457 }),
    .b({\u2_Display/n5454 ,\u2_Display/n5456 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add166/c11 ),
    .f({\u2_Display/n5471 [13],\u2_Display/n5471 [11]}),
    .fco(\u2_Display/add166/c15 ),
    .fx({\u2_Display/n5471 [14],\u2_Display/n5471 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u15_al_u4415  (
    .a({\u2_Display/n5451 ,\u2_Display/n5453 }),
    .b({\u2_Display/n5450 ,\u2_Display/n5452 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add166/c15 ),
    .f({\u2_Display/n5471 [17],\u2_Display/n5471 [15]}),
    .fco(\u2_Display/add166/c19 ),
    .fx({\u2_Display/n5471 [18],\u2_Display/n5471 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u19_al_u4416  (
    .a({\u2_Display/n5447 ,\u2_Display/n5449 }),
    .b({\u2_Display/n5446 ,\u2_Display/n5448 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add166/c19 ),
    .f({\u2_Display/n5471 [21],\u2_Display/n5471 [19]}),
    .fco(\u2_Display/add166/c23 ),
    .fx({\u2_Display/n5471 [22],\u2_Display/n5471 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u23_al_u4417  (
    .a({\u2_Display/n5443 ,\u2_Display/n5445 }),
    .b({\u2_Display/n5442 ,\u2_Display/n5444 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add166/c23 ),
    .f({\u2_Display/n5471 [25],\u2_Display/n5471 [23]}),
    .fco(\u2_Display/add166/c27 ),
    .fx({\u2_Display/n5471 [26],\u2_Display/n5471 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u27_al_u4418  (
    .a({\u2_Display/n5439 ,\u2_Display/n5441 }),
    .b({\u2_Display/n5438 ,\u2_Display/n5440 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add166/c27 ),
    .f({\u2_Display/n5471 [29],\u2_Display/n5471 [27]}),
    .fco(\u2_Display/add166/c31 ),
    .fx({\u2_Display/n5471 [30],\u2_Display/n5471 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u31_al_u4419  (
    .a({open_n10776,\u2_Display/n5437 }),
    .c(2'b00),
    .d({open_n10781,1'b1}),
    .fci(\u2_Display/add166/c31 ),
    .f({open_n10798,\u2_Display/n5471 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u3_al_u4412  (
    .a({\u2_Display/n5463 ,\u2_Display/n5465 }),
    .b({\u2_Display/n5462 ,\u2_Display/n5464 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add166/c3 ),
    .f({\u2_Display/n5471 [5],\u2_Display/n5471 [3]}),
    .fco(\u2_Display/add166/c7 ),
    .fx({\u2_Display/n5471 [6],\u2_Display/n5471 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/u7_al_u4413  (
    .a({\u2_Display/n5459 ,\u2_Display/n5461 }),
    .b({\u2_Display/n5458 ,\u2_Display/n5460 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add166/c7 ),
    .f({\u2_Display/n5471 [9],\u2_Display/n5471 [7]}),
    .fco(\u2_Display/add166/c11 ),
    .fx({\u2_Display/n5471 [10],\u2_Display/n5471 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add166/ucin_al_u4411"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add166/ucin_al_u4411  (
    .a({\u2_Display/n5467 ,1'b1}),
    .b({\u2_Display/n5466 ,\u2_Display/n5468 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5471 [1],open_n10857}),
    .fco(\u2_Display/add166/c3 ),
    .fx({\u2_Display/n5471 [2],\u2_Display/n5471 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u11_al_u4423  (
    .a({\u2_Display/n5490 ,\u2_Display/n5492 }),
    .b({\u2_Display/n5489 ,\u2_Display/n5491 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add167/c11 ),
    .f({\u2_Display/n5506 [13],\u2_Display/n5506 [11]}),
    .fco(\u2_Display/add167/c15 ),
    .fx({\u2_Display/n5506 [14],\u2_Display/n5506 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u15_al_u4424  (
    .a({\u2_Display/n5486 ,\u2_Display/n5488 }),
    .b({\u2_Display/n5485 ,\u2_Display/n5487 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add167/c15 ),
    .f({\u2_Display/n5506 [17],\u2_Display/n5506 [15]}),
    .fco(\u2_Display/add167/c19 ),
    .fx({\u2_Display/n5506 [18],\u2_Display/n5506 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u19_al_u4425  (
    .a({\u2_Display/n5482 ,\u2_Display/n5484 }),
    .b({\u2_Display/n5481 ,\u2_Display/n5483 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add167/c19 ),
    .f({\u2_Display/n5506 [21],\u2_Display/n5506 [19]}),
    .fco(\u2_Display/add167/c23 ),
    .fx({\u2_Display/n5506 [22],\u2_Display/n5506 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u23_al_u4426  (
    .a({\u2_Display/n5478 ,\u2_Display/n5480 }),
    .b({\u2_Display/n5477 ,\u2_Display/n5479 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add167/c23 ),
    .f({\u2_Display/n5506 [25],\u2_Display/n5506 [23]}),
    .fco(\u2_Display/add167/c27 ),
    .fx({\u2_Display/n5506 [26],\u2_Display/n5506 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u27_al_u4427  (
    .a({\u2_Display/n5474 ,\u2_Display/n5476 }),
    .b({\u2_Display/n5473 ,\u2_Display/n5475 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add167/c27 ),
    .f({\u2_Display/n5506 [29],\u2_Display/n5506 [27]}),
    .fco(\u2_Display/add167/c31 ),
    .fx({\u2_Display/n5506 [30],\u2_Display/n5506 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u31_al_u4428  (
    .a({open_n10950,\u2_Display/n5472 }),
    .c(2'b00),
    .d({open_n10955,1'b1}),
    .fci(\u2_Display/add167/c31 ),
    .f({open_n10972,\u2_Display/n5506 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u3_al_u4421  (
    .a({\u2_Display/n5498 ,\u2_Display/n5500 }),
    .b({\u2_Display/n5497 ,\u2_Display/n5499 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add167/c3 ),
    .f({\u2_Display/n5506 [5],\u2_Display/n5506 [3]}),
    .fco(\u2_Display/add167/c7 ),
    .fx({\u2_Display/n5506 [6],\u2_Display/n5506 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/u7_al_u4422  (
    .a({\u2_Display/n5494 ,\u2_Display/n5496 }),
    .b({\u2_Display/n5493 ,\u2_Display/n5495 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add167/c7 ),
    .f({\u2_Display/n5506 [9],\u2_Display/n5506 [7]}),
    .fco(\u2_Display/add167/c11 ),
    .fx({\u2_Display/n5506 [10],\u2_Display/n5506 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add167/ucin_al_u4420"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add167/ucin_al_u4420  (
    .a({\u2_Display/n5502 ,1'b1}),
    .b({\u2_Display/n5501 ,\u2_Display/n5503 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5506 [1],open_n11031}),
    .fco(\u2_Display/add167/c3 ),
    .fx({\u2_Display/n5506 [2],\u2_Display/n5506 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u11_al_u4432  (
    .a({\u2_Display/n5525 ,\u2_Display/n5527 }),
    .b({\u2_Display/n5524 ,\u2_Display/n5526 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add168/c11 ),
    .f({\u2_Display/n5541 [13],\u2_Display/n5541 [11]}),
    .fco(\u2_Display/add168/c15 ),
    .fx({\u2_Display/n5541 [14],\u2_Display/n5541 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u15_al_u4433  (
    .a({\u2_Display/n5521 ,\u2_Display/n5523 }),
    .b({\u2_Display/n5520 ,\u2_Display/n5522 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add168/c15 ),
    .f({\u2_Display/n5541 [17],\u2_Display/n5541 [15]}),
    .fco(\u2_Display/add168/c19 ),
    .fx({\u2_Display/n5541 [18],\u2_Display/n5541 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u19_al_u4434  (
    .a({\u2_Display/n5517 ,\u2_Display/n5519 }),
    .b({\u2_Display/n5516 ,\u2_Display/n5518 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add168/c19 ),
    .f({\u2_Display/n5541 [21],\u2_Display/n5541 [19]}),
    .fco(\u2_Display/add168/c23 ),
    .fx({\u2_Display/n5541 [22],\u2_Display/n5541 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u23_al_u4435  (
    .a({\u2_Display/n5513 ,\u2_Display/n5515 }),
    .b({\u2_Display/n5512 ,\u2_Display/n5514 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add168/c23 ),
    .f({\u2_Display/n5541 [25],\u2_Display/n5541 [23]}),
    .fco(\u2_Display/add168/c27 ),
    .fx({\u2_Display/n5541 [26],\u2_Display/n5541 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u27_al_u4436  (
    .a({\u2_Display/n5509 ,\u2_Display/n5511 }),
    .b({\u2_Display/n5508 ,\u2_Display/n5510 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add168/c27 ),
    .f({\u2_Display/n5541 [29],\u2_Display/n5541 [27]}),
    .fco(\u2_Display/add168/c31 ),
    .fx({\u2_Display/n5541 [30],\u2_Display/n5541 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u31_al_u4437  (
    .a({open_n11124,\u2_Display/n5507 }),
    .c(2'b00),
    .d({open_n11129,1'b1}),
    .fci(\u2_Display/add168/c31 ),
    .f({open_n11146,\u2_Display/n5541 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u3_al_u4430  (
    .a({\u2_Display/n5533 ,\u2_Display/n5535 }),
    .b({\u2_Display/n5532 ,\u2_Display/n5534 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add168/c3 ),
    .f({\u2_Display/n5541 [5],\u2_Display/n5541 [3]}),
    .fco(\u2_Display/add168/c7 ),
    .fx({\u2_Display/n5541 [6],\u2_Display/n5541 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/u7_al_u4431  (
    .a({\u2_Display/n5529 ,\u2_Display/n5531 }),
    .b({\u2_Display/n5528 ,\u2_Display/n5530 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add168/c7 ),
    .f({\u2_Display/n5541 [9],\u2_Display/n5541 [7]}),
    .fco(\u2_Display/add168/c11 ),
    .fx({\u2_Display/n5541 [10],\u2_Display/n5541 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add168/ucin_al_u4429"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add168/ucin_al_u4429  (
    .a({\u2_Display/n5537 ,1'b1}),
    .b({\u2_Display/n5536 ,\u2_Display/n5538 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5541 [1],open_n11205}),
    .fco(\u2_Display/add168/c3 ),
    .fx({\u2_Display/n5541 [2],\u2_Display/n5541 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u11_al_u4441  (
    .a({\u2_Display/n5560 ,\u2_Display/n5562 }),
    .b({\u2_Display/n5559 ,\u2_Display/n5561 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add169/c11 ),
    .f({\u2_Display/n5576 [13],\u2_Display/n5576 [11]}),
    .fco(\u2_Display/add169/c15 ),
    .fx({\u2_Display/n5576 [14],\u2_Display/n5576 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u15_al_u4442  (
    .a({\u2_Display/n5556 ,\u2_Display/n5558 }),
    .b({\u2_Display/n5555 ,\u2_Display/n5557 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add169/c15 ),
    .f({\u2_Display/n5576 [17],\u2_Display/n5576 [15]}),
    .fco(\u2_Display/add169/c19 ),
    .fx({\u2_Display/n5576 [18],\u2_Display/n5576 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u19_al_u4443  (
    .a({\u2_Display/n5552 ,\u2_Display/n5554 }),
    .b({\u2_Display/n5551 ,\u2_Display/n5553 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add169/c19 ),
    .f({\u2_Display/n5576 [21],\u2_Display/n5576 [19]}),
    .fco(\u2_Display/add169/c23 ),
    .fx({\u2_Display/n5576 [22],\u2_Display/n5576 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u23_al_u4444  (
    .a({\u2_Display/n5548 ,\u2_Display/n5550 }),
    .b({\u2_Display/n5547 ,\u2_Display/n5549 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add169/c23 ),
    .f({\u2_Display/n5576 [25],\u2_Display/n5576 [23]}),
    .fco(\u2_Display/add169/c27 ),
    .fx({\u2_Display/n5576 [26],\u2_Display/n5576 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u27_al_u4445  (
    .a({\u2_Display/n5544 ,\u2_Display/n5546 }),
    .b({\u2_Display/n5543 ,\u2_Display/n5545 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add169/c27 ),
    .f({\u2_Display/n5576 [29],\u2_Display/n5576 [27]}),
    .fco(\u2_Display/add169/c31 ),
    .fx({\u2_Display/n5576 [30],\u2_Display/n5576 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u31_al_u4446  (
    .a({open_n11298,\u2_Display/n5542 }),
    .c(2'b00),
    .d({open_n11303,1'b1}),
    .fci(\u2_Display/add169/c31 ),
    .f({open_n11320,\u2_Display/n5576 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u3_al_u4439  (
    .a({\u2_Display/n5568 ,\u2_Display/n5570 }),
    .b({\u2_Display/n5567 ,\u2_Display/n5569 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add169/c3 ),
    .f({\u2_Display/n5576 [5],\u2_Display/n5576 [3]}),
    .fco(\u2_Display/add169/c7 ),
    .fx({\u2_Display/n5576 [6],\u2_Display/n5576 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/u7_al_u4440  (
    .a({\u2_Display/n5564 ,\u2_Display/n5566 }),
    .b({\u2_Display/n5563 ,\u2_Display/n5565 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add169/c7 ),
    .f({\u2_Display/n5576 [9],\u2_Display/n5576 [7]}),
    .fco(\u2_Display/add169/c11 ),
    .fx({\u2_Display/n5576 [10],\u2_Display/n5576 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add169/ucin_al_u4438"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add169/ucin_al_u4438  (
    .a({\u2_Display/n5572 ,1'b1}),
    .b({\u2_Display/n5571 ,\u2_Display/n5573 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5576 [1],open_n11379}),
    .fco(\u2_Display/add169/c3 ),
    .fx({\u2_Display/n5576 [2],\u2_Display/n5576 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u11_al_u4450  (
    .a({\u2_Display/n5595 ,\u2_Display/n5597 }),
    .b({\u2_Display/n5594 ,\u2_Display/n5596 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add170/c11 ),
    .f({\u2_Display/n5611 [13],\u2_Display/n5611 [11]}),
    .fco(\u2_Display/add170/c15 ),
    .fx({\u2_Display/n5611 [14],\u2_Display/n5611 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u15_al_u4451  (
    .a({\u2_Display/n5591 ,\u2_Display/n5593 }),
    .b({\u2_Display/n5590 ,\u2_Display/n5592 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add170/c15 ),
    .f({\u2_Display/n5611 [17],\u2_Display/n5611 [15]}),
    .fco(\u2_Display/add170/c19 ),
    .fx({\u2_Display/n5611 [18],\u2_Display/n5611 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u19_al_u4452  (
    .a({\u2_Display/n5587 ,\u2_Display/n5589 }),
    .b({\u2_Display/n5586 ,\u2_Display/n5588 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add170/c19 ),
    .f({\u2_Display/n5611 [21],\u2_Display/n5611 [19]}),
    .fco(\u2_Display/add170/c23 ),
    .fx({\u2_Display/n5611 [22],\u2_Display/n5611 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u23_al_u4453  (
    .a({\u2_Display/n5583 ,\u2_Display/n5585 }),
    .b({\u2_Display/n5582 ,\u2_Display/n5584 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add170/c23 ),
    .f({\u2_Display/n5611 [25],\u2_Display/n5611 [23]}),
    .fco(\u2_Display/add170/c27 ),
    .fx({\u2_Display/n5611 [26],\u2_Display/n5611 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u27_al_u4454  (
    .a({\u2_Display/n5579 ,\u2_Display/n5581 }),
    .b({\u2_Display/n5578 ,\u2_Display/n5580 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add170/c27 ),
    .f({\u2_Display/n5611 [29],\u2_Display/n5611 [27]}),
    .fco(\u2_Display/add170/c31 ),
    .fx({\u2_Display/n5611 [30],\u2_Display/n5611 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u31_al_u4455  (
    .a({open_n11472,\u2_Display/n5577 }),
    .c(2'b00),
    .d({open_n11477,1'b1}),
    .fci(\u2_Display/add170/c31 ),
    .f({open_n11494,\u2_Display/n5611 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u3_al_u4448  (
    .a({\u2_Display/n5603 ,\u2_Display/n5605 }),
    .b({\u2_Display/n5602 ,\u2_Display/n5604 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add170/c3 ),
    .f({\u2_Display/n5611 [5],\u2_Display/n5611 [3]}),
    .fco(\u2_Display/add170/c7 ),
    .fx({\u2_Display/n5611 [6],\u2_Display/n5611 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/u7_al_u4449  (
    .a({\u2_Display/n5599 ,\u2_Display/n5601 }),
    .b({\u2_Display/n5598 ,\u2_Display/n5600 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add170/c7 ),
    .f({\u2_Display/n5611 [9],\u2_Display/n5611 [7]}),
    .fco(\u2_Display/add170/c11 ),
    .fx({\u2_Display/n5611 [10],\u2_Display/n5611 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add170/ucin_al_u4447"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add170/ucin_al_u4447  (
    .a({\u2_Display/n5607 ,1'b1}),
    .b({\u2_Display/n5606 ,\u2_Display/n5608 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5611 [1],open_n11553}),
    .fco(\u2_Display/add170/c3 ),
    .fx({\u2_Display/n5611 [2],\u2_Display/n5611 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u11_al_u4459  (
    .a({\u2_Display/n5630 ,\u2_Display/n5632 }),
    .b({\u2_Display/n5629 ,\u2_Display/n5631 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add171/c11 ),
    .f({\u2_Display/n5646 [13],\u2_Display/n5646 [11]}),
    .fco(\u2_Display/add171/c15 ),
    .fx({\u2_Display/n5646 [14],\u2_Display/n5646 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u15_al_u4460  (
    .a({\u2_Display/n5626 ,\u2_Display/n5628 }),
    .b({\u2_Display/n5625 ,\u2_Display/n5627 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add171/c15 ),
    .f({\u2_Display/n5646 [17],\u2_Display/n5646 [15]}),
    .fco(\u2_Display/add171/c19 ),
    .fx({\u2_Display/n5646 [18],\u2_Display/n5646 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u19_al_u4461  (
    .a({\u2_Display/n5622 ,\u2_Display/n5624 }),
    .b({\u2_Display/n5621 ,\u2_Display/n5623 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add171/c19 ),
    .f({\u2_Display/n5646 [21],\u2_Display/n5646 [19]}),
    .fco(\u2_Display/add171/c23 ),
    .fx({\u2_Display/n5646 [22],\u2_Display/n5646 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u23_al_u4462  (
    .a({\u2_Display/n5618 ,\u2_Display/n5620 }),
    .b({\u2_Display/n5617 ,\u2_Display/n5619 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add171/c23 ),
    .f({\u2_Display/n5646 [25],\u2_Display/n5646 [23]}),
    .fco(\u2_Display/add171/c27 ),
    .fx({\u2_Display/n5646 [26],\u2_Display/n5646 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u27_al_u4463  (
    .a({\u2_Display/n5614 ,\u2_Display/n5616 }),
    .b({\u2_Display/n5613 ,\u2_Display/n5615 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add171/c27 ),
    .f({\u2_Display/n5646 [29],\u2_Display/n5646 [27]}),
    .fco(\u2_Display/add171/c31 ),
    .fx({\u2_Display/n5646 [30],\u2_Display/n5646 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u31_al_u4464  (
    .a({open_n11646,\u2_Display/n5612 }),
    .c(2'b00),
    .d({open_n11651,1'b1}),
    .fci(\u2_Display/add171/c31 ),
    .f({open_n11668,\u2_Display/n5646 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u3_al_u4457  (
    .a({\u2_Display/n5638 ,\u2_Display/n5640 }),
    .b({\u2_Display/n5637 ,\u2_Display/n5639 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add171/c3 ),
    .f({\u2_Display/n5646 [5],\u2_Display/n5646 [3]}),
    .fco(\u2_Display/add171/c7 ),
    .fx({\u2_Display/n5646 [6],\u2_Display/n5646 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/u7_al_u4458  (
    .a({\u2_Display/n5634 ,\u2_Display/n5636 }),
    .b({\u2_Display/n5633 ,\u2_Display/n5635 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add171/c7 ),
    .f({\u2_Display/n5646 [9],\u2_Display/n5646 [7]}),
    .fco(\u2_Display/add171/c11 ),
    .fx({\u2_Display/n5646 [10],\u2_Display/n5646 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add171/ucin_al_u4456"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add171/ucin_al_u4456  (
    .a({\u2_Display/n5642 ,1'b1}),
    .b({\u2_Display/n5641 ,\u2_Display/n5643 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5646 [1],open_n11727}),
    .fco(\u2_Display/add171/c3 ),
    .fx({\u2_Display/n5646 [2],\u2_Display/n5646 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add172/ucin_al_u5049"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add172/u3_al_u5050  (
    .a({\u2_Display/n5673 ,\u2_Display/n5675 }),
    .b({\u2_Display/n5672 ,\u2_Display/n5674 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add172/c3 ),
    .f({\u2_Display/n5681 [5],\u2_Display/n5681 [3]}),
    .fco(\u2_Display/add172/c7 ),
    .fx({\u2_Display/n5681 [6],\u2_Display/n5681 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add172/ucin_al_u5049"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add172/u7_al_u5051  (
    .a({\u2_Display/n5669 ,\u2_Display/n5671 }),
    .b({open_n11748,\u2_Display/n5670 }),
    .c(2'b00),
    .d(2'b00),
    .e({open_n11751,1'b1}),
    .fci(\u2_Display/add172/c7 ),
    .f({\u2_Display/n5681 [9],\u2_Display/n5681 [7]}),
    .fx({open_n11767,\u2_Display/n5681 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add172/ucin_al_u5049"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add172/ucin_al_u5049  (
    .a({\u2_Display/n5677 ,1'b1}),
    .b({\u2_Display/n5676 ,\u2_Display/n5678 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n5681 [1],open_n11787}),
    .fco(\u2_Display/add172/c3 ),
    .fx({\u2_Display/n5681 [2],\u2_Display/n5681 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u11_al_u4468  (
    .a({\u2_Display/counta [13],\u2_Display/counta [11]}),
    .b({\u2_Display/counta [14],\u2_Display/counta [12]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add18/c11 ),
    .f({\u2_Display/n419 [13],\u2_Display/n419 [11]}),
    .fco(\u2_Display/add18/c15 ),
    .fx({\u2_Display/n419 [14],\u2_Display/n419 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u15_al_u4469  (
    .a({\u2_Display/counta [17],\u2_Display/counta [15]}),
    .b({\u2_Display/counta [18],\u2_Display/counta [16]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add18/c15 ),
    .f({\u2_Display/n419 [17],\u2_Display/n419 [15]}),
    .fco(\u2_Display/add18/c19 ),
    .fx({\u2_Display/n419 [18],\u2_Display/n419 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u19_al_u4470  (
    .a({\u2_Display/counta [21],\u2_Display/counta [19]}),
    .b({\u2_Display/counta [22],\u2_Display/counta [20]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add18/c19 ),
    .f({\u2_Display/n419 [21],\u2_Display/n419 [19]}),
    .fco(\u2_Display/add18/c23 ),
    .fx({\u2_Display/n419 [22],\u2_Display/n419 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u23_al_u4471  (
    .a({\u2_Display/counta [25],\u2_Display/counta [23]}),
    .b({\u2_Display/counta [26],\u2_Display/counta [24]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add18/c23 ),
    .f({\u2_Display/n419 [25],\u2_Display/n419 [23]}),
    .fco(\u2_Display/add18/c27 ),
    .fx({\u2_Display/n419 [26],\u2_Display/n419 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u27_al_u4472  (
    .a({\u2_Display/counta [29],\u2_Display/counta [27]}),
    .b({\u2_Display/counta [30],\u2_Display/counta [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add18/c27 ),
    .f({\u2_Display/n419 [29],\u2_Display/n419 [27]}),
    .fco(\u2_Display/add18/c31 ),
    .fx({\u2_Display/n419 [30],\u2_Display/n419 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u31_al_u4473  (
    .a({open_n11880,\u2_Display/counta [31]}),
    .c(2'b00),
    .d({open_n11885,1'b0}),
    .fci(\u2_Display/add18/c31 ),
    .f({open_n11902,\u2_Display/n419 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u3_al_u4466  (
    .a({\u2_Display/counta [5],\u2_Display/counta [3]}),
    .b({\u2_Display/counta [6],\u2_Display/counta [4]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add18/c3 ),
    .f({\u2_Display/n419 [5],\u2_Display/n419 [3]}),
    .fco(\u2_Display/add18/c7 ),
    .fx({\u2_Display/n419 [6],\u2_Display/n419 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/u7_al_u4467  (
    .a({\u2_Display/counta [9],\u2_Display/counta [7]}),
    .b({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add18/c7 ),
    .f({\u2_Display/n419 [9],\u2_Display/n419 [7]}),
    .fco(\u2_Display/add18/c11 ),
    .fx({\u2_Display/n419 [10],\u2_Display/n419 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add18/ucin_al_u4465"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add18/ucin_al_u4465  (
    .a({\u2_Display/counta [1],1'b1}),
    .b({\u2_Display/counta [2],\u2_Display/counta [0]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n419 [1],open_n11961}),
    .fco(\u2_Display/add18/c3 ),
    .fx({\u2_Display/n419 [2],\u2_Display/n419 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u11_al_u4477  (
    .a({\u2_Display/n438 ,\u2_Display/n440 }),
    .b({\u2_Display/n437 ,\u2_Display/n439 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add19/c11 ),
    .f({\u2_Display/n454 [13],\u2_Display/n454 [11]}),
    .fco(\u2_Display/add19/c15 ),
    .fx({\u2_Display/n454 [14],\u2_Display/n454 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u15_al_u4478  (
    .a({\u2_Display/n434 ,\u2_Display/n436 }),
    .b({\u2_Display/n433 ,\u2_Display/n435 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add19/c15 ),
    .f({\u2_Display/n454 [17],\u2_Display/n454 [15]}),
    .fco(\u2_Display/add19/c19 ),
    .fx({\u2_Display/n454 [18],\u2_Display/n454 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u19_al_u4479  (
    .a({\u2_Display/n430 ,\u2_Display/n432 }),
    .b({\u2_Display/n429 ,\u2_Display/n431 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add19/c19 ),
    .f({\u2_Display/n454 [21],\u2_Display/n454 [19]}),
    .fco(\u2_Display/add19/c23 ),
    .fx({\u2_Display/n454 [22],\u2_Display/n454 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u23_al_u4480  (
    .a({\u2_Display/n426 ,\u2_Display/n428 }),
    .b({\u2_Display/n425 ,\u2_Display/n427 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add19/c23 ),
    .f({\u2_Display/n454 [25],\u2_Display/n454 [23]}),
    .fco(\u2_Display/add19/c27 ),
    .fx({\u2_Display/n454 [26],\u2_Display/n454 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u27_al_u4481  (
    .a({\u2_Display/n422 ,\u2_Display/n424 }),
    .b({\u2_Display/n421 ,\u2_Display/n423 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add19/c27 ),
    .f({\u2_Display/n454 [29],\u2_Display/n454 [27]}),
    .fco(\u2_Display/add19/c31 ),
    .fx({\u2_Display/n454 [30],\u2_Display/n454 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u31_al_u4482  (
    .a({open_n12054,\u2_Display/n420 }),
    .c(2'b00),
    .d({open_n12059,1'b1}),
    .fci(\u2_Display/add19/c31 ),
    .f({open_n12076,\u2_Display/n454 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u3_al_u4475  (
    .a({\u2_Display/n446 ,\u2_Display/n448 }),
    .b({\u2_Display/n445 ,\u2_Display/n447 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add19/c3 ),
    .f({\u2_Display/n454 [5],\u2_Display/n454 [3]}),
    .fco(\u2_Display/add19/c7 ),
    .fx({\u2_Display/n454 [6],\u2_Display/n454 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/u7_al_u4476  (
    .a({\u2_Display/n442 ,\u2_Display/n444 }),
    .b({\u2_Display/n441 ,\u2_Display/n443 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add19/c7 ),
    .f({\u2_Display/n454 [9],\u2_Display/n454 [7]}),
    .fco(\u2_Display/add19/c11 ),
    .fx({\u2_Display/n454 [10],\u2_Display/n454 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add19/ucin_al_u4474"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add19/ucin_al_u4474  (
    .a({\u2_Display/n450 ,1'b1}),
    .b({\u2_Display/n449 ,\u2_Display/n451 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n454 [1],open_n12135}),
    .fco(\u2_Display/add19/c3 ),
    .fx({\u2_Display/n454 [2],\u2_Display/n454 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u11_al_u4486  (
    .a({\u2_Display/n473 ,\u2_Display/n475 }),
    .b({\u2_Display/n472 ,\u2_Display/n474 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add20/c11 ),
    .f({\u2_Display/n489 [13],\u2_Display/n489 [11]}),
    .fco(\u2_Display/add20/c15 ),
    .fx({\u2_Display/n489 [14],\u2_Display/n489 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u15_al_u4487  (
    .a({\u2_Display/n469 ,\u2_Display/n471 }),
    .b({\u2_Display/n468 ,\u2_Display/n470 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add20/c15 ),
    .f({\u2_Display/n489 [17],\u2_Display/n489 [15]}),
    .fco(\u2_Display/add20/c19 ),
    .fx({\u2_Display/n489 [18],\u2_Display/n489 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u19_al_u4488  (
    .a({\u2_Display/n465 ,\u2_Display/n467 }),
    .b({\u2_Display/n464 ,\u2_Display/n466 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add20/c19 ),
    .f({\u2_Display/n489 [21],\u2_Display/n489 [19]}),
    .fco(\u2_Display/add20/c23 ),
    .fx({\u2_Display/n489 [22],\u2_Display/n489 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u23_al_u4489  (
    .a({\u2_Display/n461 ,\u2_Display/n463 }),
    .b({\u2_Display/n460 ,\u2_Display/n462 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b01),
    .fci(\u2_Display/add20/c23 ),
    .f({\u2_Display/n489 [25],\u2_Display/n489 [23]}),
    .fco(\u2_Display/add20/c27 ),
    .fx({\u2_Display/n489 [26],\u2_Display/n489 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u27_al_u4490  (
    .a({\u2_Display/n457 ,\u2_Display/n459 }),
    .b({\u2_Display/n456 ,\u2_Display/n458 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add20/c27 ),
    .f({\u2_Display/n489 [29],\u2_Display/n489 [27]}),
    .fco(\u2_Display/add20/c31 ),
    .fx({\u2_Display/n489 [30],\u2_Display/n489 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u31_al_u4491  (
    .a({open_n12228,\u2_Display/n455 }),
    .c(2'b00),
    .d({open_n12233,1'b1}),
    .fci(\u2_Display/add20/c31 ),
    .f({open_n12250,\u2_Display/n489 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u3_al_u4484  (
    .a({\u2_Display/n481 ,\u2_Display/n483 }),
    .b({\u2_Display/n480 ,\u2_Display/n482 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add20/c3 ),
    .f({\u2_Display/n489 [5],\u2_Display/n489 [3]}),
    .fco(\u2_Display/add20/c7 ),
    .fx({\u2_Display/n489 [6],\u2_Display/n489 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/u7_al_u4485  (
    .a({\u2_Display/n477 ,\u2_Display/n479 }),
    .b({\u2_Display/n476 ,\u2_Display/n478 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add20/c7 ),
    .f({\u2_Display/n489 [9],\u2_Display/n489 [7]}),
    .fco(\u2_Display/add20/c11 ),
    .fx({\u2_Display/n489 [10],\u2_Display/n489 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add20/ucin_al_u4483"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add20/ucin_al_u4483  (
    .a({\u2_Display/n485 ,1'b1}),
    .b({\u2_Display/n484 ,\u2_Display/n486 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n489 [1],open_n12309}),
    .fco(\u2_Display/add20/c3 ),
    .fx({\u2_Display/n489 [2],\u2_Display/n489 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u11_al_u4495  (
    .a({\u2_Display/n508 ,\u2_Display/n510 }),
    .b({\u2_Display/n507 ,\u2_Display/n509 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add21/c11 ),
    .f({\u2_Display/n524 [13],\u2_Display/n524 [11]}),
    .fco(\u2_Display/add21/c15 ),
    .fx({\u2_Display/n524 [14],\u2_Display/n524 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u15_al_u4496  (
    .a({\u2_Display/n504 ,\u2_Display/n506 }),
    .b({\u2_Display/n503 ,\u2_Display/n505 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add21/c15 ),
    .f({\u2_Display/n524 [17],\u2_Display/n524 [15]}),
    .fco(\u2_Display/add21/c19 ),
    .fx({\u2_Display/n524 [18],\u2_Display/n524 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u19_al_u4497  (
    .a({\u2_Display/n500 ,\u2_Display/n502 }),
    .b({\u2_Display/n499 ,\u2_Display/n501 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add21/c19 ),
    .f({\u2_Display/n524 [21],\u2_Display/n524 [19]}),
    .fco(\u2_Display/add21/c23 ),
    .fx({\u2_Display/n524 [22],\u2_Display/n524 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u23_al_u4498  (
    .a({\u2_Display/n496 ,\u2_Display/n498 }),
    .b({\u2_Display/n495 ,\u2_Display/n497 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add21/c23 ),
    .f({\u2_Display/n524 [25],\u2_Display/n524 [23]}),
    .fco(\u2_Display/add21/c27 ),
    .fx({\u2_Display/n524 [26],\u2_Display/n524 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u27_al_u4499  (
    .a({\u2_Display/n492 ,\u2_Display/n494 }),
    .b({\u2_Display/n491 ,\u2_Display/n493 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add21/c27 ),
    .f({\u2_Display/n524 [29],\u2_Display/n524 [27]}),
    .fco(\u2_Display/add21/c31 ),
    .fx({\u2_Display/n524 [30],\u2_Display/n524 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u31_al_u4500  (
    .a({open_n12402,\u2_Display/n490 }),
    .c(2'b00),
    .d({open_n12407,1'b1}),
    .fci(\u2_Display/add21/c31 ),
    .f({open_n12424,\u2_Display/n524 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u3_al_u4493  (
    .a({\u2_Display/n516 ,\u2_Display/n518 }),
    .b({\u2_Display/n515 ,\u2_Display/n517 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add21/c3 ),
    .f({\u2_Display/n524 [5],\u2_Display/n524 [3]}),
    .fco(\u2_Display/add21/c7 ),
    .fx({\u2_Display/n524 [6],\u2_Display/n524 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/u7_al_u4494  (
    .a({\u2_Display/n512 ,\u2_Display/n514 }),
    .b({\u2_Display/n511 ,\u2_Display/n513 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add21/c7 ),
    .f({\u2_Display/n524 [9],\u2_Display/n524 [7]}),
    .fco(\u2_Display/add21/c11 ),
    .fx({\u2_Display/n524 [10],\u2_Display/n524 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add21/ucin_al_u4492"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add21/ucin_al_u4492  (
    .a({\u2_Display/n520 ,1'b1}),
    .b({\u2_Display/n519 ,\u2_Display/n521 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n524 [1],open_n12483}),
    .fco(\u2_Display/add21/c3 ),
    .fx({\u2_Display/n524 [2],\u2_Display/n524 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u11_al_u4504  (
    .a({\u2_Display/n543 ,\u2_Display/n545 }),
    .b({\u2_Display/n542 ,\u2_Display/n544 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add22/c11 ),
    .f({\u2_Display/n559 [13],\u2_Display/n559 [11]}),
    .fco(\u2_Display/add22/c15 ),
    .fx({\u2_Display/n559 [14],\u2_Display/n559 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u15_al_u4505  (
    .a({\u2_Display/n539 ,\u2_Display/n541 }),
    .b({\u2_Display/n538 ,\u2_Display/n540 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add22/c15 ),
    .f({\u2_Display/n559 [17],\u2_Display/n559 [15]}),
    .fco(\u2_Display/add22/c19 ),
    .fx({\u2_Display/n559 [18],\u2_Display/n559 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u19_al_u4506  (
    .a({\u2_Display/n535 ,\u2_Display/n537 }),
    .b({\u2_Display/n534 ,\u2_Display/n536 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add22/c19 ),
    .f({\u2_Display/n559 [21],\u2_Display/n559 [19]}),
    .fco(\u2_Display/add22/c23 ),
    .fx({\u2_Display/n559 [22],\u2_Display/n559 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u23_al_u4507  (
    .a({\u2_Display/n531 ,\u2_Display/n533 }),
    .b({\u2_Display/n530 ,\u2_Display/n532 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add22/c23 ),
    .f({\u2_Display/n559 [25],\u2_Display/n559 [23]}),
    .fco(\u2_Display/add22/c27 ),
    .fx({\u2_Display/n559 [26],\u2_Display/n559 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u27_al_u4508  (
    .a({\u2_Display/n527 ,\u2_Display/n529 }),
    .b({\u2_Display/n526 ,\u2_Display/n528 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add22/c27 ),
    .f({\u2_Display/n559 [29],\u2_Display/n559 [27]}),
    .fco(\u2_Display/add22/c31 ),
    .fx({\u2_Display/n559 [30],\u2_Display/n559 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u31_al_u4509  (
    .a({open_n12576,\u2_Display/n525 }),
    .c(2'b00),
    .d({open_n12581,1'b1}),
    .fci(\u2_Display/add22/c31 ),
    .f({open_n12598,\u2_Display/n559 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u3_al_u4502  (
    .a({\u2_Display/n551 ,\u2_Display/n553 }),
    .b({\u2_Display/n550 ,\u2_Display/n552 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add22/c3 ),
    .f({\u2_Display/n559 [5],\u2_Display/n559 [3]}),
    .fco(\u2_Display/add22/c7 ),
    .fx({\u2_Display/n559 [6],\u2_Display/n559 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/u7_al_u4503  (
    .a({\u2_Display/n547 ,\u2_Display/n549 }),
    .b({\u2_Display/n546 ,\u2_Display/n548 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add22/c7 ),
    .f({\u2_Display/n559 [9],\u2_Display/n559 [7]}),
    .fco(\u2_Display/add22/c11 ),
    .fx({\u2_Display/n559 [10],\u2_Display/n559 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add22/ucin_al_u4501"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add22/ucin_al_u4501  (
    .a({\u2_Display/n555 ,1'b1}),
    .b({\u2_Display/n554 ,\u2_Display/n556 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n559 [1],open_n12657}),
    .fco(\u2_Display/add22/c3 ),
    .fx({\u2_Display/n559 [2],\u2_Display/n559 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u11_al_u4513  (
    .a({\u2_Display/n578 ,\u2_Display/n580 }),
    .b({\u2_Display/n577 ,\u2_Display/n579 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add23/c11 ),
    .f({\u2_Display/n594 [13],\u2_Display/n594 [11]}),
    .fco(\u2_Display/add23/c15 ),
    .fx({\u2_Display/n594 [14],\u2_Display/n594 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u15_al_u4514  (
    .a({\u2_Display/n574 ,\u2_Display/n576 }),
    .b({\u2_Display/n573 ,\u2_Display/n575 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add23/c15 ),
    .f({\u2_Display/n594 [17],\u2_Display/n594 [15]}),
    .fco(\u2_Display/add23/c19 ),
    .fx({\u2_Display/n594 [18],\u2_Display/n594 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u19_al_u4515  (
    .a({\u2_Display/n570 ,\u2_Display/n572 }),
    .b({\u2_Display/n569 ,\u2_Display/n571 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add23/c19 ),
    .f({\u2_Display/n594 [21],\u2_Display/n594 [19]}),
    .fco(\u2_Display/add23/c23 ),
    .fx({\u2_Display/n594 [22],\u2_Display/n594 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u23_al_u4516  (
    .a({\u2_Display/n566 ,\u2_Display/n568 }),
    .b({\u2_Display/n565 ,\u2_Display/n567 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add23/c23 ),
    .f({\u2_Display/n594 [25],\u2_Display/n594 [23]}),
    .fco(\u2_Display/add23/c27 ),
    .fx({\u2_Display/n594 [26],\u2_Display/n594 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u27_al_u4517  (
    .a({\u2_Display/n562 ,\u2_Display/n564 }),
    .b({\u2_Display/n561 ,\u2_Display/n563 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add23/c27 ),
    .f({\u2_Display/n594 [29],\u2_Display/n594 [27]}),
    .fco(\u2_Display/add23/c31 ),
    .fx({\u2_Display/n594 [30],\u2_Display/n594 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u31_al_u4518  (
    .a({open_n12750,\u2_Display/n560 }),
    .c(2'b00),
    .d({open_n12755,1'b1}),
    .fci(\u2_Display/add23/c31 ),
    .f({open_n12772,\u2_Display/n594 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u3_al_u4511  (
    .a({\u2_Display/n586 ,\u2_Display/n588 }),
    .b({\u2_Display/n585 ,\u2_Display/n587 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add23/c3 ),
    .f({\u2_Display/n594 [5],\u2_Display/n594 [3]}),
    .fco(\u2_Display/add23/c7 ),
    .fx({\u2_Display/n594 [6],\u2_Display/n594 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/u7_al_u4512  (
    .a({\u2_Display/n582 ,\u2_Display/n584 }),
    .b({\u2_Display/n581 ,\u2_Display/n583 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add23/c7 ),
    .f({\u2_Display/n594 [9],\u2_Display/n594 [7]}),
    .fco(\u2_Display/add23/c11 ),
    .fx({\u2_Display/n594 [10],\u2_Display/n594 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add23/ucin_al_u4510"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add23/ucin_al_u4510  (
    .a({\u2_Display/n590 ,1'b1}),
    .b({\u2_Display/n589 ,\u2_Display/n591 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n594 [1],open_n12831}),
    .fco(\u2_Display/add23/c3 ),
    .fx({\u2_Display/n594 [2],\u2_Display/n594 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u11_al_u4522  (
    .a({\u2_Display/n613 ,\u2_Display/n615 }),
    .b({\u2_Display/n612 ,\u2_Display/n614 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add24/c11 ),
    .f({\u2_Display/n629 [13],\u2_Display/n629 [11]}),
    .fco(\u2_Display/add24/c15 ),
    .fx({\u2_Display/n629 [14],\u2_Display/n629 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u15_al_u4523  (
    .a({\u2_Display/n609 ,\u2_Display/n611 }),
    .b({\u2_Display/n608 ,\u2_Display/n610 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add24/c15 ),
    .f({\u2_Display/n629 [17],\u2_Display/n629 [15]}),
    .fco(\u2_Display/add24/c19 ),
    .fx({\u2_Display/n629 [18],\u2_Display/n629 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u19_al_u4524  (
    .a({\u2_Display/n605 ,\u2_Display/n607 }),
    .b({\u2_Display/n604 ,\u2_Display/n606 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b01),
    .fci(\u2_Display/add24/c19 ),
    .f({\u2_Display/n629 [21],\u2_Display/n629 [19]}),
    .fco(\u2_Display/add24/c23 ),
    .fx({\u2_Display/n629 [22],\u2_Display/n629 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u23_al_u4525  (
    .a({\u2_Display/n601 ,\u2_Display/n603 }),
    .b({\u2_Display/n600 ,\u2_Display/n602 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add24/c23 ),
    .f({\u2_Display/n629 [25],\u2_Display/n629 [23]}),
    .fco(\u2_Display/add24/c27 ),
    .fx({\u2_Display/n629 [26],\u2_Display/n629 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u27_al_u4526  (
    .a({\u2_Display/n597 ,\u2_Display/n599 }),
    .b({\u2_Display/n596 ,\u2_Display/n598 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add24/c27 ),
    .f({\u2_Display/n629 [29],\u2_Display/n629 [27]}),
    .fco(\u2_Display/add24/c31 ),
    .fx({\u2_Display/n629 [30],\u2_Display/n629 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u31_al_u4527  (
    .a({open_n12924,\u2_Display/n595 }),
    .c(2'b00),
    .d({open_n12929,1'b1}),
    .fci(\u2_Display/add24/c31 ),
    .f({open_n12946,\u2_Display/n629 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u3_al_u4520  (
    .a({\u2_Display/n621 ,\u2_Display/n623 }),
    .b({\u2_Display/n620 ,\u2_Display/n622 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add24/c3 ),
    .f({\u2_Display/n629 [5],\u2_Display/n629 [3]}),
    .fco(\u2_Display/add24/c7 ),
    .fx({\u2_Display/n629 [6],\u2_Display/n629 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/u7_al_u4521  (
    .a({\u2_Display/n617 ,\u2_Display/n619 }),
    .b({\u2_Display/n616 ,\u2_Display/n618 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add24/c7 ),
    .f({\u2_Display/n629 [9],\u2_Display/n629 [7]}),
    .fco(\u2_Display/add24/c11 ),
    .fx({\u2_Display/n629 [10],\u2_Display/n629 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add24/ucin_al_u4519"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add24/ucin_al_u4519  (
    .a({\u2_Display/n625 ,1'b1}),
    .b({\u2_Display/n624 ,\u2_Display/n626 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n629 [1],open_n13005}),
    .fco(\u2_Display/add24/c3 ),
    .fx({\u2_Display/n629 [2],\u2_Display/n629 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u11_al_u4531  (
    .a({\u2_Display/n648 ,\u2_Display/n650 }),
    .b({\u2_Display/n647 ,\u2_Display/n649 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add25/c11 ),
    .f({\u2_Display/n664 [13],\u2_Display/n664 [11]}),
    .fco(\u2_Display/add25/c15 ),
    .fx({\u2_Display/n664 [14],\u2_Display/n664 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u15_al_u4532  (
    .a({\u2_Display/n644 ,\u2_Display/n646 }),
    .b({\u2_Display/n643 ,\u2_Display/n645 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add25/c15 ),
    .f({\u2_Display/n664 [17],\u2_Display/n664 [15]}),
    .fco(\u2_Display/add25/c19 ),
    .fx({\u2_Display/n664 [18],\u2_Display/n664 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u19_al_u4533  (
    .a({\u2_Display/n640 ,\u2_Display/n642 }),
    .b({\u2_Display/n639 ,\u2_Display/n641 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add25/c19 ),
    .f({\u2_Display/n664 [21],\u2_Display/n664 [19]}),
    .fco(\u2_Display/add25/c23 ),
    .fx({\u2_Display/n664 [22],\u2_Display/n664 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u23_al_u4534  (
    .a({\u2_Display/n636 ,\u2_Display/n638 }),
    .b({\u2_Display/n635 ,\u2_Display/n637 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add25/c23 ),
    .f({\u2_Display/n664 [25],\u2_Display/n664 [23]}),
    .fco(\u2_Display/add25/c27 ),
    .fx({\u2_Display/n664 [26],\u2_Display/n664 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u27_al_u4535  (
    .a({\u2_Display/n632 ,\u2_Display/n634 }),
    .b({\u2_Display/n631 ,\u2_Display/n633 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add25/c27 ),
    .f({\u2_Display/n664 [29],\u2_Display/n664 [27]}),
    .fco(\u2_Display/add25/c31 ),
    .fx({\u2_Display/n664 [30],\u2_Display/n664 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u31_al_u4536  (
    .a({open_n13098,\u2_Display/n630 }),
    .c(2'b00),
    .d({open_n13103,1'b1}),
    .fci(\u2_Display/add25/c31 ),
    .f({open_n13120,\u2_Display/n664 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u3_al_u4529  (
    .a({\u2_Display/n656 ,\u2_Display/n658 }),
    .b({\u2_Display/n655 ,\u2_Display/n657 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add25/c3 ),
    .f({\u2_Display/n664 [5],\u2_Display/n664 [3]}),
    .fco(\u2_Display/add25/c7 ),
    .fx({\u2_Display/n664 [6],\u2_Display/n664 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/u7_al_u4530  (
    .a({\u2_Display/n652 ,\u2_Display/n654 }),
    .b({\u2_Display/n651 ,\u2_Display/n653 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add25/c7 ),
    .f({\u2_Display/n664 [9],\u2_Display/n664 [7]}),
    .fco(\u2_Display/add25/c11 ),
    .fx({\u2_Display/n664 [10],\u2_Display/n664 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add25/ucin_al_u4528"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add25/ucin_al_u4528  (
    .a({\u2_Display/n660 ,1'b1}),
    .b({\u2_Display/n659 ,\u2_Display/n661 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n664 [1],open_n13179}),
    .fco(\u2_Display/add25/c3 ),
    .fx({\u2_Display/n664 [2],\u2_Display/n664 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u11_al_u4540  (
    .a({\u2_Display/n683 ,\u2_Display/n685 }),
    .b({\u2_Display/n682 ,\u2_Display/n684 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add26/c11 ),
    .f({\u2_Display/n699 [13],\u2_Display/n699 [11]}),
    .fco(\u2_Display/add26/c15 ),
    .fx({\u2_Display/n699 [14],\u2_Display/n699 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u15_al_u4541  (
    .a({\u2_Display/n679 ,\u2_Display/n681 }),
    .b({\u2_Display/n678 ,\u2_Display/n680 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add26/c15 ),
    .f({\u2_Display/n699 [17],\u2_Display/n699 [15]}),
    .fco(\u2_Display/add26/c19 ),
    .fx({\u2_Display/n699 [18],\u2_Display/n699 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u19_al_u4542  (
    .a({\u2_Display/n675 ,\u2_Display/n677 }),
    .b({\u2_Display/n674 ,\u2_Display/n676 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add26/c19 ),
    .f({\u2_Display/n699 [21],\u2_Display/n699 [19]}),
    .fco(\u2_Display/add26/c23 ),
    .fx({\u2_Display/n699 [22],\u2_Display/n699 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u23_al_u4543  (
    .a({\u2_Display/n671 ,\u2_Display/n673 }),
    .b({\u2_Display/n670 ,\u2_Display/n672 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add26/c23 ),
    .f({\u2_Display/n699 [25],\u2_Display/n699 [23]}),
    .fco(\u2_Display/add26/c27 ),
    .fx({\u2_Display/n699 [26],\u2_Display/n699 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u27_al_u4544  (
    .a({\u2_Display/n667 ,\u2_Display/n669 }),
    .b({\u2_Display/n666 ,\u2_Display/n668 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add26/c27 ),
    .f({\u2_Display/n699 [29],\u2_Display/n699 [27]}),
    .fco(\u2_Display/add26/c31 ),
    .fx({\u2_Display/n699 [30],\u2_Display/n699 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u31_al_u4545  (
    .a({open_n13272,\u2_Display/n665 }),
    .c(2'b00),
    .d({open_n13277,1'b1}),
    .fci(\u2_Display/add26/c31 ),
    .f({open_n13294,\u2_Display/n699 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u3_al_u4538  (
    .a({\u2_Display/n691 ,\u2_Display/n693 }),
    .b({\u2_Display/n690 ,\u2_Display/n692 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add26/c3 ),
    .f({\u2_Display/n699 [5],\u2_Display/n699 [3]}),
    .fco(\u2_Display/add26/c7 ),
    .fx({\u2_Display/n699 [6],\u2_Display/n699 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/u7_al_u4539  (
    .a({\u2_Display/n687 ,\u2_Display/n689 }),
    .b({\u2_Display/n686 ,\u2_Display/n688 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add26/c7 ),
    .f({\u2_Display/n699 [9],\u2_Display/n699 [7]}),
    .fco(\u2_Display/add26/c11 ),
    .fx({\u2_Display/n699 [10],\u2_Display/n699 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add26/ucin_al_u4537"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add26/ucin_al_u4537  (
    .a({\u2_Display/n695 ,1'b1}),
    .b({\u2_Display/n694 ,\u2_Display/n696 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n699 [1],open_n13353}),
    .fco(\u2_Display/add26/c3 ),
    .fx({\u2_Display/n699 [2],\u2_Display/n699 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u11_al_u4549  (
    .a({\u2_Display/n718 ,\u2_Display/n720 }),
    .b({\u2_Display/n717 ,\u2_Display/n719 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add27/c11 ),
    .f({\u2_Display/n734 [13],\u2_Display/n734 [11]}),
    .fco(\u2_Display/add27/c15 ),
    .fx({\u2_Display/n734 [14],\u2_Display/n734 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u15_al_u4550  (
    .a({\u2_Display/n714 ,\u2_Display/n716 }),
    .b({\u2_Display/n713 ,\u2_Display/n715 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add27/c15 ),
    .f({\u2_Display/n734 [17],\u2_Display/n734 [15]}),
    .fco(\u2_Display/add27/c19 ),
    .fx({\u2_Display/n734 [18],\u2_Display/n734 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u19_al_u4551  (
    .a({\u2_Display/n710 ,\u2_Display/n712 }),
    .b({\u2_Display/n709 ,\u2_Display/n711 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add27/c19 ),
    .f({\u2_Display/n734 [21],\u2_Display/n734 [19]}),
    .fco(\u2_Display/add27/c23 ),
    .fx({\u2_Display/n734 [22],\u2_Display/n734 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u23_al_u4552  (
    .a({\u2_Display/n706 ,\u2_Display/n708 }),
    .b({\u2_Display/n705 ,\u2_Display/n707 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add27/c23 ),
    .f({\u2_Display/n734 [25],\u2_Display/n734 [23]}),
    .fco(\u2_Display/add27/c27 ),
    .fx({\u2_Display/n734 [26],\u2_Display/n734 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u27_al_u4553  (
    .a({\u2_Display/n702 ,\u2_Display/n704 }),
    .b({\u2_Display/n701 ,\u2_Display/n703 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add27/c27 ),
    .f({\u2_Display/n734 [29],\u2_Display/n734 [27]}),
    .fco(\u2_Display/add27/c31 ),
    .fx({\u2_Display/n734 [30],\u2_Display/n734 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u31_al_u4554  (
    .a({open_n13446,\u2_Display/n700 }),
    .c(2'b00),
    .d({open_n13451,1'b1}),
    .fci(\u2_Display/add27/c31 ),
    .f({open_n13468,\u2_Display/n734 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u3_al_u4547  (
    .a({\u2_Display/n726 ,\u2_Display/n728 }),
    .b({\u2_Display/n725 ,\u2_Display/n727 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add27/c3 ),
    .f({\u2_Display/n734 [5],\u2_Display/n734 [3]}),
    .fco(\u2_Display/add27/c7 ),
    .fx({\u2_Display/n734 [6],\u2_Display/n734 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/u7_al_u4548  (
    .a({\u2_Display/n722 ,\u2_Display/n724 }),
    .b({\u2_Display/n721 ,\u2_Display/n723 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add27/c7 ),
    .f({\u2_Display/n734 [9],\u2_Display/n734 [7]}),
    .fco(\u2_Display/add27/c11 ),
    .fx({\u2_Display/n734 [10],\u2_Display/n734 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add27/ucin_al_u4546"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add27/ucin_al_u4546  (
    .a({\u2_Display/n730 ,1'b1}),
    .b({\u2_Display/n729 ,\u2_Display/n731 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n734 [1],open_n13527}),
    .fco(\u2_Display/add27/c3 ),
    .fx({\u2_Display/n734 [2],\u2_Display/n734 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u11_al_u4558  (
    .a({\u2_Display/n753 ,\u2_Display/n755 }),
    .b({\u2_Display/n752 ,\u2_Display/n754 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add28/c11 ),
    .f({\u2_Display/n769 [13],\u2_Display/n769 [11]}),
    .fco(\u2_Display/add28/c15 ),
    .fx({\u2_Display/n769 [14],\u2_Display/n769 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u15_al_u4559  (
    .a({\u2_Display/n749 ,\u2_Display/n751 }),
    .b({\u2_Display/n748 ,\u2_Display/n750 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b01),
    .fci(\u2_Display/add28/c15 ),
    .f({\u2_Display/n769 [17],\u2_Display/n769 [15]}),
    .fco(\u2_Display/add28/c19 ),
    .fx({\u2_Display/n769 [18],\u2_Display/n769 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u19_al_u4560  (
    .a({\u2_Display/n745 ,\u2_Display/n747 }),
    .b({\u2_Display/n744 ,\u2_Display/n746 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add28/c19 ),
    .f({\u2_Display/n769 [21],\u2_Display/n769 [19]}),
    .fco(\u2_Display/add28/c23 ),
    .fx({\u2_Display/n769 [22],\u2_Display/n769 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u23_al_u4561  (
    .a({\u2_Display/n741 ,\u2_Display/n743 }),
    .b({\u2_Display/n740 ,\u2_Display/n742 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add28/c23 ),
    .f({\u2_Display/n769 [25],\u2_Display/n769 [23]}),
    .fco(\u2_Display/add28/c27 ),
    .fx({\u2_Display/n769 [26],\u2_Display/n769 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u27_al_u4562  (
    .a({\u2_Display/n737 ,\u2_Display/n739 }),
    .b({\u2_Display/n736 ,\u2_Display/n738 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add28/c27 ),
    .f({\u2_Display/n769 [29],\u2_Display/n769 [27]}),
    .fco(\u2_Display/add28/c31 ),
    .fx({\u2_Display/n769 [30],\u2_Display/n769 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u31_al_u4563  (
    .a({open_n13620,\u2_Display/n735 }),
    .c(2'b00),
    .d({open_n13625,1'b1}),
    .fci(\u2_Display/add28/c31 ),
    .f({open_n13642,\u2_Display/n769 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u3_al_u4556  (
    .a({\u2_Display/n761 ,\u2_Display/n763 }),
    .b({\u2_Display/n760 ,\u2_Display/n762 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add28/c3 ),
    .f({\u2_Display/n769 [5],\u2_Display/n769 [3]}),
    .fco(\u2_Display/add28/c7 ),
    .fx({\u2_Display/n769 [6],\u2_Display/n769 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/u7_al_u4557  (
    .a({\u2_Display/n757 ,\u2_Display/n759 }),
    .b({\u2_Display/n756 ,\u2_Display/n758 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add28/c7 ),
    .f({\u2_Display/n769 [9],\u2_Display/n769 [7]}),
    .fco(\u2_Display/add28/c11 ),
    .fx({\u2_Display/n769 [10],\u2_Display/n769 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add28/ucin_al_u4555"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add28/ucin_al_u4555  (
    .a({\u2_Display/n765 ,1'b1}),
    .b({\u2_Display/n764 ,\u2_Display/n766 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n769 [1],open_n13701}),
    .fco(\u2_Display/add28/c3 ),
    .fx({\u2_Display/n769 [2],\u2_Display/n769 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u11_al_u4567  (
    .a({\u2_Display/n788 ,\u2_Display/n790 }),
    .b({\u2_Display/n787 ,\u2_Display/n789 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add29/c11 ),
    .f({\u2_Display/n804 [13],\u2_Display/n804 [11]}),
    .fco(\u2_Display/add29/c15 ),
    .fx({\u2_Display/n804 [14],\u2_Display/n804 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u15_al_u4568  (
    .a({\u2_Display/n784 ,\u2_Display/n786 }),
    .b({\u2_Display/n783 ,\u2_Display/n785 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add29/c15 ),
    .f({\u2_Display/n804 [17],\u2_Display/n804 [15]}),
    .fco(\u2_Display/add29/c19 ),
    .fx({\u2_Display/n804 [18],\u2_Display/n804 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u19_al_u4569  (
    .a({\u2_Display/n780 ,\u2_Display/n782 }),
    .b({\u2_Display/n779 ,\u2_Display/n781 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add29/c19 ),
    .f({\u2_Display/n804 [21],\u2_Display/n804 [19]}),
    .fco(\u2_Display/add29/c23 ),
    .fx({\u2_Display/n804 [22],\u2_Display/n804 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u23_al_u4570  (
    .a({\u2_Display/n776 ,\u2_Display/n778 }),
    .b({\u2_Display/n775 ,\u2_Display/n777 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add29/c23 ),
    .f({\u2_Display/n804 [25],\u2_Display/n804 [23]}),
    .fco(\u2_Display/add29/c27 ),
    .fx({\u2_Display/n804 [26],\u2_Display/n804 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u27_al_u4571  (
    .a({\u2_Display/n772 ,\u2_Display/n774 }),
    .b({\u2_Display/n771 ,\u2_Display/n773 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add29/c27 ),
    .f({\u2_Display/n804 [29],\u2_Display/n804 [27]}),
    .fco(\u2_Display/add29/c31 ),
    .fx({\u2_Display/n804 [30],\u2_Display/n804 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u31_al_u4572  (
    .a({open_n13794,\u2_Display/n770 }),
    .c(2'b00),
    .d({open_n13799,1'b1}),
    .fci(\u2_Display/add29/c31 ),
    .f({open_n13816,\u2_Display/n804 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u3_al_u4565  (
    .a({\u2_Display/n796 ,\u2_Display/n798 }),
    .b({\u2_Display/n795 ,\u2_Display/n797 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add29/c3 ),
    .f({\u2_Display/n804 [5],\u2_Display/n804 [3]}),
    .fco(\u2_Display/add29/c7 ),
    .fx({\u2_Display/n804 [6],\u2_Display/n804 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/u7_al_u4566  (
    .a({\u2_Display/n792 ,\u2_Display/n794 }),
    .b({\u2_Display/n791 ,\u2_Display/n793 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add29/c7 ),
    .f({\u2_Display/n804 [9],\u2_Display/n804 [7]}),
    .fco(\u2_Display/add29/c11 ),
    .fx({\u2_Display/n804 [10],\u2_Display/n804 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add29/ucin_al_u4564"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add29/ucin_al_u4564  (
    .a({\u2_Display/n800 ,1'b1}),
    .b({\u2_Display/n799 ,\u2_Display/n801 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n804 [1],open_n13875}),
    .fco(\u2_Display/add29/c3 ),
    .fx({\u2_Display/n804 [2],\u2_Display/n804 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add2_2/u0|u2_Display/add2_2/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add2_2/u0|u2_Display/add2_2/ucin  (
    .a(2'b10),
    .b({\u2_Display/i [8],open_n13878}),
    .f({\u2_Display/n43 [0],open_n13898}),
    .fco(\u2_Display/add2_2/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add2_2/u0|u2_Display/add2_2/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add2_2/u2|u2_Display/add2_2/u1  (
    .a(2'b10),
    .b(\u2_Display/i [10:9]),
    .fci(\u2_Display/add2_2/c1 ),
    .f(\u2_Display/n43 [2:1]),
    .fco(\u2_Display/add2_2/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add2_2/u0|u2_Display/add2_2/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add2_2/ucout_al_u5058  (
    .fci(\u2_Display/add2_2/c3 ),
    .f({open_n13947,\u2_Display/add2_2_co }));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u11_al_u4576  (
    .a({\u2_Display/n823 ,\u2_Display/n825 }),
    .b({\u2_Display/n822 ,\u2_Display/n824 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add30/c11 ),
    .f({\u2_Display/n839 [13],\u2_Display/n839 [11]}),
    .fco(\u2_Display/add30/c15 ),
    .fx({\u2_Display/n839 [14],\u2_Display/n839 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u15_al_u4577  (
    .a({\u2_Display/n819 ,\u2_Display/n821 }),
    .b({\u2_Display/n818 ,\u2_Display/n820 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add30/c15 ),
    .f({\u2_Display/n839 [17],\u2_Display/n839 [15]}),
    .fco(\u2_Display/add30/c19 ),
    .fx({\u2_Display/n839 [18],\u2_Display/n839 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u19_al_u4578  (
    .a({\u2_Display/n815 ,\u2_Display/n817 }),
    .b({\u2_Display/n814 ,\u2_Display/n816 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add30/c19 ),
    .f({\u2_Display/n839 [21],\u2_Display/n839 [19]}),
    .fco(\u2_Display/add30/c23 ),
    .fx({\u2_Display/n839 [22],\u2_Display/n839 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u23_al_u4579  (
    .a({\u2_Display/n811 ,\u2_Display/n813 }),
    .b({\u2_Display/n810 ,\u2_Display/n812 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add30/c23 ),
    .f({\u2_Display/n839 [25],\u2_Display/n839 [23]}),
    .fco(\u2_Display/add30/c27 ),
    .fx({\u2_Display/n839 [26],\u2_Display/n839 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u27_al_u4580  (
    .a({\u2_Display/n807 ,\u2_Display/n809 }),
    .b({\u2_Display/n806 ,\u2_Display/n808 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add30/c27 ),
    .f({\u2_Display/n839 [29],\u2_Display/n839 [27]}),
    .fco(\u2_Display/add30/c31 ),
    .fx({\u2_Display/n839 [30],\u2_Display/n839 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u31_al_u4581  (
    .a({open_n14043,\u2_Display/n805 }),
    .c(2'b00),
    .d({open_n14048,1'b1}),
    .fci(\u2_Display/add30/c31 ),
    .f({open_n14065,\u2_Display/n839 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u3_al_u4574  (
    .a({\u2_Display/n831 ,\u2_Display/n833 }),
    .b({\u2_Display/n830 ,\u2_Display/n832 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add30/c3 ),
    .f({\u2_Display/n839 [5],\u2_Display/n839 [3]}),
    .fco(\u2_Display/add30/c7 ),
    .fx({\u2_Display/n839 [6],\u2_Display/n839 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/u7_al_u4575  (
    .a({\u2_Display/n827 ,\u2_Display/n829 }),
    .b({\u2_Display/n826 ,\u2_Display/n828 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add30/c7 ),
    .f({\u2_Display/n839 [9],\u2_Display/n839 [7]}),
    .fco(\u2_Display/add30/c11 ),
    .fx({\u2_Display/n839 [10],\u2_Display/n839 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add30/ucin_al_u4573"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add30/ucin_al_u4573  (
    .a({\u2_Display/n835 ,1'b1}),
    .b({\u2_Display/n834 ,\u2_Display/n836 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n839 [1],open_n14124}),
    .fco(\u2_Display/add30/c3 ),
    .fx({\u2_Display/n839 [2],\u2_Display/n839 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u11_al_u4585  (
    .a({\u2_Display/n858 ,\u2_Display/n860 }),
    .b({\u2_Display/n857 ,\u2_Display/n859 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add31/c11 ),
    .f({\u2_Display/n874 [13],\u2_Display/n874 [11]}),
    .fco(\u2_Display/add31/c15 ),
    .fx({\u2_Display/n874 [14],\u2_Display/n874 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u15_al_u4586  (
    .a({\u2_Display/n854 ,\u2_Display/n856 }),
    .b({\u2_Display/n853 ,\u2_Display/n855 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add31/c15 ),
    .f({\u2_Display/n874 [17],\u2_Display/n874 [15]}),
    .fco(\u2_Display/add31/c19 ),
    .fx({\u2_Display/n874 [18],\u2_Display/n874 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u19_al_u4587  (
    .a({\u2_Display/n850 ,\u2_Display/n852 }),
    .b({\u2_Display/n849 ,\u2_Display/n851 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add31/c19 ),
    .f({\u2_Display/n874 [21],\u2_Display/n874 [19]}),
    .fco(\u2_Display/add31/c23 ),
    .fx({\u2_Display/n874 [22],\u2_Display/n874 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u23_al_u4588  (
    .a({\u2_Display/n846 ,\u2_Display/n848 }),
    .b({\u2_Display/n845 ,\u2_Display/n847 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add31/c23 ),
    .f({\u2_Display/n874 [25],\u2_Display/n874 [23]}),
    .fco(\u2_Display/add31/c27 ),
    .fx({\u2_Display/n874 [26],\u2_Display/n874 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u27_al_u4589  (
    .a({\u2_Display/n842 ,\u2_Display/n844 }),
    .b({\u2_Display/n841 ,\u2_Display/n843 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add31/c27 ),
    .f({\u2_Display/n874 [29],\u2_Display/n874 [27]}),
    .fco(\u2_Display/add31/c31 ),
    .fx({\u2_Display/n874 [30],\u2_Display/n874 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u31_al_u4590  (
    .a({open_n14217,\u2_Display/n840 }),
    .c(2'b00),
    .d({open_n14222,1'b1}),
    .fci(\u2_Display/add31/c31 ),
    .f({open_n14239,\u2_Display/n874 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u3_al_u4583  (
    .a({\u2_Display/n866 ,\u2_Display/n868 }),
    .b({\u2_Display/n865 ,\u2_Display/n867 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add31/c3 ),
    .f({\u2_Display/n874 [5],\u2_Display/n874 [3]}),
    .fco(\u2_Display/add31/c7 ),
    .fx({\u2_Display/n874 [6],\u2_Display/n874 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/u7_al_u4584  (
    .a({\u2_Display/n862 ,\u2_Display/n864 }),
    .b({\u2_Display/n861 ,\u2_Display/n863 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add31/c7 ),
    .f({\u2_Display/n874 [9],\u2_Display/n874 [7]}),
    .fco(\u2_Display/add31/c11 ),
    .fx({\u2_Display/n874 [10],\u2_Display/n874 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add31/ucin_al_u4582"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add31/ucin_al_u4582  (
    .a({\u2_Display/n870 ,1'b1}),
    .b({\u2_Display/n869 ,\u2_Display/n871 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n874 [1],open_n14298}),
    .fco(\u2_Display/add31/c3 ),
    .fx({\u2_Display/n874 [2],\u2_Display/n874 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u11_al_u4594  (
    .a({\u2_Display/n893 ,\u2_Display/n895 }),
    .b({\u2_Display/n892 ,\u2_Display/n894 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b01),
    .fci(\u2_Display/add32/c11 ),
    .f({\u2_Display/n909 [13],\u2_Display/n909 [11]}),
    .fco(\u2_Display/add32/c15 ),
    .fx({\u2_Display/n909 [14],\u2_Display/n909 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u15_al_u4595  (
    .a({\u2_Display/n889 ,\u2_Display/n891 }),
    .b({\u2_Display/n888 ,\u2_Display/n890 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add32/c15 ),
    .f({\u2_Display/n909 [17],\u2_Display/n909 [15]}),
    .fco(\u2_Display/add32/c19 ),
    .fx({\u2_Display/n909 [18],\u2_Display/n909 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u19_al_u4596  (
    .a({\u2_Display/n885 ,\u2_Display/n887 }),
    .b({\u2_Display/n884 ,\u2_Display/n886 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add32/c19 ),
    .f({\u2_Display/n909 [21],\u2_Display/n909 [19]}),
    .fco(\u2_Display/add32/c23 ),
    .fx({\u2_Display/n909 [22],\u2_Display/n909 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u23_al_u4597  (
    .a({\u2_Display/n881 ,\u2_Display/n883 }),
    .b({\u2_Display/n880 ,\u2_Display/n882 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add32/c23 ),
    .f({\u2_Display/n909 [25],\u2_Display/n909 [23]}),
    .fco(\u2_Display/add32/c27 ),
    .fx({\u2_Display/n909 [26],\u2_Display/n909 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u27_al_u4598  (
    .a({\u2_Display/n877 ,\u2_Display/n879 }),
    .b({\u2_Display/n876 ,\u2_Display/n878 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add32/c27 ),
    .f({\u2_Display/n909 [29],\u2_Display/n909 [27]}),
    .fco(\u2_Display/add32/c31 ),
    .fx({\u2_Display/n909 [30],\u2_Display/n909 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u31_al_u4599  (
    .a({open_n14391,\u2_Display/n875 }),
    .c(2'b00),
    .d({open_n14396,1'b1}),
    .fci(\u2_Display/add32/c31 ),
    .f({open_n14413,\u2_Display/n909 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u3_al_u4592  (
    .a({\u2_Display/n901 ,\u2_Display/n903 }),
    .b({\u2_Display/n900 ,\u2_Display/n902 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add32/c3 ),
    .f({\u2_Display/n909 [5],\u2_Display/n909 [3]}),
    .fco(\u2_Display/add32/c7 ),
    .fx({\u2_Display/n909 [6],\u2_Display/n909 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/u7_al_u4593  (
    .a({\u2_Display/n897 ,\u2_Display/n899 }),
    .b({\u2_Display/n896 ,\u2_Display/n898 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add32/c7 ),
    .f({\u2_Display/n909 [9],\u2_Display/n909 [7]}),
    .fco(\u2_Display/add32/c11 ),
    .fx({\u2_Display/n909 [10],\u2_Display/n909 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add32/ucin_al_u4591"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add32/ucin_al_u4591  (
    .a({\u2_Display/n905 ,1'b1}),
    .b({\u2_Display/n904 ,\u2_Display/n906 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n909 [1],open_n14472}),
    .fco(\u2_Display/add32/c3 ),
    .fx({\u2_Display/n909 [2],\u2_Display/n909 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u11_al_u4603  (
    .a({\u2_Display/n928 ,\u2_Display/n930 }),
    .b({\u2_Display/n927 ,\u2_Display/n929 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add33/c11 ),
    .f({\u2_Display/n944 [13],\u2_Display/n944 [11]}),
    .fco(\u2_Display/add33/c15 ),
    .fx({\u2_Display/n944 [14],\u2_Display/n944 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u15_al_u4604  (
    .a({\u2_Display/n924 ,\u2_Display/n926 }),
    .b({\u2_Display/n923 ,\u2_Display/n925 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add33/c15 ),
    .f({\u2_Display/n944 [17],\u2_Display/n944 [15]}),
    .fco(\u2_Display/add33/c19 ),
    .fx({\u2_Display/n944 [18],\u2_Display/n944 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u19_al_u4605  (
    .a({\u2_Display/n920 ,\u2_Display/n922 }),
    .b({\u2_Display/n919 ,\u2_Display/n921 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add33/c19 ),
    .f({\u2_Display/n944 [21],\u2_Display/n944 [19]}),
    .fco(\u2_Display/add33/c23 ),
    .fx({\u2_Display/n944 [22],\u2_Display/n944 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u23_al_u4606  (
    .a({\u2_Display/n916 ,\u2_Display/n918 }),
    .b({\u2_Display/n915 ,\u2_Display/n917 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add33/c23 ),
    .f({\u2_Display/n944 [25],\u2_Display/n944 [23]}),
    .fco(\u2_Display/add33/c27 ),
    .fx({\u2_Display/n944 [26],\u2_Display/n944 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u27_al_u4607  (
    .a({\u2_Display/n912 ,\u2_Display/n914 }),
    .b({\u2_Display/n911 ,\u2_Display/n913 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add33/c27 ),
    .f({\u2_Display/n944 [29],\u2_Display/n944 [27]}),
    .fco(\u2_Display/add33/c31 ),
    .fx({\u2_Display/n944 [30],\u2_Display/n944 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u31_al_u4608  (
    .a({open_n14565,\u2_Display/n910 }),
    .c(2'b00),
    .d({open_n14570,1'b1}),
    .fci(\u2_Display/add33/c31 ),
    .f({open_n14587,\u2_Display/n944 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u3_al_u4601  (
    .a({\u2_Display/n936 ,\u2_Display/n938 }),
    .b({\u2_Display/n935 ,\u2_Display/n937 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add33/c3 ),
    .f({\u2_Display/n944 [5],\u2_Display/n944 [3]}),
    .fco(\u2_Display/add33/c7 ),
    .fx({\u2_Display/n944 [6],\u2_Display/n944 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/u7_al_u4602  (
    .a({\u2_Display/n932 ,\u2_Display/n934 }),
    .b({\u2_Display/n931 ,\u2_Display/n933 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add33/c7 ),
    .f({\u2_Display/n944 [9],\u2_Display/n944 [7]}),
    .fco(\u2_Display/add33/c11 ),
    .fx({\u2_Display/n944 [10],\u2_Display/n944 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add33/ucin_al_u4600"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add33/ucin_al_u4600  (
    .a({\u2_Display/n940 ,1'b1}),
    .b({\u2_Display/n939 ,\u2_Display/n941 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n944 [1],open_n14646}),
    .fco(\u2_Display/add33/c3 ),
    .fx({\u2_Display/n944 [2],\u2_Display/n944 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u11_al_u4612  (
    .a({\u2_Display/n963 ,\u2_Display/n965 }),
    .b({\u2_Display/n962 ,\u2_Display/n964 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add34/c11 ),
    .f({\u2_Display/n979 [13],\u2_Display/n979 [11]}),
    .fco(\u2_Display/add34/c15 ),
    .fx({\u2_Display/n979 [14],\u2_Display/n979 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u15_al_u4613  (
    .a({\u2_Display/n959 ,\u2_Display/n961 }),
    .b({\u2_Display/n958 ,\u2_Display/n960 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add34/c15 ),
    .f({\u2_Display/n979 [17],\u2_Display/n979 [15]}),
    .fco(\u2_Display/add34/c19 ),
    .fx({\u2_Display/n979 [18],\u2_Display/n979 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u19_al_u4614  (
    .a({\u2_Display/n955 ,\u2_Display/n957 }),
    .b({\u2_Display/n954 ,\u2_Display/n956 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add34/c19 ),
    .f({\u2_Display/n979 [21],\u2_Display/n979 [19]}),
    .fco(\u2_Display/add34/c23 ),
    .fx({\u2_Display/n979 [22],\u2_Display/n979 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u23_al_u4615  (
    .a({\u2_Display/n951 ,\u2_Display/n953 }),
    .b({\u2_Display/n950 ,\u2_Display/n952 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add34/c23 ),
    .f({\u2_Display/n979 [25],\u2_Display/n979 [23]}),
    .fco(\u2_Display/add34/c27 ),
    .fx({\u2_Display/n979 [26],\u2_Display/n979 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u27_al_u4616  (
    .a({\u2_Display/n947 ,\u2_Display/n949 }),
    .b({\u2_Display/n946 ,\u2_Display/n948 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add34/c27 ),
    .f({\u2_Display/n979 [29],\u2_Display/n979 [27]}),
    .fco(\u2_Display/add34/c31 ),
    .fx({\u2_Display/n979 [30],\u2_Display/n979 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u31_al_u4617  (
    .a({open_n14739,\u2_Display/n945 }),
    .c(2'b00),
    .d({open_n14744,1'b1}),
    .fci(\u2_Display/add34/c31 ),
    .f({open_n14761,\u2_Display/n979 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u3_al_u4610  (
    .a({\u2_Display/n971 ,\u2_Display/n973 }),
    .b({\u2_Display/n970 ,\u2_Display/n972 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add34/c3 ),
    .f({\u2_Display/n979 [5],\u2_Display/n979 [3]}),
    .fco(\u2_Display/add34/c7 ),
    .fx({\u2_Display/n979 [6],\u2_Display/n979 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/u7_al_u4611  (
    .a({\u2_Display/n967 ,\u2_Display/n969 }),
    .b({\u2_Display/n966 ,\u2_Display/n968 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add34/c7 ),
    .f({\u2_Display/n979 [9],\u2_Display/n979 [7]}),
    .fco(\u2_Display/add34/c11 ),
    .fx({\u2_Display/n979 [10],\u2_Display/n979 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add34/ucin_al_u4609"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add34/ucin_al_u4609  (
    .a({\u2_Display/n975 ,1'b1}),
    .b({\u2_Display/n974 ,\u2_Display/n976 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n979 [1],open_n14820}),
    .fco(\u2_Display/add34/c3 ),
    .fx({\u2_Display/n979 [2],\u2_Display/n979 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u11_al_u4621  (
    .a({\u2_Display/n998 ,\u2_Display/n1000 }),
    .b({\u2_Display/n997 ,\u2_Display/n999 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add35/c11 ),
    .f({\u2_Display/n1014 [13],\u2_Display/n1014 [11]}),
    .fco(\u2_Display/add35/c15 ),
    .fx({\u2_Display/n1014 [14],\u2_Display/n1014 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u15_al_u4622  (
    .a({\u2_Display/n994 ,\u2_Display/n996 }),
    .b({\u2_Display/n993 ,\u2_Display/n995 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add35/c15 ),
    .f({\u2_Display/n1014 [17],\u2_Display/n1014 [15]}),
    .fco(\u2_Display/add35/c19 ),
    .fx({\u2_Display/n1014 [18],\u2_Display/n1014 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u19_al_u4623  (
    .a({\u2_Display/n990 ,\u2_Display/n992 }),
    .b({\u2_Display/n989 ,\u2_Display/n991 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add35/c19 ),
    .f({\u2_Display/n1014 [21],\u2_Display/n1014 [19]}),
    .fco(\u2_Display/add35/c23 ),
    .fx({\u2_Display/n1014 [22],\u2_Display/n1014 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u23_al_u4624  (
    .a({\u2_Display/n986 ,\u2_Display/n988 }),
    .b({\u2_Display/n985 ,\u2_Display/n987 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add35/c23 ),
    .f({\u2_Display/n1014 [25],\u2_Display/n1014 [23]}),
    .fco(\u2_Display/add35/c27 ),
    .fx({\u2_Display/n1014 [26],\u2_Display/n1014 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u27_al_u4625  (
    .a({\u2_Display/n982 ,\u2_Display/n984 }),
    .b({\u2_Display/n981 ,\u2_Display/n983 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add35/c27 ),
    .f({\u2_Display/n1014 [29],\u2_Display/n1014 [27]}),
    .fco(\u2_Display/add35/c31 ),
    .fx({\u2_Display/n1014 [30],\u2_Display/n1014 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u31_al_u4626  (
    .a({open_n14913,\u2_Display/n980 }),
    .c(2'b00),
    .d({open_n14918,1'b1}),
    .fci(\u2_Display/add35/c31 ),
    .f({open_n14935,\u2_Display/n1014 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u3_al_u4619  (
    .a({\u2_Display/n1006 ,\u2_Display/n1008 }),
    .b({\u2_Display/n1005 ,\u2_Display/n1007 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add35/c3 ),
    .f({\u2_Display/n1014 [5],\u2_Display/n1014 [3]}),
    .fco(\u2_Display/add35/c7 ),
    .fx({\u2_Display/n1014 [6],\u2_Display/n1014 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/u7_al_u4620  (
    .a({\u2_Display/n1002 ,\u2_Display/n1004 }),
    .b({\u2_Display/n1001 ,\u2_Display/n1003 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add35/c7 ),
    .f({\u2_Display/n1014 [9],\u2_Display/n1014 [7]}),
    .fco(\u2_Display/add35/c11 ),
    .fx({\u2_Display/n1014 [10],\u2_Display/n1014 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add35/ucin_al_u4618"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add35/ucin_al_u4618  (
    .a({\u2_Display/n1010 ,1'b1}),
    .b({\u2_Display/n1009 ,\u2_Display/n1011 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1014 [1],open_n14994}),
    .fco(\u2_Display/add35/c3 ),
    .fx({\u2_Display/n1014 [2],\u2_Display/n1014 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u11_al_u4630  (
    .a({\u2_Display/n1033 ,\u2_Display/n1035 }),
    .b({\u2_Display/n1032 ,\u2_Display/n1034 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add36/c11 ),
    .f({\u2_Display/n1049 [13],\u2_Display/n1049 [11]}),
    .fco(\u2_Display/add36/c15 ),
    .fx({\u2_Display/n1049 [14],\u2_Display/n1049 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u15_al_u4631  (
    .a({\u2_Display/n1029 ,\u2_Display/n1031 }),
    .b({\u2_Display/n1028 ,\u2_Display/n1030 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add36/c15 ),
    .f({\u2_Display/n1049 [17],\u2_Display/n1049 [15]}),
    .fco(\u2_Display/add36/c19 ),
    .fx({\u2_Display/n1049 [18],\u2_Display/n1049 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u19_al_u4632  (
    .a({\u2_Display/n1025 ,\u2_Display/n1027 }),
    .b({\u2_Display/n1024 ,\u2_Display/n1026 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add36/c19 ),
    .f({\u2_Display/n1049 [21],\u2_Display/n1049 [19]}),
    .fco(\u2_Display/add36/c23 ),
    .fx({\u2_Display/n1049 [22],\u2_Display/n1049 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u23_al_u4633  (
    .a({\u2_Display/n1021 ,\u2_Display/n1023 }),
    .b({\u2_Display/n1020 ,\u2_Display/n1022 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add36/c23 ),
    .f({\u2_Display/n1049 [25],\u2_Display/n1049 [23]}),
    .fco(\u2_Display/add36/c27 ),
    .fx({\u2_Display/n1049 [26],\u2_Display/n1049 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u27_al_u4634  (
    .a({\u2_Display/n1017 ,\u2_Display/n1019 }),
    .b({\u2_Display/n1016 ,\u2_Display/n1018 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add36/c27 ),
    .f({\u2_Display/n1049 [29],\u2_Display/n1049 [27]}),
    .fco(\u2_Display/add36/c31 ),
    .fx({\u2_Display/n1049 [30],\u2_Display/n1049 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u31_al_u4635  (
    .a({open_n15087,\u2_Display/n1015 }),
    .c(2'b00),
    .d({open_n15092,1'b1}),
    .fci(\u2_Display/add36/c31 ),
    .f({open_n15109,\u2_Display/n1049 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u3_al_u4628  (
    .a({\u2_Display/n1041 ,\u2_Display/n1043 }),
    .b({\u2_Display/n1040 ,\u2_Display/n1042 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add36/c3 ),
    .f({\u2_Display/n1049 [5],\u2_Display/n1049 [3]}),
    .fco(\u2_Display/add36/c7 ),
    .fx({\u2_Display/n1049 [6],\u2_Display/n1049 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/u7_al_u4629  (
    .a({\u2_Display/n1037 ,\u2_Display/n1039 }),
    .b({\u2_Display/n1036 ,\u2_Display/n1038 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b01),
    .fci(\u2_Display/add36/c7 ),
    .f({\u2_Display/n1049 [9],\u2_Display/n1049 [7]}),
    .fco(\u2_Display/add36/c11 ),
    .fx({\u2_Display/n1049 [10],\u2_Display/n1049 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add36/ucin_al_u4627"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add36/ucin_al_u4627  (
    .a({\u2_Display/n1045 ,1'b1}),
    .b({\u2_Display/n1044 ,\u2_Display/n1046 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1049 [1],open_n15168}),
    .fco(\u2_Display/add36/c3 ),
    .fx({\u2_Display/n1049 [2],\u2_Display/n1049 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u11_al_u4639  (
    .a({\u2_Display/n1068 ,\u2_Display/n1070 }),
    .b({\u2_Display/n1067 ,\u2_Display/n1069 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add37/c11 ),
    .f({\u2_Display/n1084 [13],\u2_Display/n1084 [11]}),
    .fco(\u2_Display/add37/c15 ),
    .fx({\u2_Display/n1084 [14],\u2_Display/n1084 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u15_al_u4640  (
    .a({\u2_Display/n1064 ,\u2_Display/n1066 }),
    .b({\u2_Display/n1063 ,\u2_Display/n1065 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add37/c15 ),
    .f({\u2_Display/n1084 [17],\u2_Display/n1084 [15]}),
    .fco(\u2_Display/add37/c19 ),
    .fx({\u2_Display/n1084 [18],\u2_Display/n1084 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u19_al_u4641  (
    .a({\u2_Display/n1060 ,\u2_Display/n1062 }),
    .b({\u2_Display/n1059 ,\u2_Display/n1061 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add37/c19 ),
    .f({\u2_Display/n1084 [21],\u2_Display/n1084 [19]}),
    .fco(\u2_Display/add37/c23 ),
    .fx({\u2_Display/n1084 [22],\u2_Display/n1084 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u23_al_u4642  (
    .a({\u2_Display/n1056 ,\u2_Display/n1058 }),
    .b({\u2_Display/n1055 ,\u2_Display/n1057 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add37/c23 ),
    .f({\u2_Display/n1084 [25],\u2_Display/n1084 [23]}),
    .fco(\u2_Display/add37/c27 ),
    .fx({\u2_Display/n1084 [26],\u2_Display/n1084 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u27_al_u4643  (
    .a({\u2_Display/n1052 ,\u2_Display/n1054 }),
    .b({\u2_Display/n1051 ,\u2_Display/n1053 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add37/c27 ),
    .f({\u2_Display/n1084 [29],\u2_Display/n1084 [27]}),
    .fco(\u2_Display/add37/c31 ),
    .fx({\u2_Display/n1084 [30],\u2_Display/n1084 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u31_al_u4644  (
    .a({open_n15261,\u2_Display/n1050 }),
    .c(2'b00),
    .d({open_n15266,1'b1}),
    .fci(\u2_Display/add37/c31 ),
    .f({open_n15283,\u2_Display/n1084 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u3_al_u4637  (
    .a({\u2_Display/n1076 ,\u2_Display/n1078 }),
    .b({\u2_Display/n1075 ,\u2_Display/n1077 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add37/c3 ),
    .f({\u2_Display/n1084 [5],\u2_Display/n1084 [3]}),
    .fco(\u2_Display/add37/c7 ),
    .fx({\u2_Display/n1084 [6],\u2_Display/n1084 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/u7_al_u4638  (
    .a({\u2_Display/n1072 ,\u2_Display/n1074 }),
    .b({\u2_Display/n1071 ,\u2_Display/n1073 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add37/c7 ),
    .f({\u2_Display/n1084 [9],\u2_Display/n1084 [7]}),
    .fco(\u2_Display/add37/c11 ),
    .fx({\u2_Display/n1084 [10],\u2_Display/n1084 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add37/ucin_al_u4636"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add37/ucin_al_u4636  (
    .a({\u2_Display/n1080 ,1'b1}),
    .b({\u2_Display/n1079 ,\u2_Display/n1081 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1084 [1],open_n15342}),
    .fco(\u2_Display/add37/c3 ),
    .fx({\u2_Display/n1084 [2],\u2_Display/n1084 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u11_al_u4648  (
    .a({\u2_Display/n1103 ,\u2_Display/n1105 }),
    .b({\u2_Display/n1102 ,\u2_Display/n1104 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add38/c11 ),
    .f({\u2_Display/n1119 [13],\u2_Display/n1119 [11]}),
    .fco(\u2_Display/add38/c15 ),
    .fx({\u2_Display/n1119 [14],\u2_Display/n1119 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u15_al_u4649  (
    .a({\u2_Display/n1099 ,\u2_Display/n1101 }),
    .b({\u2_Display/n1098 ,\u2_Display/n1100 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add38/c15 ),
    .f({\u2_Display/n1119 [17],\u2_Display/n1119 [15]}),
    .fco(\u2_Display/add38/c19 ),
    .fx({\u2_Display/n1119 [18],\u2_Display/n1119 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u19_al_u4650  (
    .a({\u2_Display/n1095 ,\u2_Display/n1097 }),
    .b({\u2_Display/n1094 ,\u2_Display/n1096 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add38/c19 ),
    .f({\u2_Display/n1119 [21],\u2_Display/n1119 [19]}),
    .fco(\u2_Display/add38/c23 ),
    .fx({\u2_Display/n1119 [22],\u2_Display/n1119 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u23_al_u4651  (
    .a({\u2_Display/n1091 ,\u2_Display/n1093 }),
    .b({\u2_Display/n1090 ,\u2_Display/n1092 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add38/c23 ),
    .f({\u2_Display/n1119 [25],\u2_Display/n1119 [23]}),
    .fco(\u2_Display/add38/c27 ),
    .fx({\u2_Display/n1119 [26],\u2_Display/n1119 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u27_al_u4652  (
    .a({\u2_Display/n1087 ,\u2_Display/n1089 }),
    .b({\u2_Display/n1086 ,\u2_Display/n1088 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add38/c27 ),
    .f({\u2_Display/n1119 [29],\u2_Display/n1119 [27]}),
    .fco(\u2_Display/add38/c31 ),
    .fx({\u2_Display/n1119 [30],\u2_Display/n1119 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u31_al_u4653  (
    .a({open_n15435,\u2_Display/n1085 }),
    .c(2'b00),
    .d({open_n15440,1'b1}),
    .fci(\u2_Display/add38/c31 ),
    .f({open_n15457,\u2_Display/n1119 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u3_al_u4646  (
    .a({\u2_Display/n1111 ,\u2_Display/n1113 }),
    .b({\u2_Display/n1110 ,\u2_Display/n1112 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add38/c3 ),
    .f({\u2_Display/n1119 [5],\u2_Display/n1119 [3]}),
    .fco(\u2_Display/add38/c7 ),
    .fx({\u2_Display/n1119 [6],\u2_Display/n1119 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/u7_al_u4647  (
    .a({\u2_Display/n1107 ,\u2_Display/n1109 }),
    .b({\u2_Display/n1106 ,\u2_Display/n1108 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add38/c7 ),
    .f({\u2_Display/n1119 [9],\u2_Display/n1119 [7]}),
    .fco(\u2_Display/add38/c11 ),
    .fx({\u2_Display/n1119 [10],\u2_Display/n1119 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add38/ucin_al_u4645"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add38/ucin_al_u4645  (
    .a({\u2_Display/n1115 ,1'b1}),
    .b({\u2_Display/n1114 ,\u2_Display/n1116 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1119 [1],open_n15516}),
    .fco(\u2_Display/add38/c3 ),
    .fx({\u2_Display/n1119 [2],\u2_Display/n1119 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u11_al_u4657  (
    .a({\u2_Display/n1138 ,\u2_Display/n1140 }),
    .b({\u2_Display/n1137 ,\u2_Display/n1139 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add39/c11 ),
    .f({\u2_Display/n1154 [13],\u2_Display/n1154 [11]}),
    .fco(\u2_Display/add39/c15 ),
    .fx({\u2_Display/n1154 [14],\u2_Display/n1154 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u15_al_u4658  (
    .a({\u2_Display/n1134 ,\u2_Display/n1136 }),
    .b({\u2_Display/n1133 ,\u2_Display/n1135 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add39/c15 ),
    .f({\u2_Display/n1154 [17],\u2_Display/n1154 [15]}),
    .fco(\u2_Display/add39/c19 ),
    .fx({\u2_Display/n1154 [18],\u2_Display/n1154 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u19_al_u4659  (
    .a({\u2_Display/n1130 ,\u2_Display/n1132 }),
    .b({\u2_Display/n1129 ,\u2_Display/n1131 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add39/c19 ),
    .f({\u2_Display/n1154 [21],\u2_Display/n1154 [19]}),
    .fco(\u2_Display/add39/c23 ),
    .fx({\u2_Display/n1154 [22],\u2_Display/n1154 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u23_al_u4660  (
    .a({\u2_Display/n1126 ,\u2_Display/n1128 }),
    .b({\u2_Display/n1125 ,\u2_Display/n1127 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add39/c23 ),
    .f({\u2_Display/n1154 [25],\u2_Display/n1154 [23]}),
    .fco(\u2_Display/add39/c27 ),
    .fx({\u2_Display/n1154 [26],\u2_Display/n1154 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u27_al_u4661  (
    .a({\u2_Display/n1122 ,\u2_Display/n1124 }),
    .b({\u2_Display/n1121 ,\u2_Display/n1123 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add39/c27 ),
    .f({\u2_Display/n1154 [29],\u2_Display/n1154 [27]}),
    .fco(\u2_Display/add39/c31 ),
    .fx({\u2_Display/n1154 [30],\u2_Display/n1154 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u31_al_u4662  (
    .a({open_n15609,\u2_Display/n1120 }),
    .c(2'b00),
    .d({open_n15614,1'b1}),
    .fci(\u2_Display/add39/c31 ),
    .f({open_n15631,\u2_Display/n1154 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u3_al_u4655  (
    .a({\u2_Display/n1146 ,\u2_Display/n1148 }),
    .b({\u2_Display/n1145 ,\u2_Display/n1147 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b00),
    .fci(\u2_Display/add39/c3 ),
    .f({\u2_Display/n1154 [5],\u2_Display/n1154 [3]}),
    .fco(\u2_Display/add39/c7 ),
    .fx({\u2_Display/n1154 [6],\u2_Display/n1154 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/u7_al_u4656  (
    .a({\u2_Display/n1142 ,\u2_Display/n1144 }),
    .b({\u2_Display/n1141 ,\u2_Display/n1143 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u2_Display/add39/c7 ),
    .f({\u2_Display/n1154 [9],\u2_Display/n1154 [7]}),
    .fco(\u2_Display/add39/c11 ),
    .fx({\u2_Display/n1154 [10],\u2_Display/n1154 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add39/ucin_al_u4654"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add39/ucin_al_u4654  (
    .a({\u2_Display/n1150 ,1'b1}),
    .b({\u2_Display/n1149 ,\u2_Display/n1151 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1154 [1],open_n15690}),
    .fco(\u2_Display/add39/c3 ),
    .fx({\u2_Display/n1154 [2],\u2_Display/n1154 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add40/ucin_al_u5052"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add40/u3_al_u5053  (
    .a({\u2_Display/n1181 ,\u2_Display/n1183 }),
    .b({\u2_Display/n1180 ,\u2_Display/n1182 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b01),
    .fci(\u2_Display/add40/c3 ),
    .f({\u2_Display/n1189 [5],\u2_Display/n1189 [3]}),
    .fco(\u2_Display/add40/c7 ),
    .fx({\u2_Display/n1189 [6],\u2_Display/n1189 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add40/ucin_al_u5052"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add40/u7_al_u5054  (
    .a({\u2_Display/n1177 ,\u2_Display/n1179 }),
    .b({open_n15711,\u2_Display/n1178 }),
    .c(2'b00),
    .d(2'b00),
    .e({open_n15714,1'b0}),
    .fci(\u2_Display/add40/c7 ),
    .f({\u2_Display/n1189 [9],\u2_Display/n1189 [7]}),
    .fx({open_n15730,\u2_Display/n1189 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add40/ucin_al_u5052"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add40/ucin_al_u5052  (
    .a({\u2_Display/n1185 ,1'b1}),
    .b({\u2_Display/n1184 ,\u2_Display/n1186 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1189 [1],open_n15750}),
    .fco(\u2_Display/add40/c3 ),
    .fx({\u2_Display/n1189 [2],\u2_Display/n1189 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add4_2/u0|u2_Display/add4_2/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add4_2/u0|u2_Display/add4_2/ucin  (
    .a(2'b10),
    .b({\u2_Display/i [7],open_n15753}),
    .f({\u2_Display/n94 [0],open_n15773}),
    .fco(\u2_Display/add4_2/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add4_2/u0|u2_Display/add4_2/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add4_2/u2|u2_Display/add4_2/u1  (
    .a(2'b10),
    .b(\u2_Display/i [9:8]),
    .fci(\u2_Display/add4_2/c1 ),
    .f(\u2_Display/n94 [2:1]),
    .fco(\u2_Display/add4_2/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add4_2/u0|u2_Display/add4_2/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add4_2/ucout|u2_Display/add4_2/u3  (
    .a({open_n15800,1'b0}),
    .b({open_n15801,\u2_Display/i [10]}),
    .fci(\u2_Display/add4_2/c3 ),
    .f({\u2_Display/add4_2_co ,\u2_Display/n94 [3]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u11_al_u4666  (
    .a({\u2_Display/counta [13],\u2_Display/counta [11]}),
    .b({\u2_Display/counta [14],\u2_Display/counta [12]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add51/c11 ),
    .f({\u2_Display/n1542 [13],\u2_Display/n1542 [11]}),
    .fco(\u2_Display/add51/c15 ),
    .fx({\u2_Display/n1542 [14],\u2_Display/n1542 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u15_al_u4667  (
    .a({\u2_Display/counta [17],\u2_Display/counta [15]}),
    .b({\u2_Display/counta [18],\u2_Display/counta [16]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add51/c15 ),
    .f({\u2_Display/n1542 [17],\u2_Display/n1542 [15]}),
    .fco(\u2_Display/add51/c19 ),
    .fx({\u2_Display/n1542 [18],\u2_Display/n1542 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u19_al_u4668  (
    .a({\u2_Display/counta [21],\u2_Display/counta [19]}),
    .b({\u2_Display/counta [22],\u2_Display/counta [20]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add51/c19 ),
    .f({\u2_Display/n1542 [21],\u2_Display/n1542 [19]}),
    .fco(\u2_Display/add51/c23 ),
    .fx({\u2_Display/n1542 [22],\u2_Display/n1542 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u23_al_u4669  (
    .a({\u2_Display/counta [25],\u2_Display/counta [23]}),
    .b({\u2_Display/counta [26],\u2_Display/counta [24]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add51/c23 ),
    .f({\u2_Display/n1542 [25],\u2_Display/n1542 [23]}),
    .fco(\u2_Display/add51/c27 ),
    .fx({\u2_Display/n1542 [26],\u2_Display/n1542 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u27_al_u4670  (
    .a({\u2_Display/counta [29],\u2_Display/counta [27]}),
    .b({\u2_Display/counta [30],\u2_Display/counta [28]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add51/c27 ),
    .f({\u2_Display/n1542 [29],\u2_Display/n1542 [27]}),
    .fco(\u2_Display/add51/c31 ),
    .fx({\u2_Display/n1542 [30],\u2_Display/n1542 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u31_al_u4671  (
    .a({open_n15915,\u2_Display/counta [31]}),
    .c(2'b00),
    .d({open_n15920,1'b0}),
    .fci(\u2_Display/add51/c31 ),
    .f({open_n15937,\u2_Display/n1542 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u3_al_u4664  (
    .a({\u2_Display/counta [5],\u2_Display/counta [3]}),
    .b({\u2_Display/counta [6],\u2_Display/counta [4]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add51/c3 ),
    .f({\u2_Display/n1542 [5],\u2_Display/n1542 [3]}),
    .fco(\u2_Display/add51/c7 ),
    .fx({\u2_Display/n1542 [6],\u2_Display/n1542 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/u7_al_u4665  (
    .a({\u2_Display/counta [9],\u2_Display/counta [7]}),
    .b({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add51/c7 ),
    .f({\u2_Display/n1542 [9],\u2_Display/n1542 [7]}),
    .fco(\u2_Display/add51/c11 ),
    .fx({\u2_Display/n1542 [10],\u2_Display/n1542 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add51/ucin_al_u4663"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add51/ucin_al_u4663  (
    .a({\u2_Display/counta [1],1'b1}),
    .b({\u2_Display/counta [2],\u2_Display/counta [0]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1542 [1],open_n15996}),
    .fco(\u2_Display/add51/c3 ),
    .fx({\u2_Display/n1542 [2],\u2_Display/n1542 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u11_al_u4675  (
    .a({\u2_Display/n1561 ,\u2_Display/n1563 }),
    .b({\u2_Display/n1560 ,\u2_Display/n1562 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add52/c11 ),
    .f({\u2_Display/n1577 [13],\u2_Display/n1577 [11]}),
    .fco(\u2_Display/add52/c15 ),
    .fx({\u2_Display/n1577 [14],\u2_Display/n1577 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u15_al_u4676  (
    .a({\u2_Display/n1557 ,\u2_Display/n1559 }),
    .b({\u2_Display/n1556 ,\u2_Display/n1558 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add52/c15 ),
    .f({\u2_Display/n1577 [17],\u2_Display/n1577 [15]}),
    .fco(\u2_Display/add52/c19 ),
    .fx({\u2_Display/n1577 [18],\u2_Display/n1577 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u19_al_u4677  (
    .a({\u2_Display/n1553 ,\u2_Display/n1555 }),
    .b({\u2_Display/n1552 ,\u2_Display/n1554 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add52/c19 ),
    .f({\u2_Display/n1577 [21],\u2_Display/n1577 [19]}),
    .fco(\u2_Display/add52/c23 ),
    .fx({\u2_Display/n1577 [22],\u2_Display/n1577 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u23_al_u4678  (
    .a({\u2_Display/n1549 ,\u2_Display/n1551 }),
    .b({\u2_Display/n1548 ,\u2_Display/n1550 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add52/c23 ),
    .f({\u2_Display/n1577 [25],\u2_Display/n1577 [23]}),
    .fco(\u2_Display/add52/c27 ),
    .fx({\u2_Display/n1577 [26],\u2_Display/n1577 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u27_al_u4679  (
    .a({\u2_Display/n1545 ,\u2_Display/n1547 }),
    .b({\u2_Display/n1544 ,\u2_Display/n1546 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add52/c27 ),
    .f({\u2_Display/n1577 [29],\u2_Display/n1577 [27]}),
    .fco(\u2_Display/add52/c31 ),
    .fx({\u2_Display/n1577 [30],\u2_Display/n1577 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u31_al_u4680  (
    .a({open_n16089,\u2_Display/n1543 }),
    .c(2'b00),
    .d({open_n16094,1'b1}),
    .fci(\u2_Display/add52/c31 ),
    .f({open_n16111,\u2_Display/n1577 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u3_al_u4673  (
    .a({\u2_Display/n1569 ,\u2_Display/n1571 }),
    .b({\u2_Display/n1568 ,\u2_Display/n1570 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add52/c3 ),
    .f({\u2_Display/n1577 [5],\u2_Display/n1577 [3]}),
    .fco(\u2_Display/add52/c7 ),
    .fx({\u2_Display/n1577 [6],\u2_Display/n1577 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/u7_al_u4674  (
    .a({\u2_Display/n1565 ,\u2_Display/n1567 }),
    .b({\u2_Display/n1564 ,\u2_Display/n1566 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add52/c7 ),
    .f({\u2_Display/n1577 [9],\u2_Display/n1577 [7]}),
    .fco(\u2_Display/add52/c11 ),
    .fx({\u2_Display/n1577 [10],\u2_Display/n1577 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add52/ucin_al_u4672"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add52/ucin_al_u4672  (
    .a({\u2_Display/n1573 ,1'b1}),
    .b({\u2_Display/n1572 ,\u2_Display/n1574 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1577 [1],open_n16170}),
    .fco(\u2_Display/add52/c3 ),
    .fx({\u2_Display/n1577 [2],\u2_Display/n1577 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u11_al_u4684  (
    .a({\u2_Display/n1596 ,\u2_Display/n1598 }),
    .b({\u2_Display/n1595 ,\u2_Display/n1597 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add53/c11 ),
    .f({\u2_Display/n1612 [13],\u2_Display/n1612 [11]}),
    .fco(\u2_Display/add53/c15 ),
    .fx({\u2_Display/n1612 [14],\u2_Display/n1612 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u15_al_u4685  (
    .a({\u2_Display/n1592 ,\u2_Display/n1594 }),
    .b({\u2_Display/n1591 ,\u2_Display/n1593 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add53/c15 ),
    .f({\u2_Display/n1612 [17],\u2_Display/n1612 [15]}),
    .fco(\u2_Display/add53/c19 ),
    .fx({\u2_Display/n1612 [18],\u2_Display/n1612 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u19_al_u4686  (
    .a({\u2_Display/n1588 ,\u2_Display/n1590 }),
    .b({\u2_Display/n1587 ,\u2_Display/n1589 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add53/c19 ),
    .f({\u2_Display/n1612 [21],\u2_Display/n1612 [19]}),
    .fco(\u2_Display/add53/c23 ),
    .fx({\u2_Display/n1612 [22],\u2_Display/n1612 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u23_al_u4687  (
    .a({\u2_Display/n1584 ,\u2_Display/n1586 }),
    .b({\u2_Display/n1583 ,\u2_Display/n1585 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add53/c23 ),
    .f({\u2_Display/n1612 [25],\u2_Display/n1612 [23]}),
    .fco(\u2_Display/add53/c27 ),
    .fx({\u2_Display/n1612 [26],\u2_Display/n1612 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u27_al_u4688  (
    .a({\u2_Display/n1580 ,\u2_Display/n1582 }),
    .b({\u2_Display/n1579 ,\u2_Display/n1581 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add53/c27 ),
    .f({\u2_Display/n1612 [29],\u2_Display/n1612 [27]}),
    .fco(\u2_Display/add53/c31 ),
    .fx({\u2_Display/n1612 [30],\u2_Display/n1612 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u31_al_u4689  (
    .a({open_n16263,\u2_Display/n1578 }),
    .c(2'b00),
    .d({open_n16268,1'b1}),
    .fci(\u2_Display/add53/c31 ),
    .f({open_n16285,\u2_Display/n1612 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u3_al_u4682  (
    .a({\u2_Display/n1604 ,\u2_Display/n1606 }),
    .b({\u2_Display/n1603 ,\u2_Display/n1605 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add53/c3 ),
    .f({\u2_Display/n1612 [5],\u2_Display/n1612 [3]}),
    .fco(\u2_Display/add53/c7 ),
    .fx({\u2_Display/n1612 [6],\u2_Display/n1612 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/u7_al_u4683  (
    .a({\u2_Display/n1600 ,\u2_Display/n1602 }),
    .b({\u2_Display/n1599 ,\u2_Display/n1601 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add53/c7 ),
    .f({\u2_Display/n1612 [9],\u2_Display/n1612 [7]}),
    .fco(\u2_Display/add53/c11 ),
    .fx({\u2_Display/n1612 [10],\u2_Display/n1612 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add53/ucin_al_u4681"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add53/ucin_al_u4681  (
    .a({\u2_Display/n1608 ,1'b1}),
    .b({\u2_Display/n1607 ,\u2_Display/n1609 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1612 [1],open_n16344}),
    .fco(\u2_Display/add53/c3 ),
    .fx({\u2_Display/n1612 [2],\u2_Display/n1612 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u11_al_u4693  (
    .a({\u2_Display/n1631 ,\u2_Display/n1633 }),
    .b({\u2_Display/n1630 ,\u2_Display/n1632 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add54/c11 ),
    .f({\u2_Display/n1647 [13],\u2_Display/n1647 [11]}),
    .fco(\u2_Display/add54/c15 ),
    .fx({\u2_Display/n1647 [14],\u2_Display/n1647 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u15_al_u4694  (
    .a({\u2_Display/n1627 ,\u2_Display/n1629 }),
    .b({\u2_Display/n1626 ,\u2_Display/n1628 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add54/c15 ),
    .f({\u2_Display/n1647 [17],\u2_Display/n1647 [15]}),
    .fco(\u2_Display/add54/c19 ),
    .fx({\u2_Display/n1647 [18],\u2_Display/n1647 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u19_al_u4695  (
    .a({\u2_Display/n1623 ,\u2_Display/n1625 }),
    .b({\u2_Display/n1622 ,\u2_Display/n1624 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add54/c19 ),
    .f({\u2_Display/n1647 [21],\u2_Display/n1647 [19]}),
    .fco(\u2_Display/add54/c23 ),
    .fx({\u2_Display/n1647 [22],\u2_Display/n1647 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u23_al_u4696  (
    .a({\u2_Display/n1619 ,\u2_Display/n1621 }),
    .b({\u2_Display/n1618 ,\u2_Display/n1620 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add54/c23 ),
    .f({\u2_Display/n1647 [25],\u2_Display/n1647 [23]}),
    .fco(\u2_Display/add54/c27 ),
    .fx({\u2_Display/n1647 [26],\u2_Display/n1647 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u27_al_u4697  (
    .a({\u2_Display/n1615 ,\u2_Display/n1617 }),
    .b({\u2_Display/n1614 ,\u2_Display/n1616 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add54/c27 ),
    .f({\u2_Display/n1647 [29],\u2_Display/n1647 [27]}),
    .fco(\u2_Display/add54/c31 ),
    .fx({\u2_Display/n1647 [30],\u2_Display/n1647 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u31_al_u4698  (
    .a({open_n16437,\u2_Display/n1613 }),
    .c(2'b00),
    .d({open_n16442,1'b1}),
    .fci(\u2_Display/add54/c31 ),
    .f({open_n16459,\u2_Display/n1647 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u3_al_u4691  (
    .a({\u2_Display/n1639 ,\u2_Display/n1641 }),
    .b({\u2_Display/n1638 ,\u2_Display/n1640 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add54/c3 ),
    .f({\u2_Display/n1647 [5],\u2_Display/n1647 [3]}),
    .fco(\u2_Display/add54/c7 ),
    .fx({\u2_Display/n1647 [6],\u2_Display/n1647 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/u7_al_u4692  (
    .a({\u2_Display/n1635 ,\u2_Display/n1637 }),
    .b({\u2_Display/n1634 ,\u2_Display/n1636 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add54/c7 ),
    .f({\u2_Display/n1647 [9],\u2_Display/n1647 [7]}),
    .fco(\u2_Display/add54/c11 ),
    .fx({\u2_Display/n1647 [10],\u2_Display/n1647 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add54/ucin_al_u4690"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add54/ucin_al_u4690  (
    .a({\u2_Display/n1643 ,1'b1}),
    .b({\u2_Display/n1642 ,\u2_Display/n1644 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1647 [1],open_n16518}),
    .fco(\u2_Display/add54/c3 ),
    .fx({\u2_Display/n1647 [2],\u2_Display/n1647 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u11_al_u4702  (
    .a({\u2_Display/n1666 ,\u2_Display/n1668 }),
    .b({\u2_Display/n1665 ,\u2_Display/n1667 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add55/c11 ),
    .f({\u2_Display/n1682 [13],\u2_Display/n1682 [11]}),
    .fco(\u2_Display/add55/c15 ),
    .fx({\u2_Display/n1682 [14],\u2_Display/n1682 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u15_al_u4703  (
    .a({\u2_Display/n1662 ,\u2_Display/n1664 }),
    .b({\u2_Display/n1661 ,\u2_Display/n1663 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add55/c15 ),
    .f({\u2_Display/n1682 [17],\u2_Display/n1682 [15]}),
    .fco(\u2_Display/add55/c19 ),
    .fx({\u2_Display/n1682 [18],\u2_Display/n1682 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u19_al_u4704  (
    .a({\u2_Display/n1658 ,\u2_Display/n1660 }),
    .b({\u2_Display/n1657 ,\u2_Display/n1659 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add55/c19 ),
    .f({\u2_Display/n1682 [21],\u2_Display/n1682 [19]}),
    .fco(\u2_Display/add55/c23 ),
    .fx({\u2_Display/n1682 [22],\u2_Display/n1682 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u23_al_u4705  (
    .a({\u2_Display/n1654 ,\u2_Display/n1656 }),
    .b({\u2_Display/n1653 ,\u2_Display/n1655 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add55/c23 ),
    .f({\u2_Display/n1682 [25],\u2_Display/n1682 [23]}),
    .fco(\u2_Display/add55/c27 ),
    .fx({\u2_Display/n1682 [26],\u2_Display/n1682 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u27_al_u4706  (
    .a({\u2_Display/n1650 ,\u2_Display/n1652 }),
    .b({\u2_Display/n1649 ,\u2_Display/n1651 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add55/c27 ),
    .f({\u2_Display/n1682 [29],\u2_Display/n1682 [27]}),
    .fco(\u2_Display/add55/c31 ),
    .fx({\u2_Display/n1682 [30],\u2_Display/n1682 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u31_al_u4707  (
    .a({open_n16611,\u2_Display/n1648 }),
    .c(2'b00),
    .d({open_n16616,1'b1}),
    .fci(\u2_Display/add55/c31 ),
    .f({open_n16633,\u2_Display/n1682 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u3_al_u4700  (
    .a({\u2_Display/n1674 ,\u2_Display/n1676 }),
    .b({\u2_Display/n1673 ,\u2_Display/n1675 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add55/c3 ),
    .f({\u2_Display/n1682 [5],\u2_Display/n1682 [3]}),
    .fco(\u2_Display/add55/c7 ),
    .fx({\u2_Display/n1682 [6],\u2_Display/n1682 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/u7_al_u4701  (
    .a({\u2_Display/n1670 ,\u2_Display/n1672 }),
    .b({\u2_Display/n1669 ,\u2_Display/n1671 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add55/c7 ),
    .f({\u2_Display/n1682 [9],\u2_Display/n1682 [7]}),
    .fco(\u2_Display/add55/c11 ),
    .fx({\u2_Display/n1682 [10],\u2_Display/n1682 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add55/ucin_al_u4699"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add55/ucin_al_u4699  (
    .a({\u2_Display/n1678 ,1'b1}),
    .b({\u2_Display/n1677 ,\u2_Display/n1679 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1682 [1],open_n16692}),
    .fco(\u2_Display/add55/c3 ),
    .fx({\u2_Display/n1682 [2],\u2_Display/n1682 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u11_al_u4711  (
    .a({\u2_Display/n1701 ,\u2_Display/n1703 }),
    .b({\u2_Display/n1700 ,\u2_Display/n1702 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add56/c11 ),
    .f({\u2_Display/n1717 [13],\u2_Display/n1717 [11]}),
    .fco(\u2_Display/add56/c15 ),
    .fx({\u2_Display/n1717 [14],\u2_Display/n1717 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u15_al_u4712  (
    .a({\u2_Display/n1697 ,\u2_Display/n1699 }),
    .b({\u2_Display/n1696 ,\u2_Display/n1698 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add56/c15 ),
    .f({\u2_Display/n1717 [17],\u2_Display/n1717 [15]}),
    .fco(\u2_Display/add56/c19 ),
    .fx({\u2_Display/n1717 [18],\u2_Display/n1717 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u19_al_u4713  (
    .a({\u2_Display/n1693 ,\u2_Display/n1695 }),
    .b({\u2_Display/n1692 ,\u2_Display/n1694 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add56/c19 ),
    .f({\u2_Display/n1717 [21],\u2_Display/n1717 [19]}),
    .fco(\u2_Display/add56/c23 ),
    .fx({\u2_Display/n1717 [22],\u2_Display/n1717 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u23_al_u4714  (
    .a({\u2_Display/n1689 ,\u2_Display/n1691 }),
    .b({\u2_Display/n1688 ,\u2_Display/n1690 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add56/c23 ),
    .f({\u2_Display/n1717 [25],\u2_Display/n1717 [23]}),
    .fco(\u2_Display/add56/c27 ),
    .fx({\u2_Display/n1717 [26],\u2_Display/n1717 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u27_al_u4715  (
    .a({\u2_Display/n1685 ,\u2_Display/n1687 }),
    .b({\u2_Display/n1684 ,\u2_Display/n1686 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add56/c27 ),
    .f({\u2_Display/n1717 [29],\u2_Display/n1717 [27]}),
    .fco(\u2_Display/add56/c31 ),
    .fx({\u2_Display/n1717 [30],\u2_Display/n1717 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u31_al_u4716  (
    .a({open_n16785,\u2_Display/n1683 }),
    .c(2'b00),
    .d({open_n16790,1'b1}),
    .fci(\u2_Display/add56/c31 ),
    .f({open_n16807,\u2_Display/n1717 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u3_al_u4709  (
    .a({\u2_Display/n1709 ,\u2_Display/n1711 }),
    .b({\u2_Display/n1708 ,\u2_Display/n1710 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add56/c3 ),
    .f({\u2_Display/n1717 [5],\u2_Display/n1717 [3]}),
    .fco(\u2_Display/add56/c7 ),
    .fx({\u2_Display/n1717 [6],\u2_Display/n1717 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/u7_al_u4710  (
    .a({\u2_Display/n1705 ,\u2_Display/n1707 }),
    .b({\u2_Display/n1704 ,\u2_Display/n1706 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add56/c7 ),
    .f({\u2_Display/n1717 [9],\u2_Display/n1717 [7]}),
    .fco(\u2_Display/add56/c11 ),
    .fx({\u2_Display/n1717 [10],\u2_Display/n1717 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add56/ucin_al_u4708"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add56/ucin_al_u4708  (
    .a({\u2_Display/n1713 ,1'b1}),
    .b({\u2_Display/n1712 ,\u2_Display/n1714 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1717 [1],open_n16866}),
    .fco(\u2_Display/add56/c3 ),
    .fx({\u2_Display/n1717 [2],\u2_Display/n1717 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u11_al_u4720  (
    .a({\u2_Display/n1736 ,\u2_Display/n1738 }),
    .b({\u2_Display/n1735 ,\u2_Display/n1737 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add57/c11 ),
    .f({\u2_Display/n1752 [13],\u2_Display/n1752 [11]}),
    .fco(\u2_Display/add57/c15 ),
    .fx({\u2_Display/n1752 [14],\u2_Display/n1752 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u15_al_u4721  (
    .a({\u2_Display/n1732 ,\u2_Display/n1734 }),
    .b({\u2_Display/n1731 ,\u2_Display/n1733 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add57/c15 ),
    .f({\u2_Display/n1752 [17],\u2_Display/n1752 [15]}),
    .fco(\u2_Display/add57/c19 ),
    .fx({\u2_Display/n1752 [18],\u2_Display/n1752 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u19_al_u4722  (
    .a({\u2_Display/n1728 ,\u2_Display/n1730 }),
    .b({\u2_Display/n1727 ,\u2_Display/n1729 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add57/c19 ),
    .f({\u2_Display/n1752 [21],\u2_Display/n1752 [19]}),
    .fco(\u2_Display/add57/c23 ),
    .fx({\u2_Display/n1752 [22],\u2_Display/n1752 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u23_al_u4723  (
    .a({\u2_Display/n1724 ,\u2_Display/n1726 }),
    .b({\u2_Display/n1723 ,\u2_Display/n1725 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add57/c23 ),
    .f({\u2_Display/n1752 [25],\u2_Display/n1752 [23]}),
    .fco(\u2_Display/add57/c27 ),
    .fx({\u2_Display/n1752 [26],\u2_Display/n1752 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u27_al_u4724  (
    .a({\u2_Display/n1720 ,\u2_Display/n1722 }),
    .b({\u2_Display/n1719 ,\u2_Display/n1721 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add57/c27 ),
    .f({\u2_Display/n1752 [29],\u2_Display/n1752 [27]}),
    .fco(\u2_Display/add57/c31 ),
    .fx({\u2_Display/n1752 [30],\u2_Display/n1752 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u31_al_u4725  (
    .a({open_n16959,\u2_Display/n1718 }),
    .c(2'b00),
    .d({open_n16964,1'b1}),
    .fci(\u2_Display/add57/c31 ),
    .f({open_n16981,\u2_Display/n1752 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u3_al_u4718  (
    .a({\u2_Display/n1744 ,\u2_Display/n1746 }),
    .b({\u2_Display/n1743 ,\u2_Display/n1745 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add57/c3 ),
    .f({\u2_Display/n1752 [5],\u2_Display/n1752 [3]}),
    .fco(\u2_Display/add57/c7 ),
    .fx({\u2_Display/n1752 [6],\u2_Display/n1752 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/u7_al_u4719  (
    .a({\u2_Display/n1740 ,\u2_Display/n1742 }),
    .b({\u2_Display/n1739 ,\u2_Display/n1741 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add57/c7 ),
    .f({\u2_Display/n1752 [9],\u2_Display/n1752 [7]}),
    .fco(\u2_Display/add57/c11 ),
    .fx({\u2_Display/n1752 [10],\u2_Display/n1752 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add57/ucin_al_u4717"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add57/ucin_al_u4717  (
    .a({\u2_Display/n1748 ,1'b1}),
    .b({\u2_Display/n1747 ,\u2_Display/n1749 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1752 [1],open_n17040}),
    .fco(\u2_Display/add57/c3 ),
    .fx({\u2_Display/n1752 [2],\u2_Display/n1752 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u11_al_u4729  (
    .a({\u2_Display/n1771 ,\u2_Display/n1773 }),
    .b({\u2_Display/n1770 ,\u2_Display/n1772 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add58/c11 ),
    .f({\u2_Display/n1787 [13],\u2_Display/n1787 [11]}),
    .fco(\u2_Display/add58/c15 ),
    .fx({\u2_Display/n1787 [14],\u2_Display/n1787 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u15_al_u4730  (
    .a({\u2_Display/n1767 ,\u2_Display/n1769 }),
    .b({\u2_Display/n1766 ,\u2_Display/n1768 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add58/c15 ),
    .f({\u2_Display/n1787 [17],\u2_Display/n1787 [15]}),
    .fco(\u2_Display/add58/c19 ),
    .fx({\u2_Display/n1787 [18],\u2_Display/n1787 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u19_al_u4731  (
    .a({\u2_Display/n1763 ,\u2_Display/n1765 }),
    .b({\u2_Display/n1762 ,\u2_Display/n1764 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add58/c19 ),
    .f({\u2_Display/n1787 [21],\u2_Display/n1787 [19]}),
    .fco(\u2_Display/add58/c23 ),
    .fx({\u2_Display/n1787 [22],\u2_Display/n1787 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u23_al_u4732  (
    .a({\u2_Display/n1759 ,\u2_Display/n1761 }),
    .b({\u2_Display/n1758 ,\u2_Display/n1760 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add58/c23 ),
    .f({\u2_Display/n1787 [25],\u2_Display/n1787 [23]}),
    .fco(\u2_Display/add58/c27 ),
    .fx({\u2_Display/n1787 [26],\u2_Display/n1787 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u27_al_u4733  (
    .a({\u2_Display/n1755 ,\u2_Display/n1757 }),
    .b({\u2_Display/n1754 ,\u2_Display/n1756 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add58/c27 ),
    .f({\u2_Display/n1787 [29],\u2_Display/n1787 [27]}),
    .fco(\u2_Display/add58/c31 ),
    .fx({\u2_Display/n1787 [30],\u2_Display/n1787 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u31_al_u4734  (
    .a({open_n17133,\u2_Display/n1753 }),
    .c(2'b00),
    .d({open_n17138,1'b1}),
    .fci(\u2_Display/add58/c31 ),
    .f({open_n17155,\u2_Display/n1787 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u3_al_u4727  (
    .a({\u2_Display/n1779 ,\u2_Display/n1781 }),
    .b({\u2_Display/n1778 ,\u2_Display/n1780 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add58/c3 ),
    .f({\u2_Display/n1787 [5],\u2_Display/n1787 [3]}),
    .fco(\u2_Display/add58/c7 ),
    .fx({\u2_Display/n1787 [6],\u2_Display/n1787 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/u7_al_u4728  (
    .a({\u2_Display/n1775 ,\u2_Display/n1777 }),
    .b({\u2_Display/n1774 ,\u2_Display/n1776 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add58/c7 ),
    .f({\u2_Display/n1787 [9],\u2_Display/n1787 [7]}),
    .fco(\u2_Display/add58/c11 ),
    .fx({\u2_Display/n1787 [10],\u2_Display/n1787 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add58/ucin_al_u4726"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add58/ucin_al_u4726  (
    .a({\u2_Display/n1783 ,1'b1}),
    .b({\u2_Display/n1782 ,\u2_Display/n1784 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1787 [1],open_n17214}),
    .fco(\u2_Display/add58/c3 ),
    .fx({\u2_Display/n1787 [2],\u2_Display/n1787 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u11_al_u4738  (
    .a({\u2_Display/n1806 ,\u2_Display/n1808 }),
    .b({\u2_Display/n1805 ,\u2_Display/n1807 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add59/c11 ),
    .f({\u2_Display/n1822 [13],\u2_Display/n1822 [11]}),
    .fco(\u2_Display/add59/c15 ),
    .fx({\u2_Display/n1822 [14],\u2_Display/n1822 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u15_al_u4739  (
    .a({\u2_Display/n1802 ,\u2_Display/n1804 }),
    .b({\u2_Display/n1801 ,\u2_Display/n1803 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add59/c15 ),
    .f({\u2_Display/n1822 [17],\u2_Display/n1822 [15]}),
    .fco(\u2_Display/add59/c19 ),
    .fx({\u2_Display/n1822 [18],\u2_Display/n1822 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u19_al_u4740  (
    .a({\u2_Display/n1798 ,\u2_Display/n1800 }),
    .b({\u2_Display/n1797 ,\u2_Display/n1799 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add59/c19 ),
    .f({\u2_Display/n1822 [21],\u2_Display/n1822 [19]}),
    .fco(\u2_Display/add59/c23 ),
    .fx({\u2_Display/n1822 [22],\u2_Display/n1822 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u23_al_u4741  (
    .a({\u2_Display/n1794 ,\u2_Display/n1796 }),
    .b({\u2_Display/n1793 ,\u2_Display/n1795 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add59/c23 ),
    .f({\u2_Display/n1822 [25],\u2_Display/n1822 [23]}),
    .fco(\u2_Display/add59/c27 ),
    .fx({\u2_Display/n1822 [26],\u2_Display/n1822 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u27_al_u4742  (
    .a({\u2_Display/n1790 ,\u2_Display/n1792 }),
    .b({\u2_Display/n1789 ,\u2_Display/n1791 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add59/c27 ),
    .f({\u2_Display/n1822 [29],\u2_Display/n1822 [27]}),
    .fco(\u2_Display/add59/c31 ),
    .fx({\u2_Display/n1822 [30],\u2_Display/n1822 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u31_al_u4743  (
    .a({open_n17307,\u2_Display/n1788 }),
    .c(2'b00),
    .d({open_n17312,1'b1}),
    .fci(\u2_Display/add59/c31 ),
    .f({open_n17329,\u2_Display/n1822 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u3_al_u4736  (
    .a({\u2_Display/n1814 ,\u2_Display/n1816 }),
    .b({\u2_Display/n1813 ,\u2_Display/n1815 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add59/c3 ),
    .f({\u2_Display/n1822 [5],\u2_Display/n1822 [3]}),
    .fco(\u2_Display/add59/c7 ),
    .fx({\u2_Display/n1822 [6],\u2_Display/n1822 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/u7_al_u4737  (
    .a({\u2_Display/n1810 ,\u2_Display/n1812 }),
    .b({\u2_Display/n1809 ,\u2_Display/n1811 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add59/c7 ),
    .f({\u2_Display/n1822 [9],\u2_Display/n1822 [7]}),
    .fco(\u2_Display/add59/c11 ),
    .fx({\u2_Display/n1822 [10],\u2_Display/n1822 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add59/ucin_al_u4735"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add59/ucin_al_u4735  (
    .a({\u2_Display/n1818 ,1'b1}),
    .b({\u2_Display/n1817 ,\u2_Display/n1819 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1822 [1],open_n17388}),
    .fco(\u2_Display/add59/c3 ),
    .fx({\u2_Display/n1822 [2],\u2_Display/n1822 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u11_al_u4747  (
    .a({\u2_Display/n1841 ,\u2_Display/n1843 }),
    .b({\u2_Display/n1840 ,\u2_Display/n1842 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add60/c11 ),
    .f({\u2_Display/n1857 [13],\u2_Display/n1857 [11]}),
    .fco(\u2_Display/add60/c15 ),
    .fx({\u2_Display/n1857 [14],\u2_Display/n1857 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u15_al_u4748  (
    .a({\u2_Display/n1837 ,\u2_Display/n1839 }),
    .b({\u2_Display/n1836 ,\u2_Display/n1838 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add60/c15 ),
    .f({\u2_Display/n1857 [17],\u2_Display/n1857 [15]}),
    .fco(\u2_Display/add60/c19 ),
    .fx({\u2_Display/n1857 [18],\u2_Display/n1857 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u19_al_u4749  (
    .a({\u2_Display/n1833 ,\u2_Display/n1835 }),
    .b({\u2_Display/n1832 ,\u2_Display/n1834 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add60/c19 ),
    .f({\u2_Display/n1857 [21],\u2_Display/n1857 [19]}),
    .fco(\u2_Display/add60/c23 ),
    .fx({\u2_Display/n1857 [22],\u2_Display/n1857 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u23_al_u4750  (
    .a({\u2_Display/n1829 ,\u2_Display/n1831 }),
    .b({\u2_Display/n1828 ,\u2_Display/n1830 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add60/c23 ),
    .f({\u2_Display/n1857 [25],\u2_Display/n1857 [23]}),
    .fco(\u2_Display/add60/c27 ),
    .fx({\u2_Display/n1857 [26],\u2_Display/n1857 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u27_al_u4751  (
    .a({\u2_Display/n1825 ,\u2_Display/n1827 }),
    .b({\u2_Display/n1824 ,\u2_Display/n1826 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add60/c27 ),
    .f({\u2_Display/n1857 [29],\u2_Display/n1857 [27]}),
    .fco(\u2_Display/add60/c31 ),
    .fx({\u2_Display/n1857 [30],\u2_Display/n1857 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u31_al_u4752  (
    .a({open_n17481,\u2_Display/n1823 }),
    .c(2'b00),
    .d({open_n17486,1'b1}),
    .fci(\u2_Display/add60/c31 ),
    .f({open_n17503,\u2_Display/n1857 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u3_al_u4745  (
    .a({\u2_Display/n1849 ,\u2_Display/n1851 }),
    .b({\u2_Display/n1848 ,\u2_Display/n1850 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add60/c3 ),
    .f({\u2_Display/n1857 [5],\u2_Display/n1857 [3]}),
    .fco(\u2_Display/add60/c7 ),
    .fx({\u2_Display/n1857 [6],\u2_Display/n1857 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/u7_al_u4746  (
    .a({\u2_Display/n1845 ,\u2_Display/n1847 }),
    .b({\u2_Display/n1844 ,\u2_Display/n1846 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add60/c7 ),
    .f({\u2_Display/n1857 [9],\u2_Display/n1857 [7]}),
    .fco(\u2_Display/add60/c11 ),
    .fx({\u2_Display/n1857 [10],\u2_Display/n1857 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add60/ucin_al_u4744"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add60/ucin_al_u4744  (
    .a({\u2_Display/n1853 ,1'b1}),
    .b({\u2_Display/n1852 ,\u2_Display/n1854 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1857 [1],open_n17562}),
    .fco(\u2_Display/add60/c3 ),
    .fx({\u2_Display/n1857 [2],\u2_Display/n1857 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u11_al_u4756  (
    .a({\u2_Display/n1876 ,\u2_Display/n1878 }),
    .b({\u2_Display/n1875 ,\u2_Display/n1877 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add61/c11 ),
    .f({\u2_Display/n1892 [13],\u2_Display/n1892 [11]}),
    .fco(\u2_Display/add61/c15 ),
    .fx({\u2_Display/n1892 [14],\u2_Display/n1892 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u15_al_u4757  (
    .a({\u2_Display/n1872 ,\u2_Display/n1874 }),
    .b({\u2_Display/n1871 ,\u2_Display/n1873 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add61/c15 ),
    .f({\u2_Display/n1892 [17],\u2_Display/n1892 [15]}),
    .fco(\u2_Display/add61/c19 ),
    .fx({\u2_Display/n1892 [18],\u2_Display/n1892 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u19_al_u4758  (
    .a({\u2_Display/n1868 ,\u2_Display/n1870 }),
    .b({\u2_Display/n1867 ,\u2_Display/n1869 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add61/c19 ),
    .f({\u2_Display/n1892 [21],\u2_Display/n1892 [19]}),
    .fco(\u2_Display/add61/c23 ),
    .fx({\u2_Display/n1892 [22],\u2_Display/n1892 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u23_al_u4759  (
    .a({\u2_Display/n1864 ,\u2_Display/n1866 }),
    .b({\u2_Display/n1863 ,\u2_Display/n1865 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add61/c23 ),
    .f({\u2_Display/n1892 [25],\u2_Display/n1892 [23]}),
    .fco(\u2_Display/add61/c27 ),
    .fx({\u2_Display/n1892 [26],\u2_Display/n1892 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u27_al_u4760  (
    .a({\u2_Display/n1860 ,\u2_Display/n1862 }),
    .b({\u2_Display/n1859 ,\u2_Display/n1861 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add61/c27 ),
    .f({\u2_Display/n1892 [29],\u2_Display/n1892 [27]}),
    .fco(\u2_Display/add61/c31 ),
    .fx({\u2_Display/n1892 [30],\u2_Display/n1892 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u31_al_u4761  (
    .a({open_n17655,\u2_Display/n1858 }),
    .c(2'b00),
    .d({open_n17660,1'b1}),
    .fci(\u2_Display/add61/c31 ),
    .f({open_n17677,\u2_Display/n1892 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u3_al_u4754  (
    .a({\u2_Display/n1884 ,\u2_Display/n1886 }),
    .b({\u2_Display/n1883 ,\u2_Display/n1885 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add61/c3 ),
    .f({\u2_Display/n1892 [5],\u2_Display/n1892 [3]}),
    .fco(\u2_Display/add61/c7 ),
    .fx({\u2_Display/n1892 [6],\u2_Display/n1892 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/u7_al_u4755  (
    .a({\u2_Display/n1880 ,\u2_Display/n1882 }),
    .b({\u2_Display/n1879 ,\u2_Display/n1881 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add61/c7 ),
    .f({\u2_Display/n1892 [9],\u2_Display/n1892 [7]}),
    .fco(\u2_Display/add61/c11 ),
    .fx({\u2_Display/n1892 [10],\u2_Display/n1892 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add61/ucin_al_u4753"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add61/ucin_al_u4753  (
    .a({\u2_Display/n1888 ,1'b1}),
    .b({\u2_Display/n1887 ,\u2_Display/n1889 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1892 [1],open_n17736}),
    .fco(\u2_Display/add61/c3 ),
    .fx({\u2_Display/n1892 [2],\u2_Display/n1892 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u11_al_u4765  (
    .a({\u2_Display/n1911 ,\u2_Display/n1913 }),
    .b({\u2_Display/n1910 ,\u2_Display/n1912 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add62/c11 ),
    .f({\u2_Display/n1927 [13],\u2_Display/n1927 [11]}),
    .fco(\u2_Display/add62/c15 ),
    .fx({\u2_Display/n1927 [14],\u2_Display/n1927 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u15_al_u4766  (
    .a({\u2_Display/n1907 ,\u2_Display/n1909 }),
    .b({\u2_Display/n1906 ,\u2_Display/n1908 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add62/c15 ),
    .f({\u2_Display/n1927 [17],\u2_Display/n1927 [15]}),
    .fco(\u2_Display/add62/c19 ),
    .fx({\u2_Display/n1927 [18],\u2_Display/n1927 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u19_al_u4767  (
    .a({\u2_Display/n1903 ,\u2_Display/n1905 }),
    .b({\u2_Display/n1902 ,\u2_Display/n1904 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add62/c19 ),
    .f({\u2_Display/n1927 [21],\u2_Display/n1927 [19]}),
    .fco(\u2_Display/add62/c23 ),
    .fx({\u2_Display/n1927 [22],\u2_Display/n1927 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u23_al_u4768  (
    .a({\u2_Display/n1899 ,\u2_Display/n1901 }),
    .b({\u2_Display/n1898 ,\u2_Display/n1900 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add62/c23 ),
    .f({\u2_Display/n1927 [25],\u2_Display/n1927 [23]}),
    .fco(\u2_Display/add62/c27 ),
    .fx({\u2_Display/n1927 [26],\u2_Display/n1927 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u27_al_u4769  (
    .a({\u2_Display/n1895 ,\u2_Display/n1897 }),
    .b({\u2_Display/n1894 ,\u2_Display/n1896 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add62/c27 ),
    .f({\u2_Display/n1927 [29],\u2_Display/n1927 [27]}),
    .fco(\u2_Display/add62/c31 ),
    .fx({\u2_Display/n1927 [30],\u2_Display/n1927 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u31_al_u4770  (
    .a({open_n17829,\u2_Display/n1893 }),
    .c(2'b00),
    .d({open_n17834,1'b1}),
    .fci(\u2_Display/add62/c31 ),
    .f({open_n17851,\u2_Display/n1927 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u3_al_u4763  (
    .a({\u2_Display/n1919 ,\u2_Display/n1921 }),
    .b({\u2_Display/n1918 ,\u2_Display/n1920 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add62/c3 ),
    .f({\u2_Display/n1927 [5],\u2_Display/n1927 [3]}),
    .fco(\u2_Display/add62/c7 ),
    .fx({\u2_Display/n1927 [6],\u2_Display/n1927 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/u7_al_u4764  (
    .a({\u2_Display/n1915 ,\u2_Display/n1917 }),
    .b({\u2_Display/n1914 ,\u2_Display/n1916 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add62/c7 ),
    .f({\u2_Display/n1927 [9],\u2_Display/n1927 [7]}),
    .fco(\u2_Display/add62/c11 ),
    .fx({\u2_Display/n1927 [10],\u2_Display/n1927 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add62/ucin_al_u4762"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add62/ucin_al_u4762  (
    .a({\u2_Display/n1923 ,1'b1}),
    .b({\u2_Display/n1922 ,\u2_Display/n1924 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1927 [1],open_n17910}),
    .fco(\u2_Display/add62/c3 ),
    .fx({\u2_Display/n1927 [2],\u2_Display/n1927 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u11_al_u4774  (
    .a({\u2_Display/n1946 ,\u2_Display/n1948 }),
    .b({\u2_Display/n1945 ,\u2_Display/n1947 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add63/c11 ),
    .f({\u2_Display/n1962 [13],\u2_Display/n1962 [11]}),
    .fco(\u2_Display/add63/c15 ),
    .fx({\u2_Display/n1962 [14],\u2_Display/n1962 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u15_al_u4775  (
    .a({\u2_Display/n1942 ,\u2_Display/n1944 }),
    .b({\u2_Display/n1941 ,\u2_Display/n1943 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add63/c15 ),
    .f({\u2_Display/n1962 [17],\u2_Display/n1962 [15]}),
    .fco(\u2_Display/add63/c19 ),
    .fx({\u2_Display/n1962 [18],\u2_Display/n1962 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u19_al_u4776  (
    .a({\u2_Display/n1938 ,\u2_Display/n1940 }),
    .b({\u2_Display/n1937 ,\u2_Display/n1939 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add63/c19 ),
    .f({\u2_Display/n1962 [21],\u2_Display/n1962 [19]}),
    .fco(\u2_Display/add63/c23 ),
    .fx({\u2_Display/n1962 [22],\u2_Display/n1962 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u23_al_u4777  (
    .a({\u2_Display/n1934 ,\u2_Display/n1936 }),
    .b({\u2_Display/n1933 ,\u2_Display/n1935 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add63/c23 ),
    .f({\u2_Display/n1962 [25],\u2_Display/n1962 [23]}),
    .fco(\u2_Display/add63/c27 ),
    .fx({\u2_Display/n1962 [26],\u2_Display/n1962 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u27_al_u4778  (
    .a({\u2_Display/n1930 ,\u2_Display/n1932 }),
    .b({\u2_Display/n1929 ,\u2_Display/n1931 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add63/c27 ),
    .f({\u2_Display/n1962 [29],\u2_Display/n1962 [27]}),
    .fco(\u2_Display/add63/c31 ),
    .fx({\u2_Display/n1962 [30],\u2_Display/n1962 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u31_al_u4779  (
    .a({open_n18003,\u2_Display/n1928 }),
    .c(2'b00),
    .d({open_n18008,1'b1}),
    .fci(\u2_Display/add63/c31 ),
    .f({open_n18025,\u2_Display/n1962 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u3_al_u4772  (
    .a({\u2_Display/n1954 ,\u2_Display/n1956 }),
    .b({\u2_Display/n1953 ,\u2_Display/n1955 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add63/c3 ),
    .f({\u2_Display/n1962 [5],\u2_Display/n1962 [3]}),
    .fco(\u2_Display/add63/c7 ),
    .fx({\u2_Display/n1962 [6],\u2_Display/n1962 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/u7_al_u4773  (
    .a({\u2_Display/n1950 ,\u2_Display/n1952 }),
    .b({\u2_Display/n1949 ,\u2_Display/n1951 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add63/c7 ),
    .f({\u2_Display/n1962 [9],\u2_Display/n1962 [7]}),
    .fco(\u2_Display/add63/c11 ),
    .fx({\u2_Display/n1962 [10],\u2_Display/n1962 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add63/ucin_al_u4771"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add63/ucin_al_u4771  (
    .a({\u2_Display/n1958 ,1'b1}),
    .b({\u2_Display/n1957 ,\u2_Display/n1959 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1962 [1],open_n18084}),
    .fco(\u2_Display/add63/c3 ),
    .fx({\u2_Display/n1962 [2],\u2_Display/n1962 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u11_al_u4783  (
    .a({\u2_Display/n1981 ,\u2_Display/n1983 }),
    .b({\u2_Display/n1980 ,\u2_Display/n1982 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add64/c11 ),
    .f({\u2_Display/n1997 [13],\u2_Display/n1997 [11]}),
    .fco(\u2_Display/add64/c15 ),
    .fx({\u2_Display/n1997 [14],\u2_Display/n1997 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u15_al_u4784  (
    .a({\u2_Display/n1977 ,\u2_Display/n1979 }),
    .b({\u2_Display/n1976 ,\u2_Display/n1978 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add64/c15 ),
    .f({\u2_Display/n1997 [17],\u2_Display/n1997 [15]}),
    .fco(\u2_Display/add64/c19 ),
    .fx({\u2_Display/n1997 [18],\u2_Display/n1997 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u19_al_u4785  (
    .a({\u2_Display/n1973 ,\u2_Display/n1975 }),
    .b({\u2_Display/n1972 ,\u2_Display/n1974 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add64/c19 ),
    .f({\u2_Display/n1997 [21],\u2_Display/n1997 [19]}),
    .fco(\u2_Display/add64/c23 ),
    .fx({\u2_Display/n1997 [22],\u2_Display/n1997 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u23_al_u4786  (
    .a({\u2_Display/n1969 ,\u2_Display/n1971 }),
    .b({\u2_Display/n1968 ,\u2_Display/n1970 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add64/c23 ),
    .f({\u2_Display/n1997 [25],\u2_Display/n1997 [23]}),
    .fco(\u2_Display/add64/c27 ),
    .fx({\u2_Display/n1997 [26],\u2_Display/n1997 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u27_al_u4787  (
    .a({\u2_Display/n1965 ,\u2_Display/n1967 }),
    .b({\u2_Display/n1964 ,\u2_Display/n1966 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add64/c27 ),
    .f({\u2_Display/n1997 [29],\u2_Display/n1997 [27]}),
    .fco(\u2_Display/add64/c31 ),
    .fx({\u2_Display/n1997 [30],\u2_Display/n1997 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u31_al_u4788  (
    .a({open_n18177,\u2_Display/n1963 }),
    .c(2'b00),
    .d({open_n18182,1'b1}),
    .fci(\u2_Display/add64/c31 ),
    .f({open_n18199,\u2_Display/n1997 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u3_al_u4781  (
    .a({\u2_Display/n1989 ,\u2_Display/n1991 }),
    .b({\u2_Display/n1988 ,\u2_Display/n1990 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add64/c3 ),
    .f({\u2_Display/n1997 [5],\u2_Display/n1997 [3]}),
    .fco(\u2_Display/add64/c7 ),
    .fx({\u2_Display/n1997 [6],\u2_Display/n1997 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/u7_al_u4782  (
    .a({\u2_Display/n1985 ,\u2_Display/n1987 }),
    .b({\u2_Display/n1984 ,\u2_Display/n1986 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add64/c7 ),
    .f({\u2_Display/n1997 [9],\u2_Display/n1997 [7]}),
    .fco(\u2_Display/add64/c11 ),
    .fx({\u2_Display/n1997 [10],\u2_Display/n1997 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add64/ucin_al_u4780"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add64/ucin_al_u4780  (
    .a({\u2_Display/n1993 ,1'b1}),
    .b({\u2_Display/n1992 ,\u2_Display/n1994 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n1997 [1],open_n18258}),
    .fco(\u2_Display/add64/c3 ),
    .fx({\u2_Display/n1997 [2],\u2_Display/n1997 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u11_al_u4792  (
    .a({\u2_Display/n2016 ,\u2_Display/n2018 }),
    .b({\u2_Display/n2015 ,\u2_Display/n2017 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add65/c11 ),
    .f({\u2_Display/n2032 [13],\u2_Display/n2032 [11]}),
    .fco(\u2_Display/add65/c15 ),
    .fx({\u2_Display/n2032 [14],\u2_Display/n2032 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u15_al_u4793  (
    .a({\u2_Display/n2012 ,\u2_Display/n2014 }),
    .b({\u2_Display/n2011 ,\u2_Display/n2013 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add65/c15 ),
    .f({\u2_Display/n2032 [17],\u2_Display/n2032 [15]}),
    .fco(\u2_Display/add65/c19 ),
    .fx({\u2_Display/n2032 [18],\u2_Display/n2032 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u19_al_u4794  (
    .a({\u2_Display/n2008 ,\u2_Display/n2010 }),
    .b({\u2_Display/n2007 ,\u2_Display/n2009 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add65/c19 ),
    .f({\u2_Display/n2032 [21],\u2_Display/n2032 [19]}),
    .fco(\u2_Display/add65/c23 ),
    .fx({\u2_Display/n2032 [22],\u2_Display/n2032 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u23_al_u4795  (
    .a({\u2_Display/n2004 ,\u2_Display/n2006 }),
    .b({\u2_Display/n2003 ,\u2_Display/n2005 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add65/c23 ),
    .f({\u2_Display/n2032 [25],\u2_Display/n2032 [23]}),
    .fco(\u2_Display/add65/c27 ),
    .fx({\u2_Display/n2032 [26],\u2_Display/n2032 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u27_al_u4796  (
    .a({\u2_Display/n2000 ,\u2_Display/n2002 }),
    .b({\u2_Display/n1999 ,\u2_Display/n2001 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add65/c27 ),
    .f({\u2_Display/n2032 [29],\u2_Display/n2032 [27]}),
    .fco(\u2_Display/add65/c31 ),
    .fx({\u2_Display/n2032 [30],\u2_Display/n2032 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u31_al_u4797  (
    .a({open_n18351,\u2_Display/n1998 }),
    .c(2'b00),
    .d({open_n18356,1'b1}),
    .fci(\u2_Display/add65/c31 ),
    .f({open_n18373,\u2_Display/n2032 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u3_al_u4790  (
    .a({\u2_Display/n2024 ,\u2_Display/n2026 }),
    .b({\u2_Display/n2023 ,\u2_Display/n2025 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add65/c3 ),
    .f({\u2_Display/n2032 [5],\u2_Display/n2032 [3]}),
    .fco(\u2_Display/add65/c7 ),
    .fx({\u2_Display/n2032 [6],\u2_Display/n2032 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/u7_al_u4791  (
    .a({\u2_Display/n2020 ,\u2_Display/n2022 }),
    .b({\u2_Display/n2019 ,\u2_Display/n2021 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add65/c7 ),
    .f({\u2_Display/n2032 [9],\u2_Display/n2032 [7]}),
    .fco(\u2_Display/add65/c11 ),
    .fx({\u2_Display/n2032 [10],\u2_Display/n2032 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add65/ucin_al_u4789"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add65/ucin_al_u4789  (
    .a({\u2_Display/n2028 ,1'b1}),
    .b({\u2_Display/n2027 ,\u2_Display/n2029 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2032 [1],open_n18432}),
    .fco(\u2_Display/add65/c3 ),
    .fx({\u2_Display/n2032 [2],\u2_Display/n2032 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u11_al_u4801  (
    .a({\u2_Display/n2051 ,\u2_Display/n2053 }),
    .b({\u2_Display/n2050 ,\u2_Display/n2052 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add66/c11 ),
    .f({\u2_Display/n2067 [13],\u2_Display/n2067 [11]}),
    .fco(\u2_Display/add66/c15 ),
    .fx({\u2_Display/n2067 [14],\u2_Display/n2067 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u15_al_u4802  (
    .a({\u2_Display/n2047 ,\u2_Display/n2049 }),
    .b({\u2_Display/n2046 ,\u2_Display/n2048 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add66/c15 ),
    .f({\u2_Display/n2067 [17],\u2_Display/n2067 [15]}),
    .fco(\u2_Display/add66/c19 ),
    .fx({\u2_Display/n2067 [18],\u2_Display/n2067 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u19_al_u4803  (
    .a({\u2_Display/n2043 ,\u2_Display/n2045 }),
    .b({\u2_Display/n2042 ,\u2_Display/n2044 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add66/c19 ),
    .f({\u2_Display/n2067 [21],\u2_Display/n2067 [19]}),
    .fco(\u2_Display/add66/c23 ),
    .fx({\u2_Display/n2067 [22],\u2_Display/n2067 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u23_al_u4804  (
    .a({\u2_Display/n2039 ,\u2_Display/n2041 }),
    .b({\u2_Display/n2038 ,\u2_Display/n2040 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add66/c23 ),
    .f({\u2_Display/n2067 [25],\u2_Display/n2067 [23]}),
    .fco(\u2_Display/add66/c27 ),
    .fx({\u2_Display/n2067 [26],\u2_Display/n2067 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u27_al_u4805  (
    .a({\u2_Display/n2035 ,\u2_Display/n2037 }),
    .b({\u2_Display/n2034 ,\u2_Display/n2036 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add66/c27 ),
    .f({\u2_Display/n2067 [29],\u2_Display/n2067 [27]}),
    .fco(\u2_Display/add66/c31 ),
    .fx({\u2_Display/n2067 [30],\u2_Display/n2067 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u31_al_u4806  (
    .a({open_n18525,\u2_Display/n2033 }),
    .c(2'b00),
    .d({open_n18530,1'b1}),
    .fci(\u2_Display/add66/c31 ),
    .f({open_n18547,\u2_Display/n2067 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u3_al_u4799  (
    .a({\u2_Display/n2059 ,\u2_Display/n2061 }),
    .b({\u2_Display/n2058 ,\u2_Display/n2060 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add66/c3 ),
    .f({\u2_Display/n2067 [5],\u2_Display/n2067 [3]}),
    .fco(\u2_Display/add66/c7 ),
    .fx({\u2_Display/n2067 [6],\u2_Display/n2067 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/u7_al_u4800  (
    .a({\u2_Display/n2055 ,\u2_Display/n2057 }),
    .b({\u2_Display/n2054 ,\u2_Display/n2056 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add66/c7 ),
    .f({\u2_Display/n2067 [9],\u2_Display/n2067 [7]}),
    .fco(\u2_Display/add66/c11 ),
    .fx({\u2_Display/n2067 [10],\u2_Display/n2067 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add66/ucin_al_u4798"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add66/ucin_al_u4798  (
    .a({\u2_Display/n2063 ,1'b1}),
    .b({\u2_Display/n2062 ,\u2_Display/n2064 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2067 [1],open_n18606}),
    .fco(\u2_Display/add66/c3 ),
    .fx({\u2_Display/n2067 [2],\u2_Display/n2067 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u11_al_u4810  (
    .a({\u2_Display/n2086 ,\u2_Display/n2088 }),
    .b({\u2_Display/n2085 ,\u2_Display/n2087 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add67/c11 ),
    .f({\u2_Display/n2102 [13],\u2_Display/n2102 [11]}),
    .fco(\u2_Display/add67/c15 ),
    .fx({\u2_Display/n2102 [14],\u2_Display/n2102 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u15_al_u4811  (
    .a({\u2_Display/n2082 ,\u2_Display/n2084 }),
    .b({\u2_Display/n2081 ,\u2_Display/n2083 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add67/c15 ),
    .f({\u2_Display/n2102 [17],\u2_Display/n2102 [15]}),
    .fco(\u2_Display/add67/c19 ),
    .fx({\u2_Display/n2102 [18],\u2_Display/n2102 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u19_al_u4812  (
    .a({\u2_Display/n2078 ,\u2_Display/n2080 }),
    .b({\u2_Display/n2077 ,\u2_Display/n2079 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add67/c19 ),
    .f({\u2_Display/n2102 [21],\u2_Display/n2102 [19]}),
    .fco(\u2_Display/add67/c23 ),
    .fx({\u2_Display/n2102 [22],\u2_Display/n2102 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u23_al_u4813  (
    .a({\u2_Display/n2074 ,\u2_Display/n2076 }),
    .b({\u2_Display/n2073 ,\u2_Display/n2075 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add67/c23 ),
    .f({\u2_Display/n2102 [25],\u2_Display/n2102 [23]}),
    .fco(\u2_Display/add67/c27 ),
    .fx({\u2_Display/n2102 [26],\u2_Display/n2102 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u27_al_u4814  (
    .a({\u2_Display/n2070 ,\u2_Display/n2072 }),
    .b({\u2_Display/n2069 ,\u2_Display/n2071 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add67/c27 ),
    .f({\u2_Display/n2102 [29],\u2_Display/n2102 [27]}),
    .fco(\u2_Display/add67/c31 ),
    .fx({\u2_Display/n2102 [30],\u2_Display/n2102 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u31_al_u4815  (
    .a({open_n18699,\u2_Display/n2068 }),
    .c(2'b00),
    .d({open_n18704,1'b1}),
    .fci(\u2_Display/add67/c31 ),
    .f({open_n18721,\u2_Display/n2102 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u3_al_u4808  (
    .a({\u2_Display/n2094 ,\u2_Display/n2096 }),
    .b({\u2_Display/n2093 ,\u2_Display/n2095 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add67/c3 ),
    .f({\u2_Display/n2102 [5],\u2_Display/n2102 [3]}),
    .fco(\u2_Display/add67/c7 ),
    .fx({\u2_Display/n2102 [6],\u2_Display/n2102 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/u7_al_u4809  (
    .a({\u2_Display/n2090 ,\u2_Display/n2092 }),
    .b({\u2_Display/n2089 ,\u2_Display/n2091 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add67/c7 ),
    .f({\u2_Display/n2102 [9],\u2_Display/n2102 [7]}),
    .fco(\u2_Display/add67/c11 ),
    .fx({\u2_Display/n2102 [10],\u2_Display/n2102 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add67/ucin_al_u4807"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add67/ucin_al_u4807  (
    .a({\u2_Display/n2098 ,1'b1}),
    .b({\u2_Display/n2097 ,\u2_Display/n2099 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2102 [1],open_n18780}),
    .fco(\u2_Display/add67/c3 ),
    .fx({\u2_Display/n2102 [2],\u2_Display/n2102 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u11_al_u4819  (
    .a({\u2_Display/n2121 ,\u2_Display/n2123 }),
    .b({\u2_Display/n2120 ,\u2_Display/n2122 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add68/c11 ),
    .f({\u2_Display/n2137 [13],\u2_Display/n2137 [11]}),
    .fco(\u2_Display/add68/c15 ),
    .fx({\u2_Display/n2137 [14],\u2_Display/n2137 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u15_al_u4820  (
    .a({\u2_Display/n2117 ,\u2_Display/n2119 }),
    .b({\u2_Display/n2116 ,\u2_Display/n2118 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add68/c15 ),
    .f({\u2_Display/n2137 [17],\u2_Display/n2137 [15]}),
    .fco(\u2_Display/add68/c19 ),
    .fx({\u2_Display/n2137 [18],\u2_Display/n2137 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u19_al_u4821  (
    .a({\u2_Display/n2113 ,\u2_Display/n2115 }),
    .b({\u2_Display/n2112 ,\u2_Display/n2114 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add68/c19 ),
    .f({\u2_Display/n2137 [21],\u2_Display/n2137 [19]}),
    .fco(\u2_Display/add68/c23 ),
    .fx({\u2_Display/n2137 [22],\u2_Display/n2137 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u23_al_u4822  (
    .a({\u2_Display/n2109 ,\u2_Display/n2111 }),
    .b({\u2_Display/n2108 ,\u2_Display/n2110 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add68/c23 ),
    .f({\u2_Display/n2137 [25],\u2_Display/n2137 [23]}),
    .fco(\u2_Display/add68/c27 ),
    .fx({\u2_Display/n2137 [26],\u2_Display/n2137 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u27_al_u4823  (
    .a({\u2_Display/n2105 ,\u2_Display/n2107 }),
    .b({\u2_Display/n2104 ,\u2_Display/n2106 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add68/c27 ),
    .f({\u2_Display/n2137 [29],\u2_Display/n2137 [27]}),
    .fco(\u2_Display/add68/c31 ),
    .fx({\u2_Display/n2137 [30],\u2_Display/n2137 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u31_al_u4824  (
    .a({open_n18873,\u2_Display/n2103 }),
    .c(2'b00),
    .d({open_n18878,1'b1}),
    .fci(\u2_Display/add68/c31 ),
    .f({open_n18895,\u2_Display/n2137 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u3_al_u4817  (
    .a({\u2_Display/n2129 ,\u2_Display/n2131 }),
    .b({\u2_Display/n2128 ,\u2_Display/n2130 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add68/c3 ),
    .f({\u2_Display/n2137 [5],\u2_Display/n2137 [3]}),
    .fco(\u2_Display/add68/c7 ),
    .fx({\u2_Display/n2137 [6],\u2_Display/n2137 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/u7_al_u4818  (
    .a({\u2_Display/n2125 ,\u2_Display/n2127 }),
    .b({\u2_Display/n2124 ,\u2_Display/n2126 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add68/c7 ),
    .f({\u2_Display/n2137 [9],\u2_Display/n2137 [7]}),
    .fco(\u2_Display/add68/c11 ),
    .fx({\u2_Display/n2137 [10],\u2_Display/n2137 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add68/ucin_al_u4816"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add68/ucin_al_u4816  (
    .a({\u2_Display/n2133 ,1'b1}),
    .b({\u2_Display/n2132 ,\u2_Display/n2134 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2137 [1],open_n18954}),
    .fco(\u2_Display/add68/c3 ),
    .fx({\u2_Display/n2137 [2],\u2_Display/n2137 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u11_al_u4828  (
    .a({\u2_Display/n2156 ,\u2_Display/n2158 }),
    .b({\u2_Display/n2155 ,\u2_Display/n2157 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b10),
    .fci(\u2_Display/add69/c11 ),
    .f({\u2_Display/n2172 [13],\u2_Display/n2172 [11]}),
    .fco(\u2_Display/add69/c15 ),
    .fx({\u2_Display/n2172 [14],\u2_Display/n2172 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u15_al_u4829  (
    .a({\u2_Display/n2152 ,\u2_Display/n2154 }),
    .b({\u2_Display/n2151 ,\u2_Display/n2153 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add69/c15 ),
    .f({\u2_Display/n2172 [17],\u2_Display/n2172 [15]}),
    .fco(\u2_Display/add69/c19 ),
    .fx({\u2_Display/n2172 [18],\u2_Display/n2172 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u19_al_u4830  (
    .a({\u2_Display/n2148 ,\u2_Display/n2150 }),
    .b({\u2_Display/n2147 ,\u2_Display/n2149 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add69/c19 ),
    .f({\u2_Display/n2172 [21],\u2_Display/n2172 [19]}),
    .fco(\u2_Display/add69/c23 ),
    .fx({\u2_Display/n2172 [22],\u2_Display/n2172 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u23_al_u4831  (
    .a({\u2_Display/n2144 ,\u2_Display/n2146 }),
    .b({\u2_Display/n2143 ,\u2_Display/n2145 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add69/c23 ),
    .f({\u2_Display/n2172 [25],\u2_Display/n2172 [23]}),
    .fco(\u2_Display/add69/c27 ),
    .fx({\u2_Display/n2172 [26],\u2_Display/n2172 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u27_al_u4832  (
    .a({\u2_Display/n2140 ,\u2_Display/n2142 }),
    .b({\u2_Display/n2139 ,\u2_Display/n2141 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add69/c27 ),
    .f({\u2_Display/n2172 [29],\u2_Display/n2172 [27]}),
    .fco(\u2_Display/add69/c31 ),
    .fx({\u2_Display/n2172 [30],\u2_Display/n2172 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u31_al_u4833  (
    .a({open_n19047,\u2_Display/n2138 }),
    .c(2'b00),
    .d({open_n19052,1'b1}),
    .fci(\u2_Display/add69/c31 ),
    .f({open_n19069,\u2_Display/n2172 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u3_al_u4826  (
    .a({\u2_Display/n2164 ,\u2_Display/n2166 }),
    .b({\u2_Display/n2163 ,\u2_Display/n2165 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add69/c3 ),
    .f({\u2_Display/n2172 [5],\u2_Display/n2172 [3]}),
    .fco(\u2_Display/add69/c7 ),
    .fx({\u2_Display/n2172 [6],\u2_Display/n2172 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/u7_al_u4827  (
    .a({\u2_Display/n2160 ,\u2_Display/n2162 }),
    .b({\u2_Display/n2159 ,\u2_Display/n2161 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add69/c7 ),
    .f({\u2_Display/n2172 [9],\u2_Display/n2172 [7]}),
    .fco(\u2_Display/add69/c11 ),
    .fx({\u2_Display/n2172 [10],\u2_Display/n2172 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add69/ucin_al_u4825"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add69/ucin_al_u4825  (
    .a({\u2_Display/n2168 ,1'b1}),
    .b({\u2_Display/n2167 ,\u2_Display/n2169 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2172 [1],open_n19128}),
    .fco(\u2_Display/add69/c3 ),
    .fx({\u2_Display/n2172 [2],\u2_Display/n2172 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add6_2/u0|u2_Display/add6_2/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add6_2/u0|u2_Display/add6_2/ucin  (
    .a(2'b10),
    .b({\u2_Display/j [7],open_n19131}),
    .f({\u2_Display/n135 [0],open_n19151}),
    .fco(\u2_Display/add6_2/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add6_2/u0|u2_Display/add6_2/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add6_2/u2|u2_Display/add6_2/u1  (
    .a(2'b10),
    .b(\u2_Display/j [9:8]),
    .fci(\u2_Display/add6_2/c1 ),
    .f(\u2_Display/n135 [2:1]),
    .fco(\u2_Display/add6_2/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/add6_2/u0|u2_Display/add6_2/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u2_Display/add6_2/ucout_al_u5059  (
    .fci(\u2_Display/add6_2/c3 ),
    .f({open_n19200,\u2_Display/add6_2_co }));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u11_al_u4837  (
    .a({\u2_Display/n2191 ,\u2_Display/n2193 }),
    .b({\u2_Display/n2190 ,\u2_Display/n2192 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b10),
    .fci(\u2_Display/add70/c11 ),
    .f({\u2_Display/n2207 [13],\u2_Display/n2207 [11]}),
    .fco(\u2_Display/add70/c15 ),
    .fx({\u2_Display/n2207 [14],\u2_Display/n2207 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u15_al_u4838  (
    .a({\u2_Display/n2187 ,\u2_Display/n2189 }),
    .b({\u2_Display/n2186 ,\u2_Display/n2188 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add70/c15 ),
    .f({\u2_Display/n2207 [17],\u2_Display/n2207 [15]}),
    .fco(\u2_Display/add70/c19 ),
    .fx({\u2_Display/n2207 [18],\u2_Display/n2207 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u19_al_u4839  (
    .a({\u2_Display/n2183 ,\u2_Display/n2185 }),
    .b({\u2_Display/n2182 ,\u2_Display/n2184 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add70/c19 ),
    .f({\u2_Display/n2207 [21],\u2_Display/n2207 [19]}),
    .fco(\u2_Display/add70/c23 ),
    .fx({\u2_Display/n2207 [22],\u2_Display/n2207 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u23_al_u4840  (
    .a({\u2_Display/n2179 ,\u2_Display/n2181 }),
    .b({\u2_Display/n2178 ,\u2_Display/n2180 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add70/c23 ),
    .f({\u2_Display/n2207 [25],\u2_Display/n2207 [23]}),
    .fco(\u2_Display/add70/c27 ),
    .fx({\u2_Display/n2207 [26],\u2_Display/n2207 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u27_al_u4841  (
    .a({\u2_Display/n2175 ,\u2_Display/n2177 }),
    .b({\u2_Display/n2174 ,\u2_Display/n2176 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add70/c27 ),
    .f({\u2_Display/n2207 [29],\u2_Display/n2207 [27]}),
    .fco(\u2_Display/add70/c31 ),
    .fx({\u2_Display/n2207 [30],\u2_Display/n2207 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u31_al_u4842  (
    .a({open_n19296,\u2_Display/n2173 }),
    .c(2'b00),
    .d({open_n19301,1'b1}),
    .fci(\u2_Display/add70/c31 ),
    .f({open_n19318,\u2_Display/n2207 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u3_al_u4835  (
    .a({\u2_Display/n2199 ,\u2_Display/n2201 }),
    .b({\u2_Display/n2198 ,\u2_Display/n2200 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add70/c3 ),
    .f({\u2_Display/n2207 [5],\u2_Display/n2207 [3]}),
    .fco(\u2_Display/add70/c7 ),
    .fx({\u2_Display/n2207 [6],\u2_Display/n2207 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/u7_al_u4836  (
    .a({\u2_Display/n2195 ,\u2_Display/n2197 }),
    .b({\u2_Display/n2194 ,\u2_Display/n2196 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add70/c7 ),
    .f({\u2_Display/n2207 [9],\u2_Display/n2207 [7]}),
    .fco(\u2_Display/add70/c11 ),
    .fx({\u2_Display/n2207 [10],\u2_Display/n2207 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add70/ucin_al_u4834"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add70/ucin_al_u4834  (
    .a({\u2_Display/n2203 ,1'b1}),
    .b({\u2_Display/n2202 ,\u2_Display/n2204 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2207 [1],open_n19377}),
    .fco(\u2_Display/add70/c3 ),
    .fx({\u2_Display/n2207 [2],\u2_Display/n2207 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u11_al_u4846  (
    .a({\u2_Display/n2226 ,\u2_Display/n2228 }),
    .b({\u2_Display/n2225 ,\u2_Display/n2227 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add71/c11 ),
    .f({\u2_Display/n2242 [13],\u2_Display/n2242 [11]}),
    .fco(\u2_Display/add71/c15 ),
    .fx({\u2_Display/n2242 [14],\u2_Display/n2242 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u15_al_u4847  (
    .a({\u2_Display/n2222 ,\u2_Display/n2224 }),
    .b({\u2_Display/n2221 ,\u2_Display/n2223 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add71/c15 ),
    .f({\u2_Display/n2242 [17],\u2_Display/n2242 [15]}),
    .fco(\u2_Display/add71/c19 ),
    .fx({\u2_Display/n2242 [18],\u2_Display/n2242 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u19_al_u4848  (
    .a({\u2_Display/n2218 ,\u2_Display/n2220 }),
    .b({\u2_Display/n2217 ,\u2_Display/n2219 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add71/c19 ),
    .f({\u2_Display/n2242 [21],\u2_Display/n2242 [19]}),
    .fco(\u2_Display/add71/c23 ),
    .fx({\u2_Display/n2242 [22],\u2_Display/n2242 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u23_al_u4849  (
    .a({\u2_Display/n2214 ,\u2_Display/n2216 }),
    .b({\u2_Display/n2213 ,\u2_Display/n2215 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add71/c23 ),
    .f({\u2_Display/n2242 [25],\u2_Display/n2242 [23]}),
    .fco(\u2_Display/add71/c27 ),
    .fx({\u2_Display/n2242 [26],\u2_Display/n2242 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u27_al_u4850  (
    .a({\u2_Display/n2210 ,\u2_Display/n2212 }),
    .b({\u2_Display/n2209 ,\u2_Display/n2211 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add71/c27 ),
    .f({\u2_Display/n2242 [29],\u2_Display/n2242 [27]}),
    .fco(\u2_Display/add71/c31 ),
    .fx({\u2_Display/n2242 [30],\u2_Display/n2242 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u31_al_u4851  (
    .a({open_n19470,\u2_Display/n2208 }),
    .c(2'b00),
    .d({open_n19475,1'b1}),
    .fci(\u2_Display/add71/c31 ),
    .f({open_n19492,\u2_Display/n2242 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u3_al_u4844  (
    .a({\u2_Display/n2234 ,\u2_Display/n2236 }),
    .b({\u2_Display/n2233 ,\u2_Display/n2235 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add71/c3 ),
    .f({\u2_Display/n2242 [5],\u2_Display/n2242 [3]}),
    .fco(\u2_Display/add71/c7 ),
    .fx({\u2_Display/n2242 [6],\u2_Display/n2242 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/u7_al_u4845  (
    .a({\u2_Display/n2230 ,\u2_Display/n2232 }),
    .b({\u2_Display/n2229 ,\u2_Display/n2231 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add71/c7 ),
    .f({\u2_Display/n2242 [9],\u2_Display/n2242 [7]}),
    .fco(\u2_Display/add71/c11 ),
    .fx({\u2_Display/n2242 [10],\u2_Display/n2242 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add71/ucin_al_u4843"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add71/ucin_al_u4843  (
    .a({\u2_Display/n2238 ,1'b1}),
    .b({\u2_Display/n2237 ,\u2_Display/n2239 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2242 [1],open_n19551}),
    .fco(\u2_Display/add71/c3 ),
    .fx({\u2_Display/n2242 [2],\u2_Display/n2242 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u11_al_u4855  (
    .a({\u2_Display/n2261 ,\u2_Display/n2263 }),
    .b({\u2_Display/n2260 ,\u2_Display/n2262 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add72/c11 ),
    .f({\u2_Display/n2277 [13],\u2_Display/n2277 [11]}),
    .fco(\u2_Display/add72/c15 ),
    .fx({\u2_Display/n2277 [14],\u2_Display/n2277 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u15_al_u4856  (
    .a({\u2_Display/n2257 ,\u2_Display/n2259 }),
    .b({\u2_Display/n2256 ,\u2_Display/n2258 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add72/c15 ),
    .f({\u2_Display/n2277 [17],\u2_Display/n2277 [15]}),
    .fco(\u2_Display/add72/c19 ),
    .fx({\u2_Display/n2277 [18],\u2_Display/n2277 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u19_al_u4857  (
    .a({\u2_Display/n2253 ,\u2_Display/n2255 }),
    .b({\u2_Display/n2252 ,\u2_Display/n2254 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add72/c19 ),
    .f({\u2_Display/n2277 [21],\u2_Display/n2277 [19]}),
    .fco(\u2_Display/add72/c23 ),
    .fx({\u2_Display/n2277 [22],\u2_Display/n2277 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u23_al_u4858  (
    .a({\u2_Display/n2249 ,\u2_Display/n2251 }),
    .b({\u2_Display/n2248 ,\u2_Display/n2250 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add72/c23 ),
    .f({\u2_Display/n2277 [25],\u2_Display/n2277 [23]}),
    .fco(\u2_Display/add72/c27 ),
    .fx({\u2_Display/n2277 [26],\u2_Display/n2277 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u27_al_u4859  (
    .a({\u2_Display/n2245 ,\u2_Display/n2247 }),
    .b({\u2_Display/n2244 ,\u2_Display/n2246 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add72/c27 ),
    .f({\u2_Display/n2277 [29],\u2_Display/n2277 [27]}),
    .fco(\u2_Display/add72/c31 ),
    .fx({\u2_Display/n2277 [30],\u2_Display/n2277 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u31_al_u4860  (
    .a({open_n19644,\u2_Display/n2243 }),
    .c(2'b00),
    .d({open_n19649,1'b1}),
    .fci(\u2_Display/add72/c31 ),
    .f({open_n19666,\u2_Display/n2277 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u3_al_u4853  (
    .a({\u2_Display/n2269 ,\u2_Display/n2271 }),
    .b({\u2_Display/n2268 ,\u2_Display/n2270 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add72/c3 ),
    .f({\u2_Display/n2277 [5],\u2_Display/n2277 [3]}),
    .fco(\u2_Display/add72/c7 ),
    .fx({\u2_Display/n2277 [6],\u2_Display/n2277 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/u7_al_u4854  (
    .a({\u2_Display/n2265 ,\u2_Display/n2267 }),
    .b({\u2_Display/n2264 ,\u2_Display/n2266 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b00),
    .fci(\u2_Display/add72/c7 ),
    .f({\u2_Display/n2277 [9],\u2_Display/n2277 [7]}),
    .fco(\u2_Display/add72/c11 ),
    .fx({\u2_Display/n2277 [10],\u2_Display/n2277 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add72/ucin_al_u4852"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add72/ucin_al_u4852  (
    .a({\u2_Display/n2273 ,1'b1}),
    .b({\u2_Display/n2272 ,\u2_Display/n2274 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2277 [1],open_n19725}),
    .fco(\u2_Display/add72/c3 ),
    .fx({\u2_Display/n2277 [2],\u2_Display/n2277 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add73/ucin_al_u5055"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add73/u3_al_u5056  (
    .a({\u2_Display/n2304 ,\u2_Display/n2306 }),
    .b({\u2_Display/n2303 ,\u2_Display/n2305 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add73/c3 ),
    .f({\u2_Display/n2312 [5],\u2_Display/n2312 [3]}),
    .fco(\u2_Display/add73/c7 ),
    .fx({\u2_Display/n2312 [6],\u2_Display/n2312 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add73/ucin_al_u5055"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add73/u7_al_u5057  (
    .a({\u2_Display/n2300 ,\u2_Display/n2302 }),
    .b({open_n19746,\u2_Display/n2301 }),
    .c(2'b00),
    .d(2'b00),
    .e({open_n19749,1'b0}),
    .fci(\u2_Display/add73/c7 ),
    .f({\u2_Display/n2312 [9],\u2_Display/n2312 [7]}),
    .fx({open_n19765,\u2_Display/n2312 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add73/ucin_al_u5055"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add73/ucin_al_u5055  (
    .a({\u2_Display/n2308 ,1'b1}),
    .b({\u2_Display/n2307 ,\u2_Display/n2309 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .f({\u2_Display/n2312 [1],open_n19785}),
    .fco(\u2_Display/add73/c3 ),
    .fx({\u2_Display/n2312 [2],\u2_Display/n2312 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u11_al_u4864  (
    .a({\u2_Display/counta [13],\u2_Display/counta [11]}),
    .b({\u2_Display/counta [14],\u2_Display/counta [12]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add84/c11 ),
    .f({\u2_Display/n2665 [13],\u2_Display/n2665 [11]}),
    .fco(\u2_Display/add84/c15 ),
    .fx({\u2_Display/n2665 [14],\u2_Display/n2665 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u15_al_u4865  (
    .a({\u2_Display/counta [17],\u2_Display/counta [15]}),
    .b({\u2_Display/counta [18],\u2_Display/counta [16]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add84/c15 ),
    .f({\u2_Display/n2665 [17],\u2_Display/n2665 [15]}),
    .fco(\u2_Display/add84/c19 ),
    .fx({\u2_Display/n2665 [18],\u2_Display/n2665 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u19_al_u4866  (
    .a({\u2_Display/counta [21],\u2_Display/counta [19]}),
    .b({\u2_Display/counta [22],\u2_Display/counta [20]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add84/c19 ),
    .f({\u2_Display/n2665 [21],\u2_Display/n2665 [19]}),
    .fco(\u2_Display/add84/c23 ),
    .fx({\u2_Display/n2665 [22],\u2_Display/n2665 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u23_al_u4867  (
    .a({\u2_Display/counta [25],\u2_Display/counta [23]}),
    .b({\u2_Display/counta [26],\u2_Display/counta [24]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add84/c23 ),
    .f({\u2_Display/n2665 [25],\u2_Display/n2665 [23]}),
    .fco(\u2_Display/add84/c27 ),
    .fx({\u2_Display/n2665 [26],\u2_Display/n2665 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u27_al_u4868  (
    .a({\u2_Display/counta [29],\u2_Display/counta [27]}),
    .b({\u2_Display/counta [30],\u2_Display/counta [28]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add84/c27 ),
    .f({\u2_Display/n2665 [29],\u2_Display/n2665 [27]}),
    .fco(\u2_Display/add84/c31 ),
    .fx({\u2_Display/n2665 [30],\u2_Display/n2665 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u31_al_u4869  (
    .a({open_n19878,\u2_Display/counta [31]}),
    .c(2'b00),
    .d({open_n19883,1'b0}),
    .fci(\u2_Display/add84/c31 ),
    .f({open_n19900,\u2_Display/n2665 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u3_al_u4862  (
    .a({\u2_Display/counta [5],\u2_Display/counta [3]}),
    .b({\u2_Display/counta [6],\u2_Display/counta [4]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add84/c3 ),
    .f({\u2_Display/n2665 [5],\u2_Display/n2665 [3]}),
    .fco(\u2_Display/add84/c7 ),
    .fx({\u2_Display/n2665 [6],\u2_Display/n2665 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/u7_al_u4863  (
    .a({\u2_Display/counta [9],\u2_Display/counta [7]}),
    .b({\u2_Display/counta [10],\u2_Display/counta [8]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add84/c7 ),
    .f({\u2_Display/n2665 [9],\u2_Display/n2665 [7]}),
    .fco(\u2_Display/add84/c11 ),
    .fx({\u2_Display/n2665 [10],\u2_Display/n2665 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add84/ucin_al_u4861"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add84/ucin_al_u4861  (
    .a({\u2_Display/counta [1],1'b1}),
    .b({\u2_Display/counta [2],\u2_Display/counta [0]}),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2665 [1],open_n19959}),
    .fco(\u2_Display/add84/c3 ),
    .fx({\u2_Display/n2665 [2],\u2_Display/n2665 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u11_al_u4873  (
    .a({\u2_Display/n2684 ,\u2_Display/n2686 }),
    .b({\u2_Display/n2683 ,\u2_Display/n2685 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add85/c11 ),
    .f({\u2_Display/n2700 [13],\u2_Display/n2700 [11]}),
    .fco(\u2_Display/add85/c15 ),
    .fx({\u2_Display/n2700 [14],\u2_Display/n2700 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u15_al_u4874  (
    .a({\u2_Display/n2680 ,\u2_Display/n2682 }),
    .b({\u2_Display/n2679 ,\u2_Display/n2681 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add85/c15 ),
    .f({\u2_Display/n2700 [17],\u2_Display/n2700 [15]}),
    .fco(\u2_Display/add85/c19 ),
    .fx({\u2_Display/n2700 [18],\u2_Display/n2700 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u19_al_u4875  (
    .a({\u2_Display/n2676 ,\u2_Display/n2678 }),
    .b({\u2_Display/n2675 ,\u2_Display/n2677 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add85/c19 ),
    .f({\u2_Display/n2700 [21],\u2_Display/n2700 [19]}),
    .fco(\u2_Display/add85/c23 ),
    .fx({\u2_Display/n2700 [22],\u2_Display/n2700 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u23_al_u4876  (
    .a({\u2_Display/n2672 ,\u2_Display/n2674 }),
    .b({\u2_Display/n2671 ,\u2_Display/n2673 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add85/c23 ),
    .f({\u2_Display/n2700 [25],\u2_Display/n2700 [23]}),
    .fco(\u2_Display/add85/c27 ),
    .fx({\u2_Display/n2700 [26],\u2_Display/n2700 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u27_al_u4877  (
    .a({\u2_Display/n2668 ,\u2_Display/n2670 }),
    .b({\u2_Display/n2667 ,\u2_Display/n2669 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add85/c27 ),
    .f({\u2_Display/n2700 [29],\u2_Display/n2700 [27]}),
    .fco(\u2_Display/add85/c31 ),
    .fx({\u2_Display/n2700 [30],\u2_Display/n2700 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u31_al_u4878  (
    .a({open_n20052,\u2_Display/n2666 }),
    .c(2'b00),
    .d({open_n20057,1'b1}),
    .fci(\u2_Display/add85/c31 ),
    .f({open_n20074,\u2_Display/n2700 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u3_al_u4871  (
    .a({\u2_Display/n2692 ,\u2_Display/n2694 }),
    .b({\u2_Display/n2691 ,\u2_Display/n2693 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add85/c3 ),
    .f({\u2_Display/n2700 [5],\u2_Display/n2700 [3]}),
    .fco(\u2_Display/add85/c7 ),
    .fx({\u2_Display/n2700 [6],\u2_Display/n2700 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/u7_al_u4872  (
    .a({\u2_Display/n2688 ,\u2_Display/n2690 }),
    .b({\u2_Display/n2687 ,\u2_Display/n2689 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add85/c7 ),
    .f({\u2_Display/n2700 [9],\u2_Display/n2700 [7]}),
    .fco(\u2_Display/add85/c11 ),
    .fx({\u2_Display/n2700 [10],\u2_Display/n2700 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add85/ucin_al_u4870"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add85/ucin_al_u4870  (
    .a({\u2_Display/n2696 ,1'b1}),
    .b({\u2_Display/n2695 ,\u2_Display/n2697 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2700 [1],open_n20133}),
    .fco(\u2_Display/add85/c3 ),
    .fx({\u2_Display/n2700 [2],\u2_Display/n2700 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u11_al_u4882  (
    .a({\u2_Display/n2719 ,\u2_Display/n2721 }),
    .b({\u2_Display/n2718 ,\u2_Display/n2720 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add86/c11 ),
    .f({\u2_Display/n2735 [13],\u2_Display/n2735 [11]}),
    .fco(\u2_Display/add86/c15 ),
    .fx({\u2_Display/n2735 [14],\u2_Display/n2735 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u15_al_u4883  (
    .a({\u2_Display/n2715 ,\u2_Display/n2717 }),
    .b({\u2_Display/n2714 ,\u2_Display/n2716 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add86/c15 ),
    .f({\u2_Display/n2735 [17],\u2_Display/n2735 [15]}),
    .fco(\u2_Display/add86/c19 ),
    .fx({\u2_Display/n2735 [18],\u2_Display/n2735 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u19_al_u4884  (
    .a({\u2_Display/n2711 ,\u2_Display/n2713 }),
    .b({\u2_Display/n2710 ,\u2_Display/n2712 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add86/c19 ),
    .f({\u2_Display/n2735 [21],\u2_Display/n2735 [19]}),
    .fco(\u2_Display/add86/c23 ),
    .fx({\u2_Display/n2735 [22],\u2_Display/n2735 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u23_al_u4885  (
    .a({\u2_Display/n2707 ,\u2_Display/n2709 }),
    .b({\u2_Display/n2706 ,\u2_Display/n2708 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b00),
    .fci(\u2_Display/add86/c23 ),
    .f({\u2_Display/n2735 [25],\u2_Display/n2735 [23]}),
    .fco(\u2_Display/add86/c27 ),
    .fx({\u2_Display/n2735 [26],\u2_Display/n2735 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u27_al_u4886  (
    .a({\u2_Display/n2703 ,\u2_Display/n2705 }),
    .b({\u2_Display/n2702 ,\u2_Display/n2704 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add86/c27 ),
    .f({\u2_Display/n2735 [29],\u2_Display/n2735 [27]}),
    .fco(\u2_Display/add86/c31 ),
    .fx({\u2_Display/n2735 [30],\u2_Display/n2735 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u31_al_u4887  (
    .a({open_n20226,\u2_Display/n2701 }),
    .c(2'b00),
    .d({open_n20231,1'b1}),
    .fci(\u2_Display/add86/c31 ),
    .f({open_n20248,\u2_Display/n2735 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u3_al_u4880  (
    .a({\u2_Display/n2727 ,\u2_Display/n2729 }),
    .b({\u2_Display/n2726 ,\u2_Display/n2728 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add86/c3 ),
    .f({\u2_Display/n2735 [5],\u2_Display/n2735 [3]}),
    .fco(\u2_Display/add86/c7 ),
    .fx({\u2_Display/n2735 [6],\u2_Display/n2735 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/u7_al_u4881  (
    .a({\u2_Display/n2723 ,\u2_Display/n2725 }),
    .b({\u2_Display/n2722 ,\u2_Display/n2724 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add86/c7 ),
    .f({\u2_Display/n2735 [9],\u2_Display/n2735 [7]}),
    .fco(\u2_Display/add86/c11 ),
    .fx({\u2_Display/n2735 [10],\u2_Display/n2735 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add86/ucin_al_u4879"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add86/ucin_al_u4879  (
    .a({\u2_Display/n2731 ,1'b1}),
    .b({\u2_Display/n2730 ,\u2_Display/n2732 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2735 [1],open_n20307}),
    .fco(\u2_Display/add86/c3 ),
    .fx({\u2_Display/n2735 [2],\u2_Display/n2735 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u11_al_u4891  (
    .a({\u2_Display/n2754 ,\u2_Display/n2756 }),
    .b({\u2_Display/n2753 ,\u2_Display/n2755 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add87/c11 ),
    .f({\u2_Display/n2770 [13],\u2_Display/n2770 [11]}),
    .fco(\u2_Display/add87/c15 ),
    .fx({\u2_Display/n2770 [14],\u2_Display/n2770 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u15_al_u4892  (
    .a({\u2_Display/n2750 ,\u2_Display/n2752 }),
    .b({\u2_Display/n2749 ,\u2_Display/n2751 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add87/c15 ),
    .f({\u2_Display/n2770 [17],\u2_Display/n2770 [15]}),
    .fco(\u2_Display/add87/c19 ),
    .fx({\u2_Display/n2770 [18],\u2_Display/n2770 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u19_al_u4893  (
    .a({\u2_Display/n2746 ,\u2_Display/n2748 }),
    .b({\u2_Display/n2745 ,\u2_Display/n2747 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add87/c19 ),
    .f({\u2_Display/n2770 [21],\u2_Display/n2770 [19]}),
    .fco(\u2_Display/add87/c23 ),
    .fx({\u2_Display/n2770 [22],\u2_Display/n2770 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u23_al_u4894  (
    .a({\u2_Display/n2742 ,\u2_Display/n2744 }),
    .b({\u2_Display/n2741 ,\u2_Display/n2743 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add87/c23 ),
    .f({\u2_Display/n2770 [25],\u2_Display/n2770 [23]}),
    .fco(\u2_Display/add87/c27 ),
    .fx({\u2_Display/n2770 [26],\u2_Display/n2770 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u27_al_u4895  (
    .a({\u2_Display/n2738 ,\u2_Display/n2740 }),
    .b({\u2_Display/n2737 ,\u2_Display/n2739 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add87/c27 ),
    .f({\u2_Display/n2770 [29],\u2_Display/n2770 [27]}),
    .fco(\u2_Display/add87/c31 ),
    .fx({\u2_Display/n2770 [30],\u2_Display/n2770 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u31_al_u4896  (
    .a({open_n20400,\u2_Display/n2736 }),
    .c(2'b00),
    .d({open_n20405,1'b1}),
    .fci(\u2_Display/add87/c31 ),
    .f({open_n20422,\u2_Display/n2770 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u3_al_u4889  (
    .a({\u2_Display/n2762 ,\u2_Display/n2764 }),
    .b({\u2_Display/n2761 ,\u2_Display/n2763 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add87/c3 ),
    .f({\u2_Display/n2770 [5],\u2_Display/n2770 [3]}),
    .fco(\u2_Display/add87/c7 ),
    .fx({\u2_Display/n2770 [6],\u2_Display/n2770 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/u7_al_u4890  (
    .a({\u2_Display/n2758 ,\u2_Display/n2760 }),
    .b({\u2_Display/n2757 ,\u2_Display/n2759 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add87/c7 ),
    .f({\u2_Display/n2770 [9],\u2_Display/n2770 [7]}),
    .fco(\u2_Display/add87/c11 ),
    .fx({\u2_Display/n2770 [10],\u2_Display/n2770 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add87/ucin_al_u4888"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add87/ucin_al_u4888  (
    .a({\u2_Display/n2766 ,1'b1}),
    .b({\u2_Display/n2765 ,\u2_Display/n2767 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2770 [1],open_n20481}),
    .fco(\u2_Display/add87/c3 ),
    .fx({\u2_Display/n2770 [2],\u2_Display/n2770 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u11_al_u4900  (
    .a({\u2_Display/n2789 ,\u2_Display/n2791 }),
    .b({\u2_Display/n2788 ,\u2_Display/n2790 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add88/c11 ),
    .f({\u2_Display/n2805 [13],\u2_Display/n2805 [11]}),
    .fco(\u2_Display/add88/c15 ),
    .fx({\u2_Display/n2805 [14],\u2_Display/n2805 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u15_al_u4901  (
    .a({\u2_Display/n2785 ,\u2_Display/n2787 }),
    .b({\u2_Display/n2784 ,\u2_Display/n2786 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add88/c15 ),
    .f({\u2_Display/n2805 [17],\u2_Display/n2805 [15]}),
    .fco(\u2_Display/add88/c19 ),
    .fx({\u2_Display/n2805 [18],\u2_Display/n2805 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u19_al_u4902  (
    .a({\u2_Display/n2781 ,\u2_Display/n2783 }),
    .b({\u2_Display/n2780 ,\u2_Display/n2782 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add88/c19 ),
    .f({\u2_Display/n2805 [21],\u2_Display/n2805 [19]}),
    .fco(\u2_Display/add88/c23 ),
    .fx({\u2_Display/n2805 [22],\u2_Display/n2805 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u23_al_u4903  (
    .a({\u2_Display/n2777 ,\u2_Display/n2779 }),
    .b({\u2_Display/n2776 ,\u2_Display/n2778 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add88/c23 ),
    .f({\u2_Display/n2805 [25],\u2_Display/n2805 [23]}),
    .fco(\u2_Display/add88/c27 ),
    .fx({\u2_Display/n2805 [26],\u2_Display/n2805 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u27_al_u4904  (
    .a({\u2_Display/n2773 ,\u2_Display/n2775 }),
    .b({\u2_Display/n2772 ,\u2_Display/n2774 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add88/c27 ),
    .f({\u2_Display/n2805 [29],\u2_Display/n2805 [27]}),
    .fco(\u2_Display/add88/c31 ),
    .fx({\u2_Display/n2805 [30],\u2_Display/n2805 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u31_al_u4905  (
    .a({open_n20574,\u2_Display/n2771 }),
    .c(2'b00),
    .d({open_n20579,1'b1}),
    .fci(\u2_Display/add88/c31 ),
    .f({open_n20596,\u2_Display/n2805 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u3_al_u4898  (
    .a({\u2_Display/n2797 ,\u2_Display/n2799 }),
    .b({\u2_Display/n2796 ,\u2_Display/n2798 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add88/c3 ),
    .f({\u2_Display/n2805 [5],\u2_Display/n2805 [3]}),
    .fco(\u2_Display/add88/c7 ),
    .fx({\u2_Display/n2805 [6],\u2_Display/n2805 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/u7_al_u4899  (
    .a({\u2_Display/n2793 ,\u2_Display/n2795 }),
    .b({\u2_Display/n2792 ,\u2_Display/n2794 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add88/c7 ),
    .f({\u2_Display/n2805 [9],\u2_Display/n2805 [7]}),
    .fco(\u2_Display/add88/c11 ),
    .fx({\u2_Display/n2805 [10],\u2_Display/n2805 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add88/ucin_al_u4897"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add88/ucin_al_u4897  (
    .a({\u2_Display/n2801 ,1'b1}),
    .b({\u2_Display/n2800 ,\u2_Display/n2802 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2805 [1],open_n20655}),
    .fco(\u2_Display/add88/c3 ),
    .fx({\u2_Display/n2805 [2],\u2_Display/n2805 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u11_al_u4909  (
    .a({\u2_Display/n2824 ,\u2_Display/n2826 }),
    .b({\u2_Display/n2823 ,\u2_Display/n2825 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add89/c11 ),
    .f({\u2_Display/n2840 [13],\u2_Display/n2840 [11]}),
    .fco(\u2_Display/add89/c15 ),
    .fx({\u2_Display/n2840 [14],\u2_Display/n2840 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u15_al_u4910  (
    .a({\u2_Display/n2820 ,\u2_Display/n2822 }),
    .b({\u2_Display/n2819 ,\u2_Display/n2821 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add89/c15 ),
    .f({\u2_Display/n2840 [17],\u2_Display/n2840 [15]}),
    .fco(\u2_Display/add89/c19 ),
    .fx({\u2_Display/n2840 [18],\u2_Display/n2840 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u19_al_u4911  (
    .a({\u2_Display/n2816 ,\u2_Display/n2818 }),
    .b({\u2_Display/n2815 ,\u2_Display/n2817 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add89/c19 ),
    .f({\u2_Display/n2840 [21],\u2_Display/n2840 [19]}),
    .fco(\u2_Display/add89/c23 ),
    .fx({\u2_Display/n2840 [22],\u2_Display/n2840 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u23_al_u4912  (
    .a({\u2_Display/n2812 ,\u2_Display/n2814 }),
    .b({\u2_Display/n2811 ,\u2_Display/n2813 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add89/c23 ),
    .f({\u2_Display/n2840 [25],\u2_Display/n2840 [23]}),
    .fco(\u2_Display/add89/c27 ),
    .fx({\u2_Display/n2840 [26],\u2_Display/n2840 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u27_al_u4913  (
    .a({\u2_Display/n2808 ,\u2_Display/n2810 }),
    .b({\u2_Display/n2807 ,\u2_Display/n2809 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add89/c27 ),
    .f({\u2_Display/n2840 [29],\u2_Display/n2840 [27]}),
    .fco(\u2_Display/add89/c31 ),
    .fx({\u2_Display/n2840 [30],\u2_Display/n2840 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u31_al_u4914  (
    .a({open_n20748,\u2_Display/n2806 }),
    .c(2'b00),
    .d({open_n20753,1'b1}),
    .fci(\u2_Display/add89/c31 ),
    .f({open_n20770,\u2_Display/n2840 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u3_al_u4907  (
    .a({\u2_Display/n2832 ,\u2_Display/n2834 }),
    .b({\u2_Display/n2831 ,\u2_Display/n2833 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add89/c3 ),
    .f({\u2_Display/n2840 [5],\u2_Display/n2840 [3]}),
    .fco(\u2_Display/add89/c7 ),
    .fx({\u2_Display/n2840 [6],\u2_Display/n2840 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/u7_al_u4908  (
    .a({\u2_Display/n2828 ,\u2_Display/n2830 }),
    .b({\u2_Display/n2827 ,\u2_Display/n2829 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add89/c7 ),
    .f({\u2_Display/n2840 [9],\u2_Display/n2840 [7]}),
    .fco(\u2_Display/add89/c11 ),
    .fx({\u2_Display/n2840 [10],\u2_Display/n2840 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add89/ucin_al_u4906"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add89/ucin_al_u4906  (
    .a({\u2_Display/n2836 ,1'b1}),
    .b({\u2_Display/n2835 ,\u2_Display/n2837 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2840 [1],open_n20829}),
    .fco(\u2_Display/add89/c3 ),
    .fx({\u2_Display/n2840 [2],\u2_Display/n2840 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u11_al_u4918  (
    .a({\u2_Display/n2859 ,\u2_Display/n2861 }),
    .b({\u2_Display/n2858 ,\u2_Display/n2860 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add90/c11 ),
    .f({\u2_Display/n2875 [13],\u2_Display/n2875 [11]}),
    .fco(\u2_Display/add90/c15 ),
    .fx({\u2_Display/n2875 [14],\u2_Display/n2875 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u15_al_u4919  (
    .a({\u2_Display/n2855 ,\u2_Display/n2857 }),
    .b({\u2_Display/n2854 ,\u2_Display/n2856 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add90/c15 ),
    .f({\u2_Display/n2875 [17],\u2_Display/n2875 [15]}),
    .fco(\u2_Display/add90/c19 ),
    .fx({\u2_Display/n2875 [18],\u2_Display/n2875 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u19_al_u4920  (
    .a({\u2_Display/n2851 ,\u2_Display/n2853 }),
    .b({\u2_Display/n2850 ,\u2_Display/n2852 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b00),
    .fci(\u2_Display/add90/c19 ),
    .f({\u2_Display/n2875 [21],\u2_Display/n2875 [19]}),
    .fco(\u2_Display/add90/c23 ),
    .fx({\u2_Display/n2875 [22],\u2_Display/n2875 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u23_al_u4921  (
    .a({\u2_Display/n2847 ,\u2_Display/n2849 }),
    .b({\u2_Display/n2846 ,\u2_Display/n2848 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add90/c23 ),
    .f({\u2_Display/n2875 [25],\u2_Display/n2875 [23]}),
    .fco(\u2_Display/add90/c27 ),
    .fx({\u2_Display/n2875 [26],\u2_Display/n2875 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u27_al_u4922  (
    .a({\u2_Display/n2843 ,\u2_Display/n2845 }),
    .b({\u2_Display/n2842 ,\u2_Display/n2844 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add90/c27 ),
    .f({\u2_Display/n2875 [29],\u2_Display/n2875 [27]}),
    .fco(\u2_Display/add90/c31 ),
    .fx({\u2_Display/n2875 [30],\u2_Display/n2875 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u31_al_u4923  (
    .a({open_n20922,\u2_Display/n2841 }),
    .c(2'b00),
    .d({open_n20927,1'b1}),
    .fci(\u2_Display/add90/c31 ),
    .f({open_n20944,\u2_Display/n2875 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u3_al_u4916  (
    .a({\u2_Display/n2867 ,\u2_Display/n2869 }),
    .b({\u2_Display/n2866 ,\u2_Display/n2868 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add90/c3 ),
    .f({\u2_Display/n2875 [5],\u2_Display/n2875 [3]}),
    .fco(\u2_Display/add90/c7 ),
    .fx({\u2_Display/n2875 [6],\u2_Display/n2875 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/u7_al_u4917  (
    .a({\u2_Display/n2863 ,\u2_Display/n2865 }),
    .b({\u2_Display/n2862 ,\u2_Display/n2864 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add90/c7 ),
    .f({\u2_Display/n2875 [9],\u2_Display/n2875 [7]}),
    .fco(\u2_Display/add90/c11 ),
    .fx({\u2_Display/n2875 [10],\u2_Display/n2875 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add90/ucin_al_u4915"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add90/ucin_al_u4915  (
    .a({\u2_Display/n2871 ,1'b1}),
    .b({\u2_Display/n2870 ,\u2_Display/n2872 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2875 [1],open_n21003}),
    .fco(\u2_Display/add90/c3 ),
    .fx({\u2_Display/n2875 [2],\u2_Display/n2875 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u11_al_u4927  (
    .a({\u2_Display/n2894 ,\u2_Display/n2896 }),
    .b({\u2_Display/n2893 ,\u2_Display/n2895 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add91/c11 ),
    .f({\u2_Display/n2910 [13],\u2_Display/n2910 [11]}),
    .fco(\u2_Display/add91/c15 ),
    .fx({\u2_Display/n2910 [14],\u2_Display/n2910 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u15_al_u4928  (
    .a({\u2_Display/n2890 ,\u2_Display/n2892 }),
    .b({\u2_Display/n2889 ,\u2_Display/n2891 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add91/c15 ),
    .f({\u2_Display/n2910 [17],\u2_Display/n2910 [15]}),
    .fco(\u2_Display/add91/c19 ),
    .fx({\u2_Display/n2910 [18],\u2_Display/n2910 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u19_al_u4929  (
    .a({\u2_Display/n2886 ,\u2_Display/n2888 }),
    .b({\u2_Display/n2885 ,\u2_Display/n2887 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add91/c19 ),
    .f({\u2_Display/n2910 [21],\u2_Display/n2910 [19]}),
    .fco(\u2_Display/add91/c23 ),
    .fx({\u2_Display/n2910 [22],\u2_Display/n2910 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u23_al_u4930  (
    .a({\u2_Display/n2882 ,\u2_Display/n2884 }),
    .b({\u2_Display/n2881 ,\u2_Display/n2883 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add91/c23 ),
    .f({\u2_Display/n2910 [25],\u2_Display/n2910 [23]}),
    .fco(\u2_Display/add91/c27 ),
    .fx({\u2_Display/n2910 [26],\u2_Display/n2910 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u27_al_u4931  (
    .a({\u2_Display/n2878 ,\u2_Display/n2880 }),
    .b({\u2_Display/n2877 ,\u2_Display/n2879 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add91/c27 ),
    .f({\u2_Display/n2910 [29],\u2_Display/n2910 [27]}),
    .fco(\u2_Display/add91/c31 ),
    .fx({\u2_Display/n2910 [30],\u2_Display/n2910 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u31_al_u4932  (
    .a({open_n21096,\u2_Display/n2876 }),
    .c(2'b00),
    .d({open_n21101,1'b1}),
    .fci(\u2_Display/add91/c31 ),
    .f({open_n21118,\u2_Display/n2910 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u3_al_u4925  (
    .a({\u2_Display/n2902 ,\u2_Display/n2904 }),
    .b({\u2_Display/n2901 ,\u2_Display/n2903 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add91/c3 ),
    .f({\u2_Display/n2910 [5],\u2_Display/n2910 [3]}),
    .fco(\u2_Display/add91/c7 ),
    .fx({\u2_Display/n2910 [6],\u2_Display/n2910 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/u7_al_u4926  (
    .a({\u2_Display/n2898 ,\u2_Display/n2900 }),
    .b({\u2_Display/n2897 ,\u2_Display/n2899 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add91/c7 ),
    .f({\u2_Display/n2910 [9],\u2_Display/n2910 [7]}),
    .fco(\u2_Display/add91/c11 ),
    .fx({\u2_Display/n2910 [10],\u2_Display/n2910 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add91/ucin_al_u4924"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add91/ucin_al_u4924  (
    .a({\u2_Display/n2906 ,1'b1}),
    .b({\u2_Display/n2905 ,\u2_Display/n2907 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2910 [1],open_n21177}),
    .fco(\u2_Display/add91/c3 ),
    .fx({\u2_Display/n2910 [2],\u2_Display/n2910 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u11_al_u4936  (
    .a({\u2_Display/n2929 ,\u2_Display/n2931 }),
    .b({\u2_Display/n2928 ,\u2_Display/n2930 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add92/c11 ),
    .f({\u2_Display/n2945 [13],\u2_Display/n2945 [11]}),
    .fco(\u2_Display/add92/c15 ),
    .fx({\u2_Display/n2945 [14],\u2_Display/n2945 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u15_al_u4937  (
    .a({\u2_Display/n2925 ,\u2_Display/n2927 }),
    .b({\u2_Display/n2924 ,\u2_Display/n2926 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add92/c15 ),
    .f({\u2_Display/n2945 [17],\u2_Display/n2945 [15]}),
    .fco(\u2_Display/add92/c19 ),
    .fx({\u2_Display/n2945 [18],\u2_Display/n2945 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u19_al_u4938  (
    .a({\u2_Display/n2921 ,\u2_Display/n2923 }),
    .b({\u2_Display/n2920 ,\u2_Display/n2922 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add92/c19 ),
    .f({\u2_Display/n2945 [21],\u2_Display/n2945 [19]}),
    .fco(\u2_Display/add92/c23 ),
    .fx({\u2_Display/n2945 [22],\u2_Display/n2945 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u23_al_u4939  (
    .a({\u2_Display/n2917 ,\u2_Display/n2919 }),
    .b({\u2_Display/n2916 ,\u2_Display/n2918 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add92/c23 ),
    .f({\u2_Display/n2945 [25],\u2_Display/n2945 [23]}),
    .fco(\u2_Display/add92/c27 ),
    .fx({\u2_Display/n2945 [26],\u2_Display/n2945 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u27_al_u4940  (
    .a({\u2_Display/n2913 ,\u2_Display/n2915 }),
    .b({\u2_Display/n2912 ,\u2_Display/n2914 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add92/c27 ),
    .f({\u2_Display/n2945 [29],\u2_Display/n2945 [27]}),
    .fco(\u2_Display/add92/c31 ),
    .fx({\u2_Display/n2945 [30],\u2_Display/n2945 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u31_al_u4941  (
    .a({open_n21270,\u2_Display/n2911 }),
    .c(2'b00),
    .d({open_n21275,1'b1}),
    .fci(\u2_Display/add92/c31 ),
    .f({open_n21292,\u2_Display/n2945 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u3_al_u4934  (
    .a({\u2_Display/n2937 ,\u2_Display/n2939 }),
    .b({\u2_Display/n2936 ,\u2_Display/n2938 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add92/c3 ),
    .f({\u2_Display/n2945 [5],\u2_Display/n2945 [3]}),
    .fco(\u2_Display/add92/c7 ),
    .fx({\u2_Display/n2945 [6],\u2_Display/n2945 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/u7_al_u4935  (
    .a({\u2_Display/n2933 ,\u2_Display/n2935 }),
    .b({\u2_Display/n2932 ,\u2_Display/n2934 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add92/c7 ),
    .f({\u2_Display/n2945 [9],\u2_Display/n2945 [7]}),
    .fco(\u2_Display/add92/c11 ),
    .fx({\u2_Display/n2945 [10],\u2_Display/n2945 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add92/ucin_al_u4933"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add92/ucin_al_u4933  (
    .a({\u2_Display/n2941 ,1'b1}),
    .b({\u2_Display/n2940 ,\u2_Display/n2942 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2945 [1],open_n21351}),
    .fco(\u2_Display/add92/c3 ),
    .fx({\u2_Display/n2945 [2],\u2_Display/n2945 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u11_al_u4945  (
    .a({\u2_Display/n2964 ,\u2_Display/n2966 }),
    .b({\u2_Display/n2963 ,\u2_Display/n2965 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add93/c11 ),
    .f({\u2_Display/n2980 [13],\u2_Display/n2980 [11]}),
    .fco(\u2_Display/add93/c15 ),
    .fx({\u2_Display/n2980 [14],\u2_Display/n2980 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u15_al_u4946  (
    .a({\u2_Display/n2960 ,\u2_Display/n2962 }),
    .b({\u2_Display/n2959 ,\u2_Display/n2961 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add93/c15 ),
    .f({\u2_Display/n2980 [17],\u2_Display/n2980 [15]}),
    .fco(\u2_Display/add93/c19 ),
    .fx({\u2_Display/n2980 [18],\u2_Display/n2980 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u19_al_u4947  (
    .a({\u2_Display/n2956 ,\u2_Display/n2958 }),
    .b({\u2_Display/n2955 ,\u2_Display/n2957 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add93/c19 ),
    .f({\u2_Display/n2980 [21],\u2_Display/n2980 [19]}),
    .fco(\u2_Display/add93/c23 ),
    .fx({\u2_Display/n2980 [22],\u2_Display/n2980 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u23_al_u4948  (
    .a({\u2_Display/n2952 ,\u2_Display/n2954 }),
    .b({\u2_Display/n2951 ,\u2_Display/n2953 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add93/c23 ),
    .f({\u2_Display/n2980 [25],\u2_Display/n2980 [23]}),
    .fco(\u2_Display/add93/c27 ),
    .fx({\u2_Display/n2980 [26],\u2_Display/n2980 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u27_al_u4949  (
    .a({\u2_Display/n2948 ,\u2_Display/n2950 }),
    .b({\u2_Display/n2947 ,\u2_Display/n2949 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add93/c27 ),
    .f({\u2_Display/n2980 [29],\u2_Display/n2980 [27]}),
    .fco(\u2_Display/add93/c31 ),
    .fx({\u2_Display/n2980 [30],\u2_Display/n2980 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u31_al_u4950  (
    .a({open_n21444,\u2_Display/n2946 }),
    .c(2'b00),
    .d({open_n21449,1'b1}),
    .fci(\u2_Display/add93/c31 ),
    .f({open_n21466,\u2_Display/n2980 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u3_al_u4943  (
    .a({\u2_Display/n2972 ,\u2_Display/n2974 }),
    .b({\u2_Display/n2971 ,\u2_Display/n2973 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add93/c3 ),
    .f({\u2_Display/n2980 [5],\u2_Display/n2980 [3]}),
    .fco(\u2_Display/add93/c7 ),
    .fx({\u2_Display/n2980 [6],\u2_Display/n2980 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/u7_al_u4944  (
    .a({\u2_Display/n2968 ,\u2_Display/n2970 }),
    .b({\u2_Display/n2967 ,\u2_Display/n2969 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add93/c7 ),
    .f({\u2_Display/n2980 [9],\u2_Display/n2980 [7]}),
    .fco(\u2_Display/add93/c11 ),
    .fx({\u2_Display/n2980 [10],\u2_Display/n2980 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add93/ucin_al_u4942"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add93/ucin_al_u4942  (
    .a({\u2_Display/n2976 ,1'b1}),
    .b({\u2_Display/n2975 ,\u2_Display/n2977 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n2980 [1],open_n21525}),
    .fco(\u2_Display/add93/c3 ),
    .fx({\u2_Display/n2980 [2],\u2_Display/n2980 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u11_al_u4954  (
    .a({\u2_Display/n2999 ,\u2_Display/n3001 }),
    .b({\u2_Display/n2998 ,\u2_Display/n3000 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add94/c11 ),
    .f({\u2_Display/n3015 [13],\u2_Display/n3015 [11]}),
    .fco(\u2_Display/add94/c15 ),
    .fx({\u2_Display/n3015 [14],\u2_Display/n3015 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u15_al_u4955  (
    .a({\u2_Display/n2995 ,\u2_Display/n2997 }),
    .b({\u2_Display/n2994 ,\u2_Display/n2996 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b00),
    .fci(\u2_Display/add94/c15 ),
    .f({\u2_Display/n3015 [17],\u2_Display/n3015 [15]}),
    .fco(\u2_Display/add94/c19 ),
    .fx({\u2_Display/n3015 [18],\u2_Display/n3015 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u19_al_u4956  (
    .a({\u2_Display/n2991 ,\u2_Display/n2993 }),
    .b({\u2_Display/n2990 ,\u2_Display/n2992 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add94/c19 ),
    .f({\u2_Display/n3015 [21],\u2_Display/n3015 [19]}),
    .fco(\u2_Display/add94/c23 ),
    .fx({\u2_Display/n3015 [22],\u2_Display/n3015 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u23_al_u4957  (
    .a({\u2_Display/n2987 ,\u2_Display/n2989 }),
    .b({\u2_Display/n2986 ,\u2_Display/n2988 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add94/c23 ),
    .f({\u2_Display/n3015 [25],\u2_Display/n3015 [23]}),
    .fco(\u2_Display/add94/c27 ),
    .fx({\u2_Display/n3015 [26],\u2_Display/n3015 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u27_al_u4958  (
    .a({\u2_Display/n2983 ,\u2_Display/n2985 }),
    .b({\u2_Display/n2982 ,\u2_Display/n2984 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add94/c27 ),
    .f({\u2_Display/n3015 [29],\u2_Display/n3015 [27]}),
    .fco(\u2_Display/add94/c31 ),
    .fx({\u2_Display/n3015 [30],\u2_Display/n3015 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u31_al_u4959  (
    .a({open_n21618,\u2_Display/n2981 }),
    .c(2'b00),
    .d({open_n21623,1'b1}),
    .fci(\u2_Display/add94/c31 ),
    .f({open_n21640,\u2_Display/n3015 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u3_al_u4952  (
    .a({\u2_Display/n3007 ,\u2_Display/n3009 }),
    .b({\u2_Display/n3006 ,\u2_Display/n3008 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add94/c3 ),
    .f({\u2_Display/n3015 [5],\u2_Display/n3015 [3]}),
    .fco(\u2_Display/add94/c7 ),
    .fx({\u2_Display/n3015 [6],\u2_Display/n3015 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/u7_al_u4953  (
    .a({\u2_Display/n3003 ,\u2_Display/n3005 }),
    .b({\u2_Display/n3002 ,\u2_Display/n3004 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add94/c7 ),
    .f({\u2_Display/n3015 [9],\u2_Display/n3015 [7]}),
    .fco(\u2_Display/add94/c11 ),
    .fx({\u2_Display/n3015 [10],\u2_Display/n3015 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add94/ucin_al_u4951"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add94/ucin_al_u4951  (
    .a({\u2_Display/n3011 ,1'b1}),
    .b({\u2_Display/n3010 ,\u2_Display/n3012 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3015 [1],open_n21699}),
    .fco(\u2_Display/add94/c3 ),
    .fx({\u2_Display/n3015 [2],\u2_Display/n3015 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u11_al_u4963  (
    .a({\u2_Display/n3034 ,\u2_Display/n3036 }),
    .b({\u2_Display/n3033 ,\u2_Display/n3035 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add95/c11 ),
    .f({\u2_Display/n3050 [13],\u2_Display/n3050 [11]}),
    .fco(\u2_Display/add95/c15 ),
    .fx({\u2_Display/n3050 [14],\u2_Display/n3050 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u15_al_u4964  (
    .a({\u2_Display/n3030 ,\u2_Display/n3032 }),
    .b({\u2_Display/n3029 ,\u2_Display/n3031 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add95/c15 ),
    .f({\u2_Display/n3050 [17],\u2_Display/n3050 [15]}),
    .fco(\u2_Display/add95/c19 ),
    .fx({\u2_Display/n3050 [18],\u2_Display/n3050 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u19_al_u4965  (
    .a({\u2_Display/n3026 ,\u2_Display/n3028 }),
    .b({\u2_Display/n3025 ,\u2_Display/n3027 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add95/c19 ),
    .f({\u2_Display/n3050 [21],\u2_Display/n3050 [19]}),
    .fco(\u2_Display/add95/c23 ),
    .fx({\u2_Display/n3050 [22],\u2_Display/n3050 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u23_al_u4966  (
    .a({\u2_Display/n3022 ,\u2_Display/n3024 }),
    .b({\u2_Display/n3021 ,\u2_Display/n3023 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add95/c23 ),
    .f({\u2_Display/n3050 [25],\u2_Display/n3050 [23]}),
    .fco(\u2_Display/add95/c27 ),
    .fx({\u2_Display/n3050 [26],\u2_Display/n3050 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u27_al_u4967  (
    .a({\u2_Display/n3018 ,\u2_Display/n3020 }),
    .b({\u2_Display/n3017 ,\u2_Display/n3019 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add95/c27 ),
    .f({\u2_Display/n3050 [29],\u2_Display/n3050 [27]}),
    .fco(\u2_Display/add95/c31 ),
    .fx({\u2_Display/n3050 [30],\u2_Display/n3050 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u31_al_u4968  (
    .a({open_n21792,\u2_Display/n3016 }),
    .c(2'b00),
    .d({open_n21797,1'b1}),
    .fci(\u2_Display/add95/c31 ),
    .f({open_n21814,\u2_Display/n3050 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u3_al_u4961  (
    .a({\u2_Display/n3042 ,\u2_Display/n3044 }),
    .b({\u2_Display/n3041 ,\u2_Display/n3043 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add95/c3 ),
    .f({\u2_Display/n3050 [5],\u2_Display/n3050 [3]}),
    .fco(\u2_Display/add95/c7 ),
    .fx({\u2_Display/n3050 [6],\u2_Display/n3050 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/u7_al_u4962  (
    .a({\u2_Display/n3038 ,\u2_Display/n3040 }),
    .b({\u2_Display/n3037 ,\u2_Display/n3039 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add95/c7 ),
    .f({\u2_Display/n3050 [9],\u2_Display/n3050 [7]}),
    .fco(\u2_Display/add95/c11 ),
    .fx({\u2_Display/n3050 [10],\u2_Display/n3050 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add95/ucin_al_u4960"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add95/ucin_al_u4960  (
    .a({\u2_Display/n3046 ,1'b1}),
    .b({\u2_Display/n3045 ,\u2_Display/n3047 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3050 [1],open_n21873}),
    .fco(\u2_Display/add95/c3 ),
    .fx({\u2_Display/n3050 [2],\u2_Display/n3050 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u11_al_u4972  (
    .a({\u2_Display/n3069 ,\u2_Display/n3071 }),
    .b({\u2_Display/n3068 ,\u2_Display/n3070 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .fci(\u2_Display/add96/c11 ),
    .f({\u2_Display/n3085 [13],\u2_Display/n3085 [11]}),
    .fco(\u2_Display/add96/c15 ),
    .fx({\u2_Display/n3085 [14],\u2_Display/n3085 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u15_al_u4973  (
    .a({\u2_Display/n3065 ,\u2_Display/n3067 }),
    .b({\u2_Display/n3064 ,\u2_Display/n3066 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add96/c15 ),
    .f({\u2_Display/n3085 [17],\u2_Display/n3085 [15]}),
    .fco(\u2_Display/add96/c19 ),
    .fx({\u2_Display/n3085 [18],\u2_Display/n3085 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u19_al_u4974  (
    .a({\u2_Display/n3061 ,\u2_Display/n3063 }),
    .b({\u2_Display/n3060 ,\u2_Display/n3062 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b11),
    .fci(\u2_Display/add96/c19 ),
    .f({\u2_Display/n3085 [21],\u2_Display/n3085 [19]}),
    .fco(\u2_Display/add96/c23 ),
    .fx({\u2_Display/n3085 [22],\u2_Display/n3085 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u23_al_u4975  (
    .a({\u2_Display/n3057 ,\u2_Display/n3059 }),
    .b({\u2_Display/n3056 ,\u2_Display/n3058 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add96/c23 ),
    .f({\u2_Display/n3085 [25],\u2_Display/n3085 [23]}),
    .fco(\u2_Display/add96/c27 ),
    .fx({\u2_Display/n3085 [26],\u2_Display/n3085 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u27_al_u4976  (
    .a({\u2_Display/n3053 ,\u2_Display/n3055 }),
    .b({\u2_Display/n3052 ,\u2_Display/n3054 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add96/c27 ),
    .f({\u2_Display/n3085 [29],\u2_Display/n3085 [27]}),
    .fco(\u2_Display/add96/c31 ),
    .fx({\u2_Display/n3085 [30],\u2_Display/n3085 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u31_al_u4977  (
    .a({open_n21966,\u2_Display/n3051 }),
    .c(2'b00),
    .d({open_n21971,1'b1}),
    .fci(\u2_Display/add96/c31 ),
    .f({open_n21988,\u2_Display/n3085 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u3_al_u4970  (
    .a({\u2_Display/n3077 ,\u2_Display/n3079 }),
    .b({\u2_Display/n3076 ,\u2_Display/n3078 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add96/c3 ),
    .f({\u2_Display/n3085 [5],\u2_Display/n3085 [3]}),
    .fco(\u2_Display/add96/c7 ),
    .fx({\u2_Display/n3085 [6],\u2_Display/n3085 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/u7_al_u4971  (
    .a({\u2_Display/n3073 ,\u2_Display/n3075 }),
    .b({\u2_Display/n3072 ,\u2_Display/n3074 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add96/c7 ),
    .f({\u2_Display/n3085 [9],\u2_Display/n3085 [7]}),
    .fco(\u2_Display/add96/c11 ),
    .fx({\u2_Display/n3085 [10],\u2_Display/n3085 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add96/ucin_al_u4969"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add96/ucin_al_u4969  (
    .a({\u2_Display/n3081 ,1'b1}),
    .b({\u2_Display/n3080 ,\u2_Display/n3082 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3085 [1],open_n22047}),
    .fco(\u2_Display/add96/c3 ),
    .fx({\u2_Display/n3085 [2],\u2_Display/n3085 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u11_al_u4981  (
    .a({\u2_Display/n3104 ,\u2_Display/n3106 }),
    .b({\u2_Display/n3103 ,\u2_Display/n3105 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b10),
    .fci(\u2_Display/add97/c11 ),
    .f({\u2_Display/n3120 [13],\u2_Display/n3120 [11]}),
    .fco(\u2_Display/add97/c15 ),
    .fx({\u2_Display/n3120 [14],\u2_Display/n3120 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u15_al_u4982  (
    .a({\u2_Display/n3100 ,\u2_Display/n3102 }),
    .b({\u2_Display/n3099 ,\u2_Display/n3101 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b01),
    .fci(\u2_Display/add97/c15 ),
    .f({\u2_Display/n3120 [17],\u2_Display/n3120 [15]}),
    .fco(\u2_Display/add97/c19 ),
    .fx({\u2_Display/n3120 [18],\u2_Display/n3120 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u19_al_u4983  (
    .a({\u2_Display/n3096 ,\u2_Display/n3098 }),
    .b({\u2_Display/n3095 ,\u2_Display/n3097 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add97/c19 ),
    .f({\u2_Display/n3120 [21],\u2_Display/n3120 [19]}),
    .fco(\u2_Display/add97/c23 ),
    .fx({\u2_Display/n3120 [22],\u2_Display/n3120 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u23_al_u4984  (
    .a({\u2_Display/n3092 ,\u2_Display/n3094 }),
    .b({\u2_Display/n3091 ,\u2_Display/n3093 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add97/c23 ),
    .f({\u2_Display/n3120 [25],\u2_Display/n3120 [23]}),
    .fco(\u2_Display/add97/c27 ),
    .fx({\u2_Display/n3120 [26],\u2_Display/n3120 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u27_al_u4985  (
    .a({\u2_Display/n3088 ,\u2_Display/n3090 }),
    .b({\u2_Display/n3087 ,\u2_Display/n3089 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add97/c27 ),
    .f({\u2_Display/n3120 [29],\u2_Display/n3120 [27]}),
    .fco(\u2_Display/add97/c31 ),
    .fx({\u2_Display/n3120 [30],\u2_Display/n3120 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u31_al_u4986  (
    .a({open_n22140,\u2_Display/n3086 }),
    .c(2'b00),
    .d({open_n22145,1'b1}),
    .fci(\u2_Display/add97/c31 ),
    .f({open_n22162,\u2_Display/n3120 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u3_al_u4979  (
    .a({\u2_Display/n3112 ,\u2_Display/n3114 }),
    .b({\u2_Display/n3111 ,\u2_Display/n3113 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add97/c3 ),
    .f({\u2_Display/n3120 [5],\u2_Display/n3120 [3]}),
    .fco(\u2_Display/add97/c7 ),
    .fx({\u2_Display/n3120 [6],\u2_Display/n3120 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/u7_al_u4980  (
    .a({\u2_Display/n3108 ,\u2_Display/n3110 }),
    .b({\u2_Display/n3107 ,\u2_Display/n3109 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add97/c7 ),
    .f({\u2_Display/n3120 [9],\u2_Display/n3120 [7]}),
    .fco(\u2_Display/add97/c11 ),
    .fx({\u2_Display/n3120 [10],\u2_Display/n3120 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add97/ucin_al_u4978"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add97/ucin_al_u4978  (
    .a({\u2_Display/n3116 ,1'b1}),
    .b({\u2_Display/n3115 ,\u2_Display/n3117 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3120 [1],open_n22221}),
    .fco(\u2_Display/add97/c3 ),
    .fx({\u2_Display/n3120 [2],\u2_Display/n3120 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u11_al_u4990  (
    .a({\u2_Display/n3139 ,\u2_Display/n3141 }),
    .b({\u2_Display/n3138 ,\u2_Display/n3140 }),
    .c(2'b00),
    .d(2'b10),
    .e(2'b00),
    .fci(\u2_Display/add98/c11 ),
    .f({\u2_Display/n3155 [13],\u2_Display/n3155 [11]}),
    .fco(\u2_Display/add98/c15 ),
    .fx({\u2_Display/n3155 [14],\u2_Display/n3155 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u15_al_u4991  (
    .a({\u2_Display/n3135 ,\u2_Display/n3137 }),
    .b({\u2_Display/n3134 ,\u2_Display/n3136 }),
    .c(2'b00),
    .d(2'b01),
    .e(2'b11),
    .fci(\u2_Display/add98/c15 ),
    .f({\u2_Display/n3155 [17],\u2_Display/n3155 [15]}),
    .fco(\u2_Display/add98/c19 ),
    .fx({\u2_Display/n3155 [18],\u2_Display/n3155 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u19_al_u4992  (
    .a({\u2_Display/n3131 ,\u2_Display/n3133 }),
    .b({\u2_Display/n3130 ,\u2_Display/n3132 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add98/c19 ),
    .f({\u2_Display/n3155 [21],\u2_Display/n3155 [19]}),
    .fco(\u2_Display/add98/c23 ),
    .fx({\u2_Display/n3155 [22],\u2_Display/n3155 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u23_al_u4993  (
    .a({\u2_Display/n3127 ,\u2_Display/n3129 }),
    .b({\u2_Display/n3126 ,\u2_Display/n3128 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add98/c23 ),
    .f({\u2_Display/n3155 [25],\u2_Display/n3155 [23]}),
    .fco(\u2_Display/add98/c27 ),
    .fx({\u2_Display/n3155 [26],\u2_Display/n3155 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u27_al_u4994  (
    .a({\u2_Display/n3123 ,\u2_Display/n3125 }),
    .b({\u2_Display/n3122 ,\u2_Display/n3124 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add98/c27 ),
    .f({\u2_Display/n3155 [29],\u2_Display/n3155 [27]}),
    .fco(\u2_Display/add98/c31 ),
    .fx({\u2_Display/n3155 [30],\u2_Display/n3155 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u31_al_u4995  (
    .a({open_n22314,\u2_Display/n3121 }),
    .c(2'b00),
    .d({open_n22319,1'b1}),
    .fci(\u2_Display/add98/c31 ),
    .f({open_n22336,\u2_Display/n3155 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u3_al_u4988  (
    .a({\u2_Display/n3147 ,\u2_Display/n3149 }),
    .b({\u2_Display/n3146 ,\u2_Display/n3148 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add98/c3 ),
    .f({\u2_Display/n3155 [5],\u2_Display/n3155 [3]}),
    .fco(\u2_Display/add98/c7 ),
    .fx({\u2_Display/n3155 [6],\u2_Display/n3155 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/u7_al_u4989  (
    .a({\u2_Display/n3143 ,\u2_Display/n3145 }),
    .b({\u2_Display/n3142 ,\u2_Display/n3144 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add98/c7 ),
    .f({\u2_Display/n3155 [9],\u2_Display/n3155 [7]}),
    .fco(\u2_Display/add98/c11 ),
    .fx({\u2_Display/n3155 [10],\u2_Display/n3155 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add98/ucin_al_u4987"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add98/ucin_al_u4987  (
    .a({\u2_Display/n3151 ,1'b1}),
    .b({\u2_Display/n3150 ,\u2_Display/n3152 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3155 [1],open_n22395}),
    .fco(\u2_Display/add98/c3 ),
    .fx({\u2_Display/n3155 [2],\u2_Display/n3155 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u11_al_u4999  (
    .a({\u2_Display/n3174 ,\u2_Display/n3176 }),
    .b({\u2_Display/n3173 ,\u2_Display/n3175 }),
    .c(2'b00),
    .d(2'b00),
    .e(2'b11),
    .fci(\u2_Display/add99/c11 ),
    .f({\u2_Display/n3190 [13],\u2_Display/n3190 [11]}),
    .fco(\u2_Display/add99/c15 ),
    .fx({\u2_Display/n3190 [14],\u2_Display/n3190 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u15_al_u5000  (
    .a({\u2_Display/n3170 ,\u2_Display/n3172 }),
    .b({\u2_Display/n3169 ,\u2_Display/n3171 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b10),
    .fci(\u2_Display/add99/c15 ),
    .f({\u2_Display/n3190 [17],\u2_Display/n3190 [15]}),
    .fco(\u2_Display/add99/c19 ),
    .fx({\u2_Display/n3190 [18],\u2_Display/n3190 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u19_al_u5001  (
    .a({\u2_Display/n3166 ,\u2_Display/n3168 }),
    .b({\u2_Display/n3165 ,\u2_Display/n3167 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add99/c19 ),
    .f({\u2_Display/n3190 [21],\u2_Display/n3190 [19]}),
    .fco(\u2_Display/add99/c23 ),
    .fx({\u2_Display/n3190 [22],\u2_Display/n3190 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u23_al_u5002  (
    .a({\u2_Display/n3162 ,\u2_Display/n3164 }),
    .b({\u2_Display/n3161 ,\u2_Display/n3163 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add99/c23 ),
    .f({\u2_Display/n3190 [25],\u2_Display/n3190 [23]}),
    .fco(\u2_Display/add99/c27 ),
    .fx({\u2_Display/n3190 [26],\u2_Display/n3190 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u27_al_u5003  (
    .a({\u2_Display/n3158 ,\u2_Display/n3160 }),
    .b({\u2_Display/n3157 ,\u2_Display/n3159 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add99/c27 ),
    .f({\u2_Display/n3190 [29],\u2_Display/n3190 [27]}),
    .fco(\u2_Display/add99/c31 ),
    .fx({\u2_Display/n3190 [30],\u2_Display/n3190 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u31_al_u5004  (
    .a({open_n22488,\u2_Display/n3156 }),
    .c(2'b00),
    .d({open_n22493,1'b1}),
    .fci(\u2_Display/add99/c31 ),
    .f({open_n22510,\u2_Display/n3190 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u3_al_u4997  (
    .a({\u2_Display/n3182 ,\u2_Display/n3184 }),
    .b({\u2_Display/n3181 ,\u2_Display/n3183 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .fci(\u2_Display/add99/c3 ),
    .f({\u2_Display/n3190 [5],\u2_Display/n3190 [3]}),
    .fco(\u2_Display/add99/c7 ),
    .fx({\u2_Display/n3190 [6],\u2_Display/n3190 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/u7_al_u4998  (
    .a({\u2_Display/n3178 ,\u2_Display/n3180 }),
    .b({\u2_Display/n3177 ,\u2_Display/n3179 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b01),
    .fci(\u2_Display/add99/c7 ),
    .f({\u2_Display/n3190 [9],\u2_Display/n3190 [7]}),
    .fco(\u2_Display/add99/c11 ),
    .fx({\u2_Display/n3190 [10],\u2_Display/n3190 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/add99/ucin_al_u4996"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/add99/ucin_al_u4996  (
    .a({\u2_Display/n3186 ,1'b1}),
    .b({\u2_Display/n3185 ,\u2_Display/n3187 }),
    .c(2'b00),
    .d(2'b11),
    .e(2'b11),
    .f({\u2_Display/n3190 [1],open_n22569}),
    .fco(\u2_Display/add99/c3 ),
    .fx({\u2_Display/n3190 [2],\u2_Display/n3190 [0]}));
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/clk1s_reg  (
    .ce(\u2_Display/n35 ),
    .clk(clk_vga),
    .d(\u2_Display/n36 ),
    .q(\u2_Display/clk1s ));  // source/rtl/Display.v(61)
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_0|u2_Display/lt0_2_cin  (
    .a({lcd_xpos[0],1'b0}),
    .b({\u2_Display/i [0],open_n22573}),
    .fco(\u2_Display/lt0_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_10|u2_Display/lt0_2_9  (
    .a(lcd_xpos[10:9]),
    .b(\u2_Display/n43 [2:1]),
    .fci(\u2_Display/lt0_2_c9 ),
    .fco(\u2_Display/lt0_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_2|u2_Display/lt0_2_1  (
    .a(lcd_xpos[2:1]),
    .b(\u2_Display/i [2:1]),
    .fci(\u2_Display/lt0_2_c1 ),
    .fco(\u2_Display/lt0_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_4|u2_Display/lt0_2_3  (
    .a(lcd_xpos[4:3]),
    .b(\u2_Display/i [4:3]),
    .fci(\u2_Display/lt0_2_c3 ),
    .fco(\u2_Display/lt0_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_6|u2_Display/lt0_2_5  (
    .a(lcd_xpos[6:5]),
    .b(\u2_Display/i [6:5]),
    .fci(\u2_Display/lt0_2_c5 ),
    .fco(\u2_Display/lt0_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_8|u2_Display/lt0_2_7  (
    .a(lcd_xpos[8:7]),
    .b({\u2_Display/n43 [0],\u2_Display/i [7]}),
    .fci(\u2_Display/lt0_2_c7 ),
    .fco(\u2_Display/lt0_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt0_2_0|u2_Display/lt0_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt0_2_cout|u2_Display/lt0_2_11  (
    .a({1'b0,lcd_xpos[11]}),
    .b({1'b1,\u2_Display/add2_2_co }),
    .fci(\u2_Display/lt0_2_c11 ),
    .f({\u2_Display/n44 ,open_n22737}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_0|u2_Display/lt100_cin  (
    .a({\u2_Display/n3082 ,1'b0}),
    .b({1'b0,open_n22743}),
    .fco(\u2_Display/lt100_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_10|u2_Display/lt100_9  (
    .a({\u2_Display/n3072 ,\u2_Display/n3073 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c9 ),
    .fco(\u2_Display/lt100_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_12|u2_Display/lt100_11  (
    .a({\u2_Display/n3070 ,\u2_Display/n3071 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c11 ),
    .fco(\u2_Display/lt100_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_14|u2_Display/lt100_13  (
    .a({\u2_Display/n3068 ,\u2_Display/n3069 }),
    .b(2'b11),
    .fci(\u2_Display/lt100_c13 ),
    .fco(\u2_Display/lt100_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_16|u2_Display/lt100_15  (
    .a({\u2_Display/n3066 ,\u2_Display/n3067 }),
    .b(2'b10),
    .fci(\u2_Display/lt100_c15 ),
    .fco(\u2_Display/lt100_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_18|u2_Display/lt100_17  (
    .a({\u2_Display/n3064 ,\u2_Display/n3065 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c17 ),
    .fco(\u2_Display/lt100_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_20|u2_Display/lt100_19  (
    .a({\u2_Display/n3062 ,\u2_Display/n3063 }),
    .b(2'b01),
    .fci(\u2_Display/lt100_c19 ),
    .fco(\u2_Display/lt100_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_22|u2_Display/lt100_21  (
    .a({\u2_Display/n3060 ,\u2_Display/n3061 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c21 ),
    .fco(\u2_Display/lt100_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_24|u2_Display/lt100_23  (
    .a({\u2_Display/n3058 ,\u2_Display/n3059 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c23 ),
    .fco(\u2_Display/lt100_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_26|u2_Display/lt100_25  (
    .a({\u2_Display/n3056 ,\u2_Display/n3057 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c25 ),
    .fco(\u2_Display/lt100_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_28|u2_Display/lt100_27  (
    .a({\u2_Display/n3054 ,\u2_Display/n3055 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c27 ),
    .fco(\u2_Display/lt100_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_2|u2_Display/lt100_1  (
    .a({\u2_Display/n3080 ,\u2_Display/n3081 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c1 ),
    .fco(\u2_Display/lt100_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_30|u2_Display/lt100_29  (
    .a({\u2_Display/n3052 ,\u2_Display/n3053 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c29 ),
    .fco(\u2_Display/lt100_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_4|u2_Display/lt100_3  (
    .a({\u2_Display/n3078 ,\u2_Display/n3079 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c3 ),
    .fco(\u2_Display/lt100_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_6|u2_Display/lt100_5  (
    .a({\u2_Display/n3076 ,\u2_Display/n3077 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c5 ),
    .fco(\u2_Display/lt100_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_8|u2_Display/lt100_7  (
    .a({\u2_Display/n3074 ,\u2_Display/n3075 }),
    .b(2'b00),
    .fci(\u2_Display/lt100_c7 ),
    .fco(\u2_Display/lt100_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt100_0|u2_Display/lt100_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt100_cout|u2_Display/lt100_31  (
    .a({1'b0,\u2_Display/n3051 }),
    .b(2'b10),
    .fci(\u2_Display/lt100_c31 ),
    .f({\u2_Display/n3083 ,open_n23147}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_0|u2_Display/lt101_cin  (
    .a({\u2_Display/n3117 ,1'b0}),
    .b({1'b0,open_n23153}),
    .fco(\u2_Display/lt101_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_10|u2_Display/lt101_9  (
    .a({\u2_Display/n3107 ,\u2_Display/n3108 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c9 ),
    .fco(\u2_Display/lt101_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_12|u2_Display/lt101_11  (
    .a({\u2_Display/n3105 ,\u2_Display/n3106 }),
    .b(2'b10),
    .fci(\u2_Display/lt101_c11 ),
    .fco(\u2_Display/lt101_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_14|u2_Display/lt101_13  (
    .a({\u2_Display/n3103 ,\u2_Display/n3104 }),
    .b(2'b01),
    .fci(\u2_Display/lt101_c13 ),
    .fco(\u2_Display/lt101_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_16|u2_Display/lt101_15  (
    .a({\u2_Display/n3101 ,\u2_Display/n3102 }),
    .b(2'b01),
    .fci(\u2_Display/lt101_c15 ),
    .fco(\u2_Display/lt101_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_18|u2_Display/lt101_17  (
    .a({\u2_Display/n3099 ,\u2_Display/n3100 }),
    .b(2'b10),
    .fci(\u2_Display/lt101_c17 ),
    .fco(\u2_Display/lt101_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_20|u2_Display/lt101_19  (
    .a({\u2_Display/n3097 ,\u2_Display/n3098 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c19 ),
    .fco(\u2_Display/lt101_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_22|u2_Display/lt101_21  (
    .a({\u2_Display/n3095 ,\u2_Display/n3096 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c21 ),
    .fco(\u2_Display/lt101_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_24|u2_Display/lt101_23  (
    .a({\u2_Display/n3093 ,\u2_Display/n3094 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c23 ),
    .fco(\u2_Display/lt101_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_26|u2_Display/lt101_25  (
    .a({\u2_Display/n3091 ,\u2_Display/n3092 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c25 ),
    .fco(\u2_Display/lt101_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_28|u2_Display/lt101_27  (
    .a({\u2_Display/n3089 ,\u2_Display/n3090 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c27 ),
    .fco(\u2_Display/lt101_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_2|u2_Display/lt101_1  (
    .a({\u2_Display/n3115 ,\u2_Display/n3116 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c1 ),
    .fco(\u2_Display/lt101_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_30|u2_Display/lt101_29  (
    .a({\u2_Display/n3087 ,\u2_Display/n3088 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c29 ),
    .fco(\u2_Display/lt101_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_4|u2_Display/lt101_3  (
    .a({\u2_Display/n3113 ,\u2_Display/n3114 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c3 ),
    .fco(\u2_Display/lt101_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_6|u2_Display/lt101_5  (
    .a({\u2_Display/n3111 ,\u2_Display/n3112 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c5 ),
    .fco(\u2_Display/lt101_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_8|u2_Display/lt101_7  (
    .a({\u2_Display/n3109 ,\u2_Display/n3110 }),
    .b(2'b00),
    .fci(\u2_Display/lt101_c7 ),
    .fco(\u2_Display/lt101_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt101_0|u2_Display/lt101_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt101_cout|u2_Display/lt101_31  (
    .a({1'b0,\u2_Display/n3086 }),
    .b(2'b10),
    .fci(\u2_Display/lt101_c31 ),
    .f({\u2_Display/n3118 ,open_n23557}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_0|u2_Display/lt102_cin  (
    .a({\u2_Display/n3152 ,1'b0}),
    .b({1'b0,open_n23563}),
    .fco(\u2_Display/lt102_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_10|u2_Display/lt102_9  (
    .a({\u2_Display/n3142 ,\u2_Display/n3143 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c9 ),
    .fco(\u2_Display/lt102_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_12|u2_Display/lt102_11  (
    .a({\u2_Display/n3140 ,\u2_Display/n3141 }),
    .b(2'b11),
    .fci(\u2_Display/lt102_c11 ),
    .fco(\u2_Display/lt102_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_14|u2_Display/lt102_13  (
    .a({\u2_Display/n3138 ,\u2_Display/n3139 }),
    .b(2'b10),
    .fci(\u2_Display/lt102_c13 ),
    .fco(\u2_Display/lt102_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_16|u2_Display/lt102_15  (
    .a({\u2_Display/n3136 ,\u2_Display/n3137 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c15 ),
    .fco(\u2_Display/lt102_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_18|u2_Display/lt102_17  (
    .a({\u2_Display/n3134 ,\u2_Display/n3135 }),
    .b(2'b01),
    .fci(\u2_Display/lt102_c17 ),
    .fco(\u2_Display/lt102_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_20|u2_Display/lt102_19  (
    .a({\u2_Display/n3132 ,\u2_Display/n3133 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c19 ),
    .fco(\u2_Display/lt102_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_22|u2_Display/lt102_21  (
    .a({\u2_Display/n3130 ,\u2_Display/n3131 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c21 ),
    .fco(\u2_Display/lt102_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_24|u2_Display/lt102_23  (
    .a({\u2_Display/n3128 ,\u2_Display/n3129 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c23 ),
    .fco(\u2_Display/lt102_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_26|u2_Display/lt102_25  (
    .a({\u2_Display/n3126 ,\u2_Display/n3127 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c25 ),
    .fco(\u2_Display/lt102_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_28|u2_Display/lt102_27  (
    .a({\u2_Display/n3124 ,\u2_Display/n3125 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c27 ),
    .fco(\u2_Display/lt102_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_2|u2_Display/lt102_1  (
    .a({\u2_Display/n3150 ,\u2_Display/n3151 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c1 ),
    .fco(\u2_Display/lt102_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_30|u2_Display/lt102_29  (
    .a({\u2_Display/n3122 ,\u2_Display/n3123 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c29 ),
    .fco(\u2_Display/lt102_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_4|u2_Display/lt102_3  (
    .a({\u2_Display/n3148 ,\u2_Display/n3149 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c3 ),
    .fco(\u2_Display/lt102_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_6|u2_Display/lt102_5  (
    .a({\u2_Display/n3146 ,\u2_Display/n3147 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c5 ),
    .fco(\u2_Display/lt102_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_8|u2_Display/lt102_7  (
    .a({\u2_Display/n3144 ,\u2_Display/n3145 }),
    .b(2'b00),
    .fci(\u2_Display/lt102_c7 ),
    .fco(\u2_Display/lt102_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt102_0|u2_Display/lt102_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt102_cout|u2_Display/lt102_31  (
    .a({1'b0,\u2_Display/n3121 }),
    .b(2'b10),
    .fci(\u2_Display/lt102_c31 ),
    .f({\u2_Display/n3153 ,open_n23967}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_0|u2_Display/lt103_cin  (
    .a({\u2_Display/n3187 ,1'b0}),
    .b({1'b0,open_n23973}),
    .fco(\u2_Display/lt103_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_10|u2_Display/lt103_9  (
    .a({\u2_Display/n3177 ,\u2_Display/n3178 }),
    .b(2'b10),
    .fci(\u2_Display/lt103_c9 ),
    .fco(\u2_Display/lt103_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_12|u2_Display/lt103_11  (
    .a({\u2_Display/n3175 ,\u2_Display/n3176 }),
    .b(2'b01),
    .fci(\u2_Display/lt103_c11 ),
    .fco(\u2_Display/lt103_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_14|u2_Display/lt103_13  (
    .a({\u2_Display/n3173 ,\u2_Display/n3174 }),
    .b(2'b01),
    .fci(\u2_Display/lt103_c13 ),
    .fco(\u2_Display/lt103_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_16|u2_Display/lt103_15  (
    .a({\u2_Display/n3171 ,\u2_Display/n3172 }),
    .b(2'b10),
    .fci(\u2_Display/lt103_c15 ),
    .fco(\u2_Display/lt103_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_18|u2_Display/lt103_17  (
    .a({\u2_Display/n3169 ,\u2_Display/n3170 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c17 ),
    .fco(\u2_Display/lt103_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_20|u2_Display/lt103_19  (
    .a({\u2_Display/n3167 ,\u2_Display/n3168 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c19 ),
    .fco(\u2_Display/lt103_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_22|u2_Display/lt103_21  (
    .a({\u2_Display/n3165 ,\u2_Display/n3166 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c21 ),
    .fco(\u2_Display/lt103_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_24|u2_Display/lt103_23  (
    .a({\u2_Display/n3163 ,\u2_Display/n3164 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c23 ),
    .fco(\u2_Display/lt103_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_26|u2_Display/lt103_25  (
    .a({\u2_Display/n3161 ,\u2_Display/n3162 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c25 ),
    .fco(\u2_Display/lt103_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_28|u2_Display/lt103_27  (
    .a({\u2_Display/n3159 ,\u2_Display/n3160 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c27 ),
    .fco(\u2_Display/lt103_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_2|u2_Display/lt103_1  (
    .a({\u2_Display/n3185 ,\u2_Display/n3186 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c1 ),
    .fco(\u2_Display/lt103_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_30|u2_Display/lt103_29  (
    .a({\u2_Display/n3157 ,\u2_Display/n3158 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c29 ),
    .fco(\u2_Display/lt103_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_4|u2_Display/lt103_3  (
    .a({\u2_Display/n3183 ,\u2_Display/n3184 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c3 ),
    .fco(\u2_Display/lt103_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_6|u2_Display/lt103_5  (
    .a({\u2_Display/n3181 ,\u2_Display/n3182 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c5 ),
    .fco(\u2_Display/lt103_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_8|u2_Display/lt103_7  (
    .a({\u2_Display/n3179 ,\u2_Display/n3180 }),
    .b(2'b00),
    .fci(\u2_Display/lt103_c7 ),
    .fco(\u2_Display/lt103_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt103_0|u2_Display/lt103_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt103_cout|u2_Display/lt103_31  (
    .a({1'b0,\u2_Display/n3156 }),
    .b(2'b10),
    .fci(\u2_Display/lt103_c31 ),
    .f({\u2_Display/n3188 ,open_n24377}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_0|u2_Display/lt104_cin  (
    .a({\u2_Display/n3222 ,1'b0}),
    .b({1'b0,open_n24383}),
    .fco(\u2_Display/lt104_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_10|u2_Display/lt104_9  (
    .a({\u2_Display/n3212 ,\u2_Display/n3213 }),
    .b(2'b11),
    .fci(\u2_Display/lt104_c9 ),
    .fco(\u2_Display/lt104_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_12|u2_Display/lt104_11  (
    .a({\u2_Display/n3210 ,\u2_Display/n3211 }),
    .b(2'b10),
    .fci(\u2_Display/lt104_c11 ),
    .fco(\u2_Display/lt104_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_14|u2_Display/lt104_13  (
    .a({\u2_Display/n3208 ,\u2_Display/n3209 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c13 ),
    .fco(\u2_Display/lt104_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_16|u2_Display/lt104_15  (
    .a({\u2_Display/n3206 ,\u2_Display/n3207 }),
    .b(2'b01),
    .fci(\u2_Display/lt104_c15 ),
    .fco(\u2_Display/lt104_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_18|u2_Display/lt104_17  (
    .a({\u2_Display/n3204 ,\u2_Display/n3205 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c17 ),
    .fco(\u2_Display/lt104_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_20|u2_Display/lt104_19  (
    .a({\u2_Display/n3202 ,\u2_Display/n3203 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c19 ),
    .fco(\u2_Display/lt104_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_22|u2_Display/lt104_21  (
    .a({\u2_Display/n3200 ,\u2_Display/n3201 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c21 ),
    .fco(\u2_Display/lt104_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_24|u2_Display/lt104_23  (
    .a({\u2_Display/n3198 ,\u2_Display/n3199 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c23 ),
    .fco(\u2_Display/lt104_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_26|u2_Display/lt104_25  (
    .a({\u2_Display/n3196 ,\u2_Display/n3197 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c25 ),
    .fco(\u2_Display/lt104_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_28|u2_Display/lt104_27  (
    .a({\u2_Display/n3194 ,\u2_Display/n3195 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c27 ),
    .fco(\u2_Display/lt104_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_2|u2_Display/lt104_1  (
    .a({\u2_Display/n3220 ,\u2_Display/n3221 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c1 ),
    .fco(\u2_Display/lt104_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_30|u2_Display/lt104_29  (
    .a({\u2_Display/n3192 ,\u2_Display/n3193 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c29 ),
    .fco(\u2_Display/lt104_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_4|u2_Display/lt104_3  (
    .a({\u2_Display/n3218 ,\u2_Display/n3219 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c3 ),
    .fco(\u2_Display/lt104_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_6|u2_Display/lt104_5  (
    .a({\u2_Display/n3216 ,\u2_Display/n3217 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c5 ),
    .fco(\u2_Display/lt104_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_8|u2_Display/lt104_7  (
    .a({\u2_Display/n3214 ,\u2_Display/n3215 }),
    .b(2'b00),
    .fci(\u2_Display/lt104_c7 ),
    .fco(\u2_Display/lt104_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt104_0|u2_Display/lt104_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt104_cout|u2_Display/lt104_31  (
    .a({1'b0,\u2_Display/n3191 }),
    .b(2'b10),
    .fci(\u2_Display/lt104_c31 ),
    .f({\u2_Display/n3223 ,open_n24787}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_0|u2_Display/lt105_cin  (
    .a({\u2_Display/n3257 ,1'b0}),
    .b({1'b0,open_n24793}),
    .fco(\u2_Display/lt105_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_10|u2_Display/lt105_9  (
    .a({\u2_Display/n3247 ,\u2_Display/n3248 }),
    .b(2'b01),
    .fci(\u2_Display/lt105_c9 ),
    .fco(\u2_Display/lt105_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_12|u2_Display/lt105_11  (
    .a({\u2_Display/n3245 ,\u2_Display/n3246 }),
    .b(2'b01),
    .fci(\u2_Display/lt105_c11 ),
    .fco(\u2_Display/lt105_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_14|u2_Display/lt105_13  (
    .a({\u2_Display/n3243 ,\u2_Display/n3244 }),
    .b(2'b10),
    .fci(\u2_Display/lt105_c13 ),
    .fco(\u2_Display/lt105_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_16|u2_Display/lt105_15  (
    .a({\u2_Display/n3241 ,\u2_Display/n3242 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c15 ),
    .fco(\u2_Display/lt105_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_18|u2_Display/lt105_17  (
    .a({\u2_Display/n3239 ,\u2_Display/n3240 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c17 ),
    .fco(\u2_Display/lt105_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_20|u2_Display/lt105_19  (
    .a({\u2_Display/n3237 ,\u2_Display/n3238 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c19 ),
    .fco(\u2_Display/lt105_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_22|u2_Display/lt105_21  (
    .a({\u2_Display/n3235 ,\u2_Display/n3236 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c21 ),
    .fco(\u2_Display/lt105_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_24|u2_Display/lt105_23  (
    .a({\u2_Display/n3233 ,\u2_Display/n3234 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c23 ),
    .fco(\u2_Display/lt105_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_26|u2_Display/lt105_25  (
    .a({\u2_Display/n3231 ,\u2_Display/n3232 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c25 ),
    .fco(\u2_Display/lt105_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_28|u2_Display/lt105_27  (
    .a({\u2_Display/n3229 ,\u2_Display/n3230 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c27 ),
    .fco(\u2_Display/lt105_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_2|u2_Display/lt105_1  (
    .a({\u2_Display/n3255 ,\u2_Display/n3256 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c1 ),
    .fco(\u2_Display/lt105_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_30|u2_Display/lt105_29  (
    .a({\u2_Display/n3227 ,\u2_Display/n3228 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c29 ),
    .fco(\u2_Display/lt105_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_4|u2_Display/lt105_3  (
    .a({\u2_Display/n3253 ,\u2_Display/n3254 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c3 ),
    .fco(\u2_Display/lt105_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_6|u2_Display/lt105_5  (
    .a({\u2_Display/n3251 ,\u2_Display/n3252 }),
    .b(2'b00),
    .fci(\u2_Display/lt105_c5 ),
    .fco(\u2_Display/lt105_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_8|u2_Display/lt105_7  (
    .a({\u2_Display/n3249 ,\u2_Display/n3250 }),
    .b(2'b10),
    .fci(\u2_Display/lt105_c7 ),
    .fco(\u2_Display/lt105_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt105_0|u2_Display/lt105_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt105_cout|u2_Display/lt105_31  (
    .a({1'b0,\u2_Display/n3226 }),
    .b(2'b10),
    .fci(\u2_Display/lt105_c31 ),
    .f({\u2_Display/n3258 ,open_n25197}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_0|u2_Display/lt106_cin  (
    .a({\u2_Display/n3292 ,1'b0}),
    .b({1'b0,open_n25203}),
    .fco(\u2_Display/lt106_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_10|u2_Display/lt106_9  (
    .a({\u2_Display/n3282 ,\u2_Display/n3283 }),
    .b(2'b10),
    .fci(\u2_Display/lt106_c9 ),
    .fco(\u2_Display/lt106_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_12|u2_Display/lt106_11  (
    .a({\u2_Display/n3280 ,\u2_Display/n3281 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c11 ),
    .fco(\u2_Display/lt106_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_14|u2_Display/lt106_13  (
    .a({\u2_Display/n3278 ,\u2_Display/n3279 }),
    .b(2'b01),
    .fci(\u2_Display/lt106_c13 ),
    .fco(\u2_Display/lt106_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_16|u2_Display/lt106_15  (
    .a({\u2_Display/n3276 ,\u2_Display/n3277 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c15 ),
    .fco(\u2_Display/lt106_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_18|u2_Display/lt106_17  (
    .a({\u2_Display/n3274 ,\u2_Display/n3275 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c17 ),
    .fco(\u2_Display/lt106_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_20|u2_Display/lt106_19  (
    .a({\u2_Display/n3272 ,\u2_Display/n3273 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c19 ),
    .fco(\u2_Display/lt106_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_22|u2_Display/lt106_21  (
    .a({\u2_Display/n3270 ,\u2_Display/n3271 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c21 ),
    .fco(\u2_Display/lt106_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_24|u2_Display/lt106_23  (
    .a({\u2_Display/n3268 ,\u2_Display/n3269 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c23 ),
    .fco(\u2_Display/lt106_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_26|u2_Display/lt106_25  (
    .a({\u2_Display/n3266 ,\u2_Display/n3267 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c25 ),
    .fco(\u2_Display/lt106_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_28|u2_Display/lt106_27  (
    .a({\u2_Display/n3264 ,\u2_Display/n3265 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c27 ),
    .fco(\u2_Display/lt106_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_2|u2_Display/lt106_1  (
    .a({\u2_Display/n3290 ,\u2_Display/n3291 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c1 ),
    .fco(\u2_Display/lt106_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_30|u2_Display/lt106_29  (
    .a({\u2_Display/n3262 ,\u2_Display/n3263 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c29 ),
    .fco(\u2_Display/lt106_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_4|u2_Display/lt106_3  (
    .a({\u2_Display/n3288 ,\u2_Display/n3289 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c3 ),
    .fco(\u2_Display/lt106_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_6|u2_Display/lt106_5  (
    .a({\u2_Display/n3286 ,\u2_Display/n3287 }),
    .b(2'b00),
    .fci(\u2_Display/lt106_c5 ),
    .fco(\u2_Display/lt106_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_8|u2_Display/lt106_7  (
    .a({\u2_Display/n3284 ,\u2_Display/n3285 }),
    .b(2'b11),
    .fci(\u2_Display/lt106_c7 ),
    .fco(\u2_Display/lt106_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt106_0|u2_Display/lt106_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt106_cout|u2_Display/lt106_31  (
    .a({1'b0,\u2_Display/n3261 }),
    .b(2'b10),
    .fci(\u2_Display/lt106_c31 ),
    .f({\u2_Display/n3293 ,open_n25607}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_0|u2_Display/lt107_cin  (
    .a({\u2_Display/n3327 ,1'b0}),
    .b({1'b0,open_n25613}),
    .fco(\u2_Display/lt107_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_10|u2_Display/lt107_9  (
    .a({\u2_Display/n3317 ,\u2_Display/n3318 }),
    .b(2'b01),
    .fci(\u2_Display/lt107_c9 ),
    .fco(\u2_Display/lt107_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_12|u2_Display/lt107_11  (
    .a({\u2_Display/n3315 ,\u2_Display/n3316 }),
    .b(2'b10),
    .fci(\u2_Display/lt107_c11 ),
    .fco(\u2_Display/lt107_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_14|u2_Display/lt107_13  (
    .a({\u2_Display/n3313 ,\u2_Display/n3314 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c13 ),
    .fco(\u2_Display/lt107_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_16|u2_Display/lt107_15  (
    .a({\u2_Display/n3311 ,\u2_Display/n3312 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c15 ),
    .fco(\u2_Display/lt107_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_18|u2_Display/lt107_17  (
    .a({\u2_Display/n3309 ,\u2_Display/n3310 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c17 ),
    .fco(\u2_Display/lt107_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_20|u2_Display/lt107_19  (
    .a({\u2_Display/n3307 ,\u2_Display/n3308 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c19 ),
    .fco(\u2_Display/lt107_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_22|u2_Display/lt107_21  (
    .a({\u2_Display/n3305 ,\u2_Display/n3306 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c21 ),
    .fco(\u2_Display/lt107_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_24|u2_Display/lt107_23  (
    .a({\u2_Display/n3303 ,\u2_Display/n3304 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c23 ),
    .fco(\u2_Display/lt107_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_26|u2_Display/lt107_25  (
    .a({\u2_Display/n3301 ,\u2_Display/n3302 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c25 ),
    .fco(\u2_Display/lt107_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_28|u2_Display/lt107_27  (
    .a({\u2_Display/n3299 ,\u2_Display/n3300 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c27 ),
    .fco(\u2_Display/lt107_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_2|u2_Display/lt107_1  (
    .a({\u2_Display/n3325 ,\u2_Display/n3326 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c1 ),
    .fco(\u2_Display/lt107_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_30|u2_Display/lt107_29  (
    .a({\u2_Display/n3297 ,\u2_Display/n3298 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c29 ),
    .fco(\u2_Display/lt107_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_4|u2_Display/lt107_3  (
    .a({\u2_Display/n3323 ,\u2_Display/n3324 }),
    .b(2'b00),
    .fci(\u2_Display/lt107_c3 ),
    .fco(\u2_Display/lt107_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_6|u2_Display/lt107_5  (
    .a({\u2_Display/n3321 ,\u2_Display/n3322 }),
    .b(2'b10),
    .fci(\u2_Display/lt107_c5 ),
    .fco(\u2_Display/lt107_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_8|u2_Display/lt107_7  (
    .a({\u2_Display/n3319 ,\u2_Display/n3320 }),
    .b(2'b01),
    .fci(\u2_Display/lt107_c7 ),
    .fco(\u2_Display/lt107_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt107_0|u2_Display/lt107_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt107_cout|u2_Display/lt107_31  (
    .a({1'b0,\u2_Display/n3296 }),
    .b(2'b10),
    .fci(\u2_Display/lt107_c31 ),
    .f({\u2_Display/n3328 ,open_n26017}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_0|u2_Display/lt108_cin  (
    .a({\u2_Display/n3362 ,1'b0}),
    .b({1'b0,open_n26023}),
    .fco(\u2_Display/lt108_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_10|u2_Display/lt108_9  (
    .a({\u2_Display/n3352 ,\u2_Display/n3353 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c9 ),
    .fco(\u2_Display/lt108_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_12|u2_Display/lt108_11  (
    .a({\u2_Display/n3350 ,\u2_Display/n3351 }),
    .b(2'b01),
    .fci(\u2_Display/lt108_c11 ),
    .fco(\u2_Display/lt108_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_14|u2_Display/lt108_13  (
    .a({\u2_Display/n3348 ,\u2_Display/n3349 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c13 ),
    .fco(\u2_Display/lt108_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_16|u2_Display/lt108_15  (
    .a({\u2_Display/n3346 ,\u2_Display/n3347 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c15 ),
    .fco(\u2_Display/lt108_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_18|u2_Display/lt108_17  (
    .a({\u2_Display/n3344 ,\u2_Display/n3345 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c17 ),
    .fco(\u2_Display/lt108_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_20|u2_Display/lt108_19  (
    .a({\u2_Display/n3342 ,\u2_Display/n3343 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c19 ),
    .fco(\u2_Display/lt108_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_22|u2_Display/lt108_21  (
    .a({\u2_Display/n3340 ,\u2_Display/n3341 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c21 ),
    .fco(\u2_Display/lt108_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_24|u2_Display/lt108_23  (
    .a({\u2_Display/n3338 ,\u2_Display/n3339 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c23 ),
    .fco(\u2_Display/lt108_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_26|u2_Display/lt108_25  (
    .a({\u2_Display/n3336 ,\u2_Display/n3337 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c25 ),
    .fco(\u2_Display/lt108_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_28|u2_Display/lt108_27  (
    .a({\u2_Display/n3334 ,\u2_Display/n3335 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c27 ),
    .fco(\u2_Display/lt108_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_2|u2_Display/lt108_1  (
    .a({\u2_Display/n3360 ,\u2_Display/n3361 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c1 ),
    .fco(\u2_Display/lt108_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_30|u2_Display/lt108_29  (
    .a({\u2_Display/n3332 ,\u2_Display/n3333 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c29 ),
    .fco(\u2_Display/lt108_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_4|u2_Display/lt108_3  (
    .a({\u2_Display/n3358 ,\u2_Display/n3359 }),
    .b(2'b00),
    .fci(\u2_Display/lt108_c3 ),
    .fco(\u2_Display/lt108_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_6|u2_Display/lt108_5  (
    .a({\u2_Display/n3356 ,\u2_Display/n3357 }),
    .b(2'b11),
    .fci(\u2_Display/lt108_c5 ),
    .fco(\u2_Display/lt108_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_8|u2_Display/lt108_7  (
    .a({\u2_Display/n3354 ,\u2_Display/n3355 }),
    .b(2'b10),
    .fci(\u2_Display/lt108_c7 ),
    .fco(\u2_Display/lt108_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt108_0|u2_Display/lt108_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt108_cout|u2_Display/lt108_31  (
    .a({1'b0,\u2_Display/n3331 }),
    .b(2'b10),
    .fci(\u2_Display/lt108_c31 ),
    .f({\u2_Display/n3363 ,open_n26427}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_0|u2_Display/lt109_cin  (
    .a({\u2_Display/n3397 ,1'b0}),
    .b({1'b0,open_n26433}),
    .fco(\u2_Display/lt109_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_10|u2_Display/lt109_9  (
    .a({\u2_Display/n3387 ,\u2_Display/n3388 }),
    .b(2'b10),
    .fci(\u2_Display/lt109_c9 ),
    .fco(\u2_Display/lt109_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_12|u2_Display/lt109_11  (
    .a({\u2_Display/n3385 ,\u2_Display/n3386 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c11 ),
    .fco(\u2_Display/lt109_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_14|u2_Display/lt109_13  (
    .a({\u2_Display/n3383 ,\u2_Display/n3384 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c13 ),
    .fco(\u2_Display/lt109_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_16|u2_Display/lt109_15  (
    .a({\u2_Display/n3381 ,\u2_Display/n3382 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c15 ),
    .fco(\u2_Display/lt109_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_18|u2_Display/lt109_17  (
    .a({\u2_Display/n3379 ,\u2_Display/n3380 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c17 ),
    .fco(\u2_Display/lt109_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_20|u2_Display/lt109_19  (
    .a({\u2_Display/n3377 ,\u2_Display/n3378 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c19 ),
    .fco(\u2_Display/lt109_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_22|u2_Display/lt109_21  (
    .a({\u2_Display/n3375 ,\u2_Display/n3376 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c21 ),
    .fco(\u2_Display/lt109_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_24|u2_Display/lt109_23  (
    .a({\u2_Display/n3373 ,\u2_Display/n3374 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c23 ),
    .fco(\u2_Display/lt109_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_26|u2_Display/lt109_25  (
    .a({\u2_Display/n3371 ,\u2_Display/n3372 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c25 ),
    .fco(\u2_Display/lt109_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_28|u2_Display/lt109_27  (
    .a({\u2_Display/n3369 ,\u2_Display/n3370 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c27 ),
    .fco(\u2_Display/lt109_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_2|u2_Display/lt109_1  (
    .a({\u2_Display/n3395 ,\u2_Display/n3396 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c1 ),
    .fco(\u2_Display/lt109_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_30|u2_Display/lt109_29  (
    .a({\u2_Display/n3367 ,\u2_Display/n3368 }),
    .b(2'b00),
    .fci(\u2_Display/lt109_c29 ),
    .fco(\u2_Display/lt109_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_4|u2_Display/lt109_3  (
    .a({\u2_Display/n3393 ,\u2_Display/n3394 }),
    .b(2'b10),
    .fci(\u2_Display/lt109_c3 ),
    .fco(\u2_Display/lt109_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_6|u2_Display/lt109_5  (
    .a({\u2_Display/n3391 ,\u2_Display/n3392 }),
    .b(2'b01),
    .fci(\u2_Display/lt109_c5 ),
    .fco(\u2_Display/lt109_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_8|u2_Display/lt109_7  (
    .a({\u2_Display/n3389 ,\u2_Display/n3390 }),
    .b(2'b01),
    .fci(\u2_Display/lt109_c7 ),
    .fco(\u2_Display/lt109_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt109_0|u2_Display/lt109_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt109_cout|u2_Display/lt109_31  (
    .a({1'b0,\u2_Display/n3366 }),
    .b(2'b10),
    .fci(\u2_Display/lt109_c31 ),
    .f({\u2_Display/n3398 ,open_n26837}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_0|u2_Display/lt10_2_cin  (
    .a({lcd_ypos[0],1'b0}),
    .b({\u2_Display/i [0],open_n26843}),
    .fco(\u2_Display/lt10_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_10|u2_Display/lt10_2_9  (
    .a(lcd_ypos[10:9]),
    .b(\u2_Display/n140 [1:0]),
    .fci(\u2_Display/lt10_2_c9 ),
    .fco(\u2_Display/lt10_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_2|u2_Display/lt10_2_1  (
    .a(lcd_ypos[2:1]),
    .b(\u2_Display/i [2:1]),
    .fci(\u2_Display/lt10_2_c1 ),
    .fco(\u2_Display/lt10_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_4|u2_Display/lt10_2_3  (
    .a(lcd_ypos[4:3]),
    .b(\u2_Display/i [4:3]),
    .fci(\u2_Display/lt10_2_c3 ),
    .fco(\u2_Display/lt10_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_6|u2_Display/lt10_2_5  (
    .a(lcd_ypos[6:5]),
    .b(\u2_Display/i [6:5]),
    .fci(\u2_Display/lt10_2_c5 ),
    .fco(\u2_Display/lt10_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_8|u2_Display/lt10_2_7  (
    .a(lcd_ypos[8:7]),
    .b(\u2_Display/i [8:7]),
    .fci(\u2_Display/lt10_2_c7 ),
    .fco(\u2_Display/lt10_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt10_2_0|u2_Display/lt10_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt10_2_cout|u2_Display/lt10_2_11  (
    .a({1'b0,lcd_ypos[11]}),
    .b({1'b1,\u2_Display/add7_2_co }),
    .fci(\u2_Display/lt10_2_c11 ),
    .f({\u2_Display/n141 ,open_n27007}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_0|u2_Display/lt110_cin  (
    .a({\u2_Display/n3432 ,1'b0}),
    .b({1'b0,open_n27013}),
    .fco(\u2_Display/lt110_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_10|u2_Display/lt110_9  (
    .a({\u2_Display/n3422 ,\u2_Display/n3423 }),
    .b(2'b01),
    .fci(\u2_Display/lt110_c9 ),
    .fco(\u2_Display/lt110_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_12|u2_Display/lt110_11  (
    .a({\u2_Display/n3420 ,\u2_Display/n3421 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c11 ),
    .fco(\u2_Display/lt110_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_14|u2_Display/lt110_13  (
    .a({\u2_Display/n3418 ,\u2_Display/n3419 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c13 ),
    .fco(\u2_Display/lt110_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_16|u2_Display/lt110_15  (
    .a({\u2_Display/n3416 ,\u2_Display/n3417 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c15 ),
    .fco(\u2_Display/lt110_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_18|u2_Display/lt110_17  (
    .a({\u2_Display/n3414 ,\u2_Display/n3415 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c17 ),
    .fco(\u2_Display/lt110_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_20|u2_Display/lt110_19  (
    .a({\u2_Display/n3412 ,\u2_Display/n3413 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c19 ),
    .fco(\u2_Display/lt110_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_22|u2_Display/lt110_21  (
    .a({\u2_Display/n3410 ,\u2_Display/n3411 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c21 ),
    .fco(\u2_Display/lt110_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_24|u2_Display/lt110_23  (
    .a({\u2_Display/n3408 ,\u2_Display/n3409 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c23 ),
    .fco(\u2_Display/lt110_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_26|u2_Display/lt110_25  (
    .a({\u2_Display/n3406 ,\u2_Display/n3407 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c25 ),
    .fco(\u2_Display/lt110_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_28|u2_Display/lt110_27  (
    .a({\u2_Display/n3404 ,\u2_Display/n3405 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c27 ),
    .fco(\u2_Display/lt110_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_2|u2_Display/lt110_1  (
    .a({\u2_Display/n3430 ,\u2_Display/n3431 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c1 ),
    .fco(\u2_Display/lt110_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_30|u2_Display/lt110_29  (
    .a({\u2_Display/n3402 ,\u2_Display/n3403 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c29 ),
    .fco(\u2_Display/lt110_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_4|u2_Display/lt110_3  (
    .a({\u2_Display/n3428 ,\u2_Display/n3429 }),
    .b(2'b11),
    .fci(\u2_Display/lt110_c3 ),
    .fco(\u2_Display/lt110_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_6|u2_Display/lt110_5  (
    .a({\u2_Display/n3426 ,\u2_Display/n3427 }),
    .b(2'b10),
    .fci(\u2_Display/lt110_c5 ),
    .fco(\u2_Display/lt110_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_8|u2_Display/lt110_7  (
    .a({\u2_Display/n3424 ,\u2_Display/n3425 }),
    .b(2'b00),
    .fci(\u2_Display/lt110_c7 ),
    .fco(\u2_Display/lt110_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt110_0|u2_Display/lt110_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt110_cout|u2_Display/lt110_31  (
    .a({1'b0,\u2_Display/n3401 }),
    .b(2'b10),
    .fci(\u2_Display/lt110_c31 ),
    .f({\u2_Display/n3433 ,open_n27417}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_0|u2_Display/lt11_2_cin  (
    .a({\u2_Display/n143 [0],1'b0}),
    .b({lcd_ypos[0],open_n27423}),
    .fco(\u2_Display/lt11_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_10|u2_Display/lt11_2_9  (
    .a(\u2_Display/n143 [10:9]),
    .b(lcd_ypos[10:9]),
    .fci(\u2_Display/lt11_2_c9 ),
    .fco(\u2_Display/lt11_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_12|u2_Display/lt11_2_11  (
    .a({\u2_Display/n143 [31],\u2_Display/n143 [31]}),
    .b({1'b0,lcd_ypos[11]}),
    .fci(\u2_Display/lt11_2_c11 ),
    .fco(\u2_Display/lt11_2_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_2|u2_Display/lt11_2_1  (
    .a(\u2_Display/n143 [2:1]),
    .b(lcd_ypos[2:1]),
    .fci(\u2_Display/lt11_2_c1 ),
    .fco(\u2_Display/lt11_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_4|u2_Display/lt11_2_3  (
    .a(\u2_Display/n143 [4:3]),
    .b(lcd_ypos[4:3]),
    .fci(\u2_Display/lt11_2_c3 ),
    .fco(\u2_Display/lt11_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_6|u2_Display/lt11_2_5  (
    .a(\u2_Display/n143 [6:5]),
    .b(lcd_ypos[6:5]),
    .fci(\u2_Display/lt11_2_c5 ),
    .fco(\u2_Display/lt11_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_8|u2_Display/lt11_2_7  (
    .a(\u2_Display/n143 [8:7]),
    .b(lcd_ypos[8:7]),
    .fci(\u2_Display/lt11_2_c7 ),
    .fco(\u2_Display/lt11_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt11_2_0|u2_Display/lt11_2_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt11_2_cout_al_u5060  (
    .a({open_n27593,1'b0}),
    .b({open_n27594,1'b1}),
    .fci(\u2_Display/lt11_2_c13 ),
    .f({open_n27613,\u2_Display/n144 }));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_0|u2_Display/lt121_cin  (
    .a({\u2_Display/counta [0],1'b0}),
    .b({1'b0,open_n27619}),
    .fco(\u2_Display/lt121_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_10|u2_Display/lt121_9  (
    .a(\u2_Display/counta [10:9]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c9 ),
    .fco(\u2_Display/lt121_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_12|u2_Display/lt121_11  (
    .a(\u2_Display/counta [12:11]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c11 ),
    .fco(\u2_Display/lt121_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_14|u2_Display/lt121_13  (
    .a(\u2_Display/counta [14:13]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c13 ),
    .fco(\u2_Display/lt121_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_16|u2_Display/lt121_15  (
    .a(\u2_Display/counta [16:15]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c15 ),
    .fco(\u2_Display/lt121_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_18|u2_Display/lt121_17  (
    .a(\u2_Display/counta [18:17]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c17 ),
    .fco(\u2_Display/lt121_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_20|u2_Display/lt121_19  (
    .a(\u2_Display/counta [20:19]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c19 ),
    .fco(\u2_Display/lt121_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_22|u2_Display/lt121_21  (
    .a(\u2_Display/counta [22:21]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c21 ),
    .fco(\u2_Display/lt121_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_24|u2_Display/lt121_23  (
    .a(\u2_Display/counta [24:23]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c23 ),
    .fco(\u2_Display/lt121_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_26|u2_Display/lt121_25  (
    .a(\u2_Display/counta [26:25]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c25 ),
    .fco(\u2_Display/lt121_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_28|u2_Display/lt121_27  (
    .a(\u2_Display/counta [28:27]),
    .b(2'b01),
    .fci(\u2_Display/lt121_c27 ),
    .fco(\u2_Display/lt121_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_2|u2_Display/lt121_1  (
    .a(\u2_Display/counta [2:1]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c1 ),
    .fco(\u2_Display/lt121_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_30|u2_Display/lt121_29  (
    .a(\u2_Display/counta [30:29]),
    .b(2'b10),
    .fci(\u2_Display/lt121_c29 ),
    .fco(\u2_Display/lt121_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_4|u2_Display/lt121_3  (
    .a(\u2_Display/counta [4:3]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c3 ),
    .fco(\u2_Display/lt121_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_6|u2_Display/lt121_5  (
    .a(\u2_Display/counta [6:5]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c5 ),
    .fco(\u2_Display/lt121_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_8|u2_Display/lt121_7  (
    .a(\u2_Display/counta [8:7]),
    .b(2'b00),
    .fci(\u2_Display/lt121_c7 ),
    .fco(\u2_Display/lt121_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt121_0|u2_Display/lt121_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt121_cout|u2_Display/lt121_31  (
    .a({1'b0,\u2_Display/counta [31]}),
    .b(2'b11),
    .fci(\u2_Display/lt121_c31 ),
    .f({\u2_Display/n3786 ,open_n28023}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_0|u2_Display/lt122_cin  (
    .a({\u2_Display/n3820 ,1'b0}),
    .b({1'b0,open_n28029}),
    .fco(\u2_Display/lt122_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_10|u2_Display/lt122_9  (
    .a({\u2_Display/n3810 ,\u2_Display/n3811 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c9 ),
    .fco(\u2_Display/lt122_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_12|u2_Display/lt122_11  (
    .a({\u2_Display/n3808 ,\u2_Display/n3809 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c11 ),
    .fco(\u2_Display/lt122_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_14|u2_Display/lt122_13  (
    .a({\u2_Display/n3806 ,\u2_Display/n3807 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c13 ),
    .fco(\u2_Display/lt122_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_16|u2_Display/lt122_15  (
    .a({\u2_Display/n3804 ,\u2_Display/n3805 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c15 ),
    .fco(\u2_Display/lt122_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_18|u2_Display/lt122_17  (
    .a({\u2_Display/n3802 ,\u2_Display/n3803 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c17 ),
    .fco(\u2_Display/lt122_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_20|u2_Display/lt122_19  (
    .a({\u2_Display/n3800 ,\u2_Display/n3801 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c19 ),
    .fco(\u2_Display/lt122_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_22|u2_Display/lt122_21  (
    .a({\u2_Display/n3798 ,\u2_Display/n3799 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c21 ),
    .fco(\u2_Display/lt122_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_24|u2_Display/lt122_23  (
    .a({\u2_Display/n3796 ,\u2_Display/n3797 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c23 ),
    .fco(\u2_Display/lt122_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_26|u2_Display/lt122_25  (
    .a({\u2_Display/n3794 ,\u2_Display/n3795 }),
    .b(2'b10),
    .fci(\u2_Display/lt122_c25 ),
    .fco(\u2_Display/lt122_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_28|u2_Display/lt122_27  (
    .a({\u2_Display/n3792 ,\u2_Display/n3793 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c27 ),
    .fco(\u2_Display/lt122_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_2|u2_Display/lt122_1  (
    .a({\u2_Display/n3818 ,\u2_Display/n3819 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c1 ),
    .fco(\u2_Display/lt122_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_30|u2_Display/lt122_29  (
    .a({\u2_Display/n3790 ,\u2_Display/n3791 }),
    .b(2'b11),
    .fci(\u2_Display/lt122_c29 ),
    .fco(\u2_Display/lt122_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_4|u2_Display/lt122_3  (
    .a({\u2_Display/n3816 ,\u2_Display/n3817 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c3 ),
    .fco(\u2_Display/lt122_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_6|u2_Display/lt122_5  (
    .a({\u2_Display/n3814 ,\u2_Display/n3815 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c5 ),
    .fco(\u2_Display/lt122_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_8|u2_Display/lt122_7  (
    .a({\u2_Display/n3812 ,\u2_Display/n3813 }),
    .b(2'b00),
    .fci(\u2_Display/lt122_c7 ),
    .fco(\u2_Display/lt122_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt122_0|u2_Display/lt122_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt122_cout|u2_Display/lt122_31  (
    .a({1'b0,\u2_Display/n3789 }),
    .b(2'b10),
    .fci(\u2_Display/lt122_c31 ),
    .f({\u2_Display/n3821 ,open_n28433}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_0|u2_Display/lt123_cin  (
    .a({\u2_Display/n3855 ,1'b0}),
    .b({1'b0,open_n28439}),
    .fco(\u2_Display/lt123_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_10|u2_Display/lt123_9  (
    .a({\u2_Display/n3845 ,\u2_Display/n3846 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c9 ),
    .fco(\u2_Display/lt123_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_12|u2_Display/lt123_11  (
    .a({\u2_Display/n3843 ,\u2_Display/n3844 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c11 ),
    .fco(\u2_Display/lt123_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_14|u2_Display/lt123_13  (
    .a({\u2_Display/n3841 ,\u2_Display/n3842 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c13 ),
    .fco(\u2_Display/lt123_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_16|u2_Display/lt123_15  (
    .a({\u2_Display/n3839 ,\u2_Display/n3840 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c15 ),
    .fco(\u2_Display/lt123_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_18|u2_Display/lt123_17  (
    .a({\u2_Display/n3837 ,\u2_Display/n3838 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c17 ),
    .fco(\u2_Display/lt123_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_20|u2_Display/lt123_19  (
    .a({\u2_Display/n3835 ,\u2_Display/n3836 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c19 ),
    .fco(\u2_Display/lt123_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_22|u2_Display/lt123_21  (
    .a({\u2_Display/n3833 ,\u2_Display/n3834 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c21 ),
    .fco(\u2_Display/lt123_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_24|u2_Display/lt123_23  (
    .a({\u2_Display/n3831 ,\u2_Display/n3832 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c23 ),
    .fco(\u2_Display/lt123_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_26|u2_Display/lt123_25  (
    .a({\u2_Display/n3829 ,\u2_Display/n3830 }),
    .b(2'b01),
    .fci(\u2_Display/lt123_c25 ),
    .fco(\u2_Display/lt123_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_28|u2_Display/lt123_27  (
    .a({\u2_Display/n3827 ,\u2_Display/n3828 }),
    .b(2'b10),
    .fci(\u2_Display/lt123_c27 ),
    .fco(\u2_Display/lt123_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_2|u2_Display/lt123_1  (
    .a({\u2_Display/n3853 ,\u2_Display/n3854 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c1 ),
    .fco(\u2_Display/lt123_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_30|u2_Display/lt123_29  (
    .a({\u2_Display/n3825 ,\u2_Display/n3826 }),
    .b(2'b01),
    .fci(\u2_Display/lt123_c29 ),
    .fco(\u2_Display/lt123_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_4|u2_Display/lt123_3  (
    .a({\u2_Display/n3851 ,\u2_Display/n3852 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c3 ),
    .fco(\u2_Display/lt123_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_6|u2_Display/lt123_5  (
    .a({\u2_Display/n3849 ,\u2_Display/n3850 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c5 ),
    .fco(\u2_Display/lt123_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_8|u2_Display/lt123_7  (
    .a({\u2_Display/n3847 ,\u2_Display/n3848 }),
    .b(2'b00),
    .fci(\u2_Display/lt123_c7 ),
    .fco(\u2_Display/lt123_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt123_0|u2_Display/lt123_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt123_cout|u2_Display/lt123_31  (
    .a({1'b0,\u2_Display/n3824 }),
    .b(2'b10),
    .fci(\u2_Display/lt123_c31 ),
    .f({\u2_Display/n3856 ,open_n28843}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_0|u2_Display/lt124_cin  (
    .a({\u2_Display/n3890 ,1'b0}),
    .b({1'b0,open_n28849}),
    .fco(\u2_Display/lt124_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_10|u2_Display/lt124_9  (
    .a({\u2_Display/n3880 ,\u2_Display/n3881 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c9 ),
    .fco(\u2_Display/lt124_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_12|u2_Display/lt124_11  (
    .a({\u2_Display/n3878 ,\u2_Display/n3879 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c11 ),
    .fco(\u2_Display/lt124_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_14|u2_Display/lt124_13  (
    .a({\u2_Display/n3876 ,\u2_Display/n3877 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c13 ),
    .fco(\u2_Display/lt124_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_16|u2_Display/lt124_15  (
    .a({\u2_Display/n3874 ,\u2_Display/n3875 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c15 ),
    .fco(\u2_Display/lt124_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_18|u2_Display/lt124_17  (
    .a({\u2_Display/n3872 ,\u2_Display/n3873 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c17 ),
    .fco(\u2_Display/lt124_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_20|u2_Display/lt124_19  (
    .a({\u2_Display/n3870 ,\u2_Display/n3871 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c19 ),
    .fco(\u2_Display/lt124_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_22|u2_Display/lt124_21  (
    .a({\u2_Display/n3868 ,\u2_Display/n3869 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c21 ),
    .fco(\u2_Display/lt124_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_24|u2_Display/lt124_23  (
    .a({\u2_Display/n3866 ,\u2_Display/n3867 }),
    .b(2'b10),
    .fci(\u2_Display/lt124_c23 ),
    .fco(\u2_Display/lt124_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_26|u2_Display/lt124_25  (
    .a({\u2_Display/n3864 ,\u2_Display/n3865 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c25 ),
    .fco(\u2_Display/lt124_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_28|u2_Display/lt124_27  (
    .a({\u2_Display/n3862 ,\u2_Display/n3863 }),
    .b(2'b11),
    .fci(\u2_Display/lt124_c27 ),
    .fco(\u2_Display/lt124_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_2|u2_Display/lt124_1  (
    .a({\u2_Display/n3888 ,\u2_Display/n3889 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c1 ),
    .fco(\u2_Display/lt124_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_30|u2_Display/lt124_29  (
    .a({\u2_Display/n3860 ,\u2_Display/n3861 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c29 ),
    .fco(\u2_Display/lt124_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_4|u2_Display/lt124_3  (
    .a({\u2_Display/n3886 ,\u2_Display/n3887 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c3 ),
    .fco(\u2_Display/lt124_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_6|u2_Display/lt124_5  (
    .a({\u2_Display/n3884 ,\u2_Display/n3885 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c5 ),
    .fco(\u2_Display/lt124_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_8|u2_Display/lt124_7  (
    .a({\u2_Display/n3882 ,\u2_Display/n3883 }),
    .b(2'b00),
    .fci(\u2_Display/lt124_c7 ),
    .fco(\u2_Display/lt124_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt124_0|u2_Display/lt124_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt124_cout|u2_Display/lt124_31  (
    .a({1'b0,\u2_Display/n3859 }),
    .b(2'b10),
    .fci(\u2_Display/lt124_c31 ),
    .f({\u2_Display/n3891 ,open_n29253}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_0|u2_Display/lt125_cin  (
    .a({\u2_Display/n3925 ,1'b0}),
    .b({1'b0,open_n29259}),
    .fco(\u2_Display/lt125_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_10|u2_Display/lt125_9  (
    .a({\u2_Display/n3915 ,\u2_Display/n3916 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c9 ),
    .fco(\u2_Display/lt125_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_12|u2_Display/lt125_11  (
    .a({\u2_Display/n3913 ,\u2_Display/n3914 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c11 ),
    .fco(\u2_Display/lt125_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_14|u2_Display/lt125_13  (
    .a({\u2_Display/n3911 ,\u2_Display/n3912 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c13 ),
    .fco(\u2_Display/lt125_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_16|u2_Display/lt125_15  (
    .a({\u2_Display/n3909 ,\u2_Display/n3910 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c15 ),
    .fco(\u2_Display/lt125_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_18|u2_Display/lt125_17  (
    .a({\u2_Display/n3907 ,\u2_Display/n3908 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c17 ),
    .fco(\u2_Display/lt125_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_20|u2_Display/lt125_19  (
    .a({\u2_Display/n3905 ,\u2_Display/n3906 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c19 ),
    .fco(\u2_Display/lt125_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_22|u2_Display/lt125_21  (
    .a({\u2_Display/n3903 ,\u2_Display/n3904 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c21 ),
    .fco(\u2_Display/lt125_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_24|u2_Display/lt125_23  (
    .a({\u2_Display/n3901 ,\u2_Display/n3902 }),
    .b(2'b01),
    .fci(\u2_Display/lt125_c23 ),
    .fco(\u2_Display/lt125_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_26|u2_Display/lt125_25  (
    .a({\u2_Display/n3899 ,\u2_Display/n3900 }),
    .b(2'b10),
    .fci(\u2_Display/lt125_c25 ),
    .fco(\u2_Display/lt125_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_28|u2_Display/lt125_27  (
    .a({\u2_Display/n3897 ,\u2_Display/n3898 }),
    .b(2'b01),
    .fci(\u2_Display/lt125_c27 ),
    .fco(\u2_Display/lt125_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_2|u2_Display/lt125_1  (
    .a({\u2_Display/n3923 ,\u2_Display/n3924 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c1 ),
    .fco(\u2_Display/lt125_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_30|u2_Display/lt125_29  (
    .a({\u2_Display/n3895 ,\u2_Display/n3896 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c29 ),
    .fco(\u2_Display/lt125_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_4|u2_Display/lt125_3  (
    .a({\u2_Display/n3921 ,\u2_Display/n3922 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c3 ),
    .fco(\u2_Display/lt125_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_6|u2_Display/lt125_5  (
    .a({\u2_Display/n3919 ,\u2_Display/n3920 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c5 ),
    .fco(\u2_Display/lt125_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_8|u2_Display/lt125_7  (
    .a({\u2_Display/n3917 ,\u2_Display/n3918 }),
    .b(2'b00),
    .fci(\u2_Display/lt125_c7 ),
    .fco(\u2_Display/lt125_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt125_0|u2_Display/lt125_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt125_cout|u2_Display/lt125_31  (
    .a({1'b0,\u2_Display/n3894 }),
    .b(2'b10),
    .fci(\u2_Display/lt125_c31 ),
    .f({\u2_Display/n3926 ,open_n29663}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_0|u2_Display/lt126_cin  (
    .a({\u2_Display/n3960 ,1'b0}),
    .b({1'b0,open_n29669}),
    .fco(\u2_Display/lt126_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_10|u2_Display/lt126_9  (
    .a({\u2_Display/n3950 ,\u2_Display/n3951 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c9 ),
    .fco(\u2_Display/lt126_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_12|u2_Display/lt126_11  (
    .a({\u2_Display/n3948 ,\u2_Display/n3949 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c11 ),
    .fco(\u2_Display/lt126_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_14|u2_Display/lt126_13  (
    .a({\u2_Display/n3946 ,\u2_Display/n3947 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c13 ),
    .fco(\u2_Display/lt126_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_16|u2_Display/lt126_15  (
    .a({\u2_Display/n3944 ,\u2_Display/n3945 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c15 ),
    .fco(\u2_Display/lt126_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_18|u2_Display/lt126_17  (
    .a({\u2_Display/n3942 ,\u2_Display/n3943 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c17 ),
    .fco(\u2_Display/lt126_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_20|u2_Display/lt126_19  (
    .a({\u2_Display/n3940 ,\u2_Display/n3941 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c19 ),
    .fco(\u2_Display/lt126_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_22|u2_Display/lt126_21  (
    .a({\u2_Display/n3938 ,\u2_Display/n3939 }),
    .b(2'b10),
    .fci(\u2_Display/lt126_c21 ),
    .fco(\u2_Display/lt126_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_24|u2_Display/lt126_23  (
    .a({\u2_Display/n3936 ,\u2_Display/n3937 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c23 ),
    .fco(\u2_Display/lt126_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_26|u2_Display/lt126_25  (
    .a({\u2_Display/n3934 ,\u2_Display/n3935 }),
    .b(2'b11),
    .fci(\u2_Display/lt126_c25 ),
    .fco(\u2_Display/lt126_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_28|u2_Display/lt126_27  (
    .a({\u2_Display/n3932 ,\u2_Display/n3933 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c27 ),
    .fco(\u2_Display/lt126_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_2|u2_Display/lt126_1  (
    .a({\u2_Display/n3958 ,\u2_Display/n3959 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c1 ),
    .fco(\u2_Display/lt126_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_30|u2_Display/lt126_29  (
    .a({\u2_Display/n3930 ,\u2_Display/n3931 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c29 ),
    .fco(\u2_Display/lt126_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_4|u2_Display/lt126_3  (
    .a({\u2_Display/n3956 ,\u2_Display/n3957 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c3 ),
    .fco(\u2_Display/lt126_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_6|u2_Display/lt126_5  (
    .a({\u2_Display/n3954 ,\u2_Display/n3955 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c5 ),
    .fco(\u2_Display/lt126_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_8|u2_Display/lt126_7  (
    .a({\u2_Display/n3952 ,\u2_Display/n3953 }),
    .b(2'b00),
    .fci(\u2_Display/lt126_c7 ),
    .fco(\u2_Display/lt126_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt126_0|u2_Display/lt126_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt126_cout|u2_Display/lt126_31  (
    .a({1'b0,\u2_Display/n3929 }),
    .b(2'b10),
    .fci(\u2_Display/lt126_c31 ),
    .f({\u2_Display/n3961 ,open_n30073}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_0|u2_Display/lt127_cin  (
    .a({\u2_Display/n3995 ,1'b0}),
    .b({1'b0,open_n30079}),
    .fco(\u2_Display/lt127_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_10|u2_Display/lt127_9  (
    .a({\u2_Display/n3985 ,\u2_Display/n3986 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c9 ),
    .fco(\u2_Display/lt127_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_12|u2_Display/lt127_11  (
    .a({\u2_Display/n3983 ,\u2_Display/n3984 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c11 ),
    .fco(\u2_Display/lt127_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_14|u2_Display/lt127_13  (
    .a({\u2_Display/n3981 ,\u2_Display/n3982 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c13 ),
    .fco(\u2_Display/lt127_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_16|u2_Display/lt127_15  (
    .a({\u2_Display/n3979 ,\u2_Display/n3980 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c15 ),
    .fco(\u2_Display/lt127_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_18|u2_Display/lt127_17  (
    .a({\u2_Display/n3977 ,\u2_Display/n3978 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c17 ),
    .fco(\u2_Display/lt127_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_20|u2_Display/lt127_19  (
    .a({\u2_Display/n3975 ,\u2_Display/n3976 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c19 ),
    .fco(\u2_Display/lt127_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_22|u2_Display/lt127_21  (
    .a({\u2_Display/n3973 ,\u2_Display/n3974 }),
    .b(2'b01),
    .fci(\u2_Display/lt127_c21 ),
    .fco(\u2_Display/lt127_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_24|u2_Display/lt127_23  (
    .a({\u2_Display/n3971 ,\u2_Display/n3972 }),
    .b(2'b10),
    .fci(\u2_Display/lt127_c23 ),
    .fco(\u2_Display/lt127_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_26|u2_Display/lt127_25  (
    .a({\u2_Display/n3969 ,\u2_Display/n3970 }),
    .b(2'b01),
    .fci(\u2_Display/lt127_c25 ),
    .fco(\u2_Display/lt127_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_28|u2_Display/lt127_27  (
    .a({\u2_Display/n3967 ,\u2_Display/n3968 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c27 ),
    .fco(\u2_Display/lt127_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_2|u2_Display/lt127_1  (
    .a({\u2_Display/n3993 ,\u2_Display/n3994 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c1 ),
    .fco(\u2_Display/lt127_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_30|u2_Display/lt127_29  (
    .a({\u2_Display/n3965 ,\u2_Display/n3966 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c29 ),
    .fco(\u2_Display/lt127_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_4|u2_Display/lt127_3  (
    .a({\u2_Display/n3991 ,\u2_Display/n3992 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c3 ),
    .fco(\u2_Display/lt127_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_6|u2_Display/lt127_5  (
    .a({\u2_Display/n3989 ,\u2_Display/n3990 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c5 ),
    .fco(\u2_Display/lt127_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_8|u2_Display/lt127_7  (
    .a({\u2_Display/n3987 ,\u2_Display/n3988 }),
    .b(2'b00),
    .fci(\u2_Display/lt127_c7 ),
    .fco(\u2_Display/lt127_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt127_0|u2_Display/lt127_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt127_cout|u2_Display/lt127_31  (
    .a({1'b0,\u2_Display/n3964 }),
    .b(2'b10),
    .fci(\u2_Display/lt127_c31 ),
    .f({\u2_Display/n3996 ,open_n30483}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_0|u2_Display/lt128_cin  (
    .a({\u2_Display/n4030 ,1'b0}),
    .b({1'b0,open_n30489}),
    .fco(\u2_Display/lt128_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_10|u2_Display/lt128_9  (
    .a({\u2_Display/n4020 ,\u2_Display/n4021 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c9 ),
    .fco(\u2_Display/lt128_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_12|u2_Display/lt128_11  (
    .a({\u2_Display/n4018 ,\u2_Display/n4019 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c11 ),
    .fco(\u2_Display/lt128_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_14|u2_Display/lt128_13  (
    .a({\u2_Display/n4016 ,\u2_Display/n4017 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c13 ),
    .fco(\u2_Display/lt128_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_16|u2_Display/lt128_15  (
    .a({\u2_Display/n4014 ,\u2_Display/n4015 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c15 ),
    .fco(\u2_Display/lt128_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_18|u2_Display/lt128_17  (
    .a({\u2_Display/n4012 ,\u2_Display/n4013 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c17 ),
    .fco(\u2_Display/lt128_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_20|u2_Display/lt128_19  (
    .a({\u2_Display/n4010 ,\u2_Display/n4011 }),
    .b(2'b10),
    .fci(\u2_Display/lt128_c19 ),
    .fco(\u2_Display/lt128_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_22|u2_Display/lt128_21  (
    .a({\u2_Display/n4008 ,\u2_Display/n4009 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c21 ),
    .fco(\u2_Display/lt128_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_24|u2_Display/lt128_23  (
    .a({\u2_Display/n4006 ,\u2_Display/n4007 }),
    .b(2'b11),
    .fci(\u2_Display/lt128_c23 ),
    .fco(\u2_Display/lt128_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_26|u2_Display/lt128_25  (
    .a({\u2_Display/n4004 ,\u2_Display/n4005 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c25 ),
    .fco(\u2_Display/lt128_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_28|u2_Display/lt128_27  (
    .a({\u2_Display/n4002 ,\u2_Display/n4003 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c27 ),
    .fco(\u2_Display/lt128_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_2|u2_Display/lt128_1  (
    .a({\u2_Display/n4028 ,\u2_Display/n4029 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c1 ),
    .fco(\u2_Display/lt128_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_30|u2_Display/lt128_29  (
    .a({\u2_Display/n4000 ,\u2_Display/n4001 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c29 ),
    .fco(\u2_Display/lt128_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_4|u2_Display/lt128_3  (
    .a({\u2_Display/n4026 ,\u2_Display/n4027 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c3 ),
    .fco(\u2_Display/lt128_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_6|u2_Display/lt128_5  (
    .a({\u2_Display/n4024 ,\u2_Display/n4025 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c5 ),
    .fco(\u2_Display/lt128_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_8|u2_Display/lt128_7  (
    .a({\u2_Display/n4022 ,\u2_Display/n4023 }),
    .b(2'b00),
    .fci(\u2_Display/lt128_c7 ),
    .fco(\u2_Display/lt128_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt128_0|u2_Display/lt128_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt128_cout|u2_Display/lt128_31  (
    .a({1'b0,\u2_Display/n3999 }),
    .b(2'b10),
    .fci(\u2_Display/lt128_c31 ),
    .f({\u2_Display/n4031 ,open_n30893}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_0|u2_Display/lt129_cin  (
    .a({\u2_Display/n4065 ,1'b0}),
    .b({1'b0,open_n30899}),
    .fco(\u2_Display/lt129_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_10|u2_Display/lt129_9  (
    .a({\u2_Display/n4055 ,\u2_Display/n4056 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c9 ),
    .fco(\u2_Display/lt129_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_12|u2_Display/lt129_11  (
    .a({\u2_Display/n4053 ,\u2_Display/n4054 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c11 ),
    .fco(\u2_Display/lt129_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_14|u2_Display/lt129_13  (
    .a({\u2_Display/n4051 ,\u2_Display/n4052 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c13 ),
    .fco(\u2_Display/lt129_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_16|u2_Display/lt129_15  (
    .a({\u2_Display/n4049 ,\u2_Display/n4050 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c15 ),
    .fco(\u2_Display/lt129_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_18|u2_Display/lt129_17  (
    .a({\u2_Display/n4047 ,\u2_Display/n4048 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c17 ),
    .fco(\u2_Display/lt129_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_20|u2_Display/lt129_19  (
    .a({\u2_Display/n4045 ,\u2_Display/n4046 }),
    .b(2'b01),
    .fci(\u2_Display/lt129_c19 ),
    .fco(\u2_Display/lt129_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_22|u2_Display/lt129_21  (
    .a({\u2_Display/n4043 ,\u2_Display/n4044 }),
    .b(2'b10),
    .fci(\u2_Display/lt129_c21 ),
    .fco(\u2_Display/lt129_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_24|u2_Display/lt129_23  (
    .a({\u2_Display/n4041 ,\u2_Display/n4042 }),
    .b(2'b01),
    .fci(\u2_Display/lt129_c23 ),
    .fco(\u2_Display/lt129_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_26|u2_Display/lt129_25  (
    .a({\u2_Display/n4039 ,\u2_Display/n4040 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c25 ),
    .fco(\u2_Display/lt129_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_28|u2_Display/lt129_27  (
    .a({\u2_Display/n4037 ,\u2_Display/n4038 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c27 ),
    .fco(\u2_Display/lt129_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_2|u2_Display/lt129_1  (
    .a({\u2_Display/n4063 ,\u2_Display/n4064 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c1 ),
    .fco(\u2_Display/lt129_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_30|u2_Display/lt129_29  (
    .a({\u2_Display/n4035 ,\u2_Display/n4036 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c29 ),
    .fco(\u2_Display/lt129_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_4|u2_Display/lt129_3  (
    .a({\u2_Display/n4061 ,\u2_Display/n4062 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c3 ),
    .fco(\u2_Display/lt129_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_6|u2_Display/lt129_5  (
    .a({\u2_Display/n4059 ,\u2_Display/n4060 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c5 ),
    .fco(\u2_Display/lt129_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_8|u2_Display/lt129_7  (
    .a({\u2_Display/n4057 ,\u2_Display/n4058 }),
    .b(2'b00),
    .fci(\u2_Display/lt129_c7 ),
    .fco(\u2_Display/lt129_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt129_0|u2_Display/lt129_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt129_cout|u2_Display/lt129_31  (
    .a({1'b0,\u2_Display/n4034 }),
    .b(2'b10),
    .fci(\u2_Display/lt129_c31 ),
    .f({\u2_Display/n4066 ,open_n31303}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_0|u2_Display/lt130_cin  (
    .a({\u2_Display/n4100 ,1'b0}),
    .b({1'b0,open_n31309}),
    .fco(\u2_Display/lt130_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_10|u2_Display/lt130_9  (
    .a({\u2_Display/n4090 ,\u2_Display/n4091 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c9 ),
    .fco(\u2_Display/lt130_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_12|u2_Display/lt130_11  (
    .a({\u2_Display/n4088 ,\u2_Display/n4089 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c11 ),
    .fco(\u2_Display/lt130_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_14|u2_Display/lt130_13  (
    .a({\u2_Display/n4086 ,\u2_Display/n4087 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c13 ),
    .fco(\u2_Display/lt130_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_16|u2_Display/lt130_15  (
    .a({\u2_Display/n4084 ,\u2_Display/n4085 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c15 ),
    .fco(\u2_Display/lt130_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_18|u2_Display/lt130_17  (
    .a({\u2_Display/n4082 ,\u2_Display/n4083 }),
    .b(2'b10),
    .fci(\u2_Display/lt130_c17 ),
    .fco(\u2_Display/lt130_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_20|u2_Display/lt130_19  (
    .a({\u2_Display/n4080 ,\u2_Display/n4081 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c19 ),
    .fco(\u2_Display/lt130_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_22|u2_Display/lt130_21  (
    .a({\u2_Display/n4078 ,\u2_Display/n4079 }),
    .b(2'b11),
    .fci(\u2_Display/lt130_c21 ),
    .fco(\u2_Display/lt130_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_24|u2_Display/lt130_23  (
    .a({\u2_Display/n4076 ,\u2_Display/n4077 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c23 ),
    .fco(\u2_Display/lt130_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_26|u2_Display/lt130_25  (
    .a({\u2_Display/n4074 ,\u2_Display/n4075 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c25 ),
    .fco(\u2_Display/lt130_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_28|u2_Display/lt130_27  (
    .a({\u2_Display/n4072 ,\u2_Display/n4073 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c27 ),
    .fco(\u2_Display/lt130_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_2|u2_Display/lt130_1  (
    .a({\u2_Display/n4098 ,\u2_Display/n4099 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c1 ),
    .fco(\u2_Display/lt130_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_30|u2_Display/lt130_29  (
    .a({\u2_Display/n4070 ,\u2_Display/n4071 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c29 ),
    .fco(\u2_Display/lt130_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_4|u2_Display/lt130_3  (
    .a({\u2_Display/n4096 ,\u2_Display/n4097 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c3 ),
    .fco(\u2_Display/lt130_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_6|u2_Display/lt130_5  (
    .a({\u2_Display/n4094 ,\u2_Display/n4095 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c5 ),
    .fco(\u2_Display/lt130_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_8|u2_Display/lt130_7  (
    .a({\u2_Display/n4092 ,\u2_Display/n4093 }),
    .b(2'b00),
    .fci(\u2_Display/lt130_c7 ),
    .fco(\u2_Display/lt130_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt130_0|u2_Display/lt130_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt130_cout|u2_Display/lt130_31  (
    .a({1'b0,\u2_Display/n4069 }),
    .b(2'b10),
    .fci(\u2_Display/lt130_c31 ),
    .f({\u2_Display/n4101 ,open_n31713}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_0|u2_Display/lt131_cin  (
    .a({\u2_Display/n4135 ,1'b0}),
    .b({1'b0,open_n31719}),
    .fco(\u2_Display/lt131_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_10|u2_Display/lt131_9  (
    .a({\u2_Display/n4125 ,\u2_Display/n4126 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c9 ),
    .fco(\u2_Display/lt131_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_12|u2_Display/lt131_11  (
    .a({\u2_Display/n4123 ,\u2_Display/n4124 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c11 ),
    .fco(\u2_Display/lt131_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_14|u2_Display/lt131_13  (
    .a({\u2_Display/n4121 ,\u2_Display/n4122 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c13 ),
    .fco(\u2_Display/lt131_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_16|u2_Display/lt131_15  (
    .a({\u2_Display/n4119 ,\u2_Display/n4120 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c15 ),
    .fco(\u2_Display/lt131_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_18|u2_Display/lt131_17  (
    .a({\u2_Display/n4117 ,\u2_Display/n4118 }),
    .b(2'b01),
    .fci(\u2_Display/lt131_c17 ),
    .fco(\u2_Display/lt131_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_20|u2_Display/lt131_19  (
    .a({\u2_Display/n4115 ,\u2_Display/n4116 }),
    .b(2'b10),
    .fci(\u2_Display/lt131_c19 ),
    .fco(\u2_Display/lt131_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_22|u2_Display/lt131_21  (
    .a({\u2_Display/n4113 ,\u2_Display/n4114 }),
    .b(2'b01),
    .fci(\u2_Display/lt131_c21 ),
    .fco(\u2_Display/lt131_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_24|u2_Display/lt131_23  (
    .a({\u2_Display/n4111 ,\u2_Display/n4112 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c23 ),
    .fco(\u2_Display/lt131_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_26|u2_Display/lt131_25  (
    .a({\u2_Display/n4109 ,\u2_Display/n4110 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c25 ),
    .fco(\u2_Display/lt131_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_28|u2_Display/lt131_27  (
    .a({\u2_Display/n4107 ,\u2_Display/n4108 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c27 ),
    .fco(\u2_Display/lt131_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_2|u2_Display/lt131_1  (
    .a({\u2_Display/n4133 ,\u2_Display/n4134 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c1 ),
    .fco(\u2_Display/lt131_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_30|u2_Display/lt131_29  (
    .a({\u2_Display/n4105 ,\u2_Display/n4106 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c29 ),
    .fco(\u2_Display/lt131_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_4|u2_Display/lt131_3  (
    .a({\u2_Display/n4131 ,\u2_Display/n4132 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c3 ),
    .fco(\u2_Display/lt131_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_6|u2_Display/lt131_5  (
    .a({\u2_Display/n4129 ,\u2_Display/n4130 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c5 ),
    .fco(\u2_Display/lt131_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_8|u2_Display/lt131_7  (
    .a({\u2_Display/n4127 ,\u2_Display/n4128 }),
    .b(2'b00),
    .fci(\u2_Display/lt131_c7 ),
    .fco(\u2_Display/lt131_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt131_0|u2_Display/lt131_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt131_cout|u2_Display/lt131_31  (
    .a({1'b0,\u2_Display/n4104 }),
    .b(2'b10),
    .fci(\u2_Display/lt131_c31 ),
    .f({\u2_Display/n4136 ,open_n32123}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_0|u2_Display/lt132_cin  (
    .a({\u2_Display/n4170 ,1'b0}),
    .b({1'b0,open_n32129}),
    .fco(\u2_Display/lt132_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_10|u2_Display/lt132_9  (
    .a({\u2_Display/n4160 ,\u2_Display/n4161 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c9 ),
    .fco(\u2_Display/lt132_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_12|u2_Display/lt132_11  (
    .a({\u2_Display/n4158 ,\u2_Display/n4159 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c11 ),
    .fco(\u2_Display/lt132_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_14|u2_Display/lt132_13  (
    .a({\u2_Display/n4156 ,\u2_Display/n4157 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c13 ),
    .fco(\u2_Display/lt132_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_16|u2_Display/lt132_15  (
    .a({\u2_Display/n4154 ,\u2_Display/n4155 }),
    .b(2'b10),
    .fci(\u2_Display/lt132_c15 ),
    .fco(\u2_Display/lt132_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_18|u2_Display/lt132_17  (
    .a({\u2_Display/n4152 ,\u2_Display/n4153 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c17 ),
    .fco(\u2_Display/lt132_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_20|u2_Display/lt132_19  (
    .a({\u2_Display/n4150 ,\u2_Display/n4151 }),
    .b(2'b11),
    .fci(\u2_Display/lt132_c19 ),
    .fco(\u2_Display/lt132_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_22|u2_Display/lt132_21  (
    .a({\u2_Display/n4148 ,\u2_Display/n4149 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c21 ),
    .fco(\u2_Display/lt132_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_24|u2_Display/lt132_23  (
    .a({\u2_Display/n4146 ,\u2_Display/n4147 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c23 ),
    .fco(\u2_Display/lt132_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_26|u2_Display/lt132_25  (
    .a({\u2_Display/n4144 ,\u2_Display/n4145 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c25 ),
    .fco(\u2_Display/lt132_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_28|u2_Display/lt132_27  (
    .a({\u2_Display/n4142 ,\u2_Display/n4143 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c27 ),
    .fco(\u2_Display/lt132_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_2|u2_Display/lt132_1  (
    .a({\u2_Display/n4168 ,\u2_Display/n4169 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c1 ),
    .fco(\u2_Display/lt132_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_30|u2_Display/lt132_29  (
    .a({\u2_Display/n4140 ,\u2_Display/n4141 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c29 ),
    .fco(\u2_Display/lt132_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_4|u2_Display/lt132_3  (
    .a({\u2_Display/n4166 ,\u2_Display/n4167 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c3 ),
    .fco(\u2_Display/lt132_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_6|u2_Display/lt132_5  (
    .a({\u2_Display/n4164 ,\u2_Display/n4165 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c5 ),
    .fco(\u2_Display/lt132_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_8|u2_Display/lt132_7  (
    .a({\u2_Display/n4162 ,\u2_Display/n4163 }),
    .b(2'b00),
    .fci(\u2_Display/lt132_c7 ),
    .fco(\u2_Display/lt132_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt132_0|u2_Display/lt132_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt132_cout|u2_Display/lt132_31  (
    .a({1'b0,\u2_Display/n4139 }),
    .b(2'b10),
    .fci(\u2_Display/lt132_c31 ),
    .f({\u2_Display/n4171 ,open_n32533}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_0|u2_Display/lt133_cin  (
    .a({\u2_Display/n4205 ,1'b0}),
    .b({1'b0,open_n32539}),
    .fco(\u2_Display/lt133_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_10|u2_Display/lt133_9  (
    .a({\u2_Display/n4195 ,\u2_Display/n4196 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c9 ),
    .fco(\u2_Display/lt133_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_12|u2_Display/lt133_11  (
    .a({\u2_Display/n4193 ,\u2_Display/n4194 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c11 ),
    .fco(\u2_Display/lt133_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_14|u2_Display/lt133_13  (
    .a({\u2_Display/n4191 ,\u2_Display/n4192 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c13 ),
    .fco(\u2_Display/lt133_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_16|u2_Display/lt133_15  (
    .a({\u2_Display/n4189 ,\u2_Display/n4190 }),
    .b(2'b01),
    .fci(\u2_Display/lt133_c15 ),
    .fco(\u2_Display/lt133_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_18|u2_Display/lt133_17  (
    .a({\u2_Display/n4187 ,\u2_Display/n4188 }),
    .b(2'b10),
    .fci(\u2_Display/lt133_c17 ),
    .fco(\u2_Display/lt133_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_20|u2_Display/lt133_19  (
    .a({\u2_Display/n4185 ,\u2_Display/n4186 }),
    .b(2'b01),
    .fci(\u2_Display/lt133_c19 ),
    .fco(\u2_Display/lt133_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_22|u2_Display/lt133_21  (
    .a({\u2_Display/n4183 ,\u2_Display/n4184 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c21 ),
    .fco(\u2_Display/lt133_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_24|u2_Display/lt133_23  (
    .a({\u2_Display/n4181 ,\u2_Display/n4182 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c23 ),
    .fco(\u2_Display/lt133_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_26|u2_Display/lt133_25  (
    .a({\u2_Display/n4179 ,\u2_Display/n4180 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c25 ),
    .fco(\u2_Display/lt133_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_28|u2_Display/lt133_27  (
    .a({\u2_Display/n4177 ,\u2_Display/n4178 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c27 ),
    .fco(\u2_Display/lt133_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_2|u2_Display/lt133_1  (
    .a({\u2_Display/n4203 ,\u2_Display/n4204 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c1 ),
    .fco(\u2_Display/lt133_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_30|u2_Display/lt133_29  (
    .a({\u2_Display/n4175 ,\u2_Display/n4176 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c29 ),
    .fco(\u2_Display/lt133_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_4|u2_Display/lt133_3  (
    .a({\u2_Display/n4201 ,\u2_Display/n4202 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c3 ),
    .fco(\u2_Display/lt133_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_6|u2_Display/lt133_5  (
    .a({\u2_Display/n4199 ,\u2_Display/n4200 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c5 ),
    .fco(\u2_Display/lt133_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_8|u2_Display/lt133_7  (
    .a({\u2_Display/n4197 ,\u2_Display/n4198 }),
    .b(2'b00),
    .fci(\u2_Display/lt133_c7 ),
    .fco(\u2_Display/lt133_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt133_0|u2_Display/lt133_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt133_cout|u2_Display/lt133_31  (
    .a({1'b0,\u2_Display/n4174 }),
    .b(2'b10),
    .fci(\u2_Display/lt133_c31 ),
    .f({\u2_Display/n4206 ,open_n32943}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_0|u2_Display/lt134_cin  (
    .a({\u2_Display/n4240 ,1'b0}),
    .b({1'b0,open_n32949}),
    .fco(\u2_Display/lt134_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_10|u2_Display/lt134_9  (
    .a({\u2_Display/n4230 ,\u2_Display/n4231 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c9 ),
    .fco(\u2_Display/lt134_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_12|u2_Display/lt134_11  (
    .a({\u2_Display/n4228 ,\u2_Display/n4229 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c11 ),
    .fco(\u2_Display/lt134_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_14|u2_Display/lt134_13  (
    .a({\u2_Display/n4226 ,\u2_Display/n4227 }),
    .b(2'b10),
    .fci(\u2_Display/lt134_c13 ),
    .fco(\u2_Display/lt134_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_16|u2_Display/lt134_15  (
    .a({\u2_Display/n4224 ,\u2_Display/n4225 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c15 ),
    .fco(\u2_Display/lt134_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_18|u2_Display/lt134_17  (
    .a({\u2_Display/n4222 ,\u2_Display/n4223 }),
    .b(2'b11),
    .fci(\u2_Display/lt134_c17 ),
    .fco(\u2_Display/lt134_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_20|u2_Display/lt134_19  (
    .a({\u2_Display/n4220 ,\u2_Display/n4221 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c19 ),
    .fco(\u2_Display/lt134_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_22|u2_Display/lt134_21  (
    .a({\u2_Display/n4218 ,\u2_Display/n4219 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c21 ),
    .fco(\u2_Display/lt134_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_24|u2_Display/lt134_23  (
    .a({\u2_Display/n4216 ,\u2_Display/n4217 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c23 ),
    .fco(\u2_Display/lt134_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_26|u2_Display/lt134_25  (
    .a({\u2_Display/n4214 ,\u2_Display/n4215 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c25 ),
    .fco(\u2_Display/lt134_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_28|u2_Display/lt134_27  (
    .a({\u2_Display/n4212 ,\u2_Display/n4213 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c27 ),
    .fco(\u2_Display/lt134_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_2|u2_Display/lt134_1  (
    .a({\u2_Display/n4238 ,\u2_Display/n4239 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c1 ),
    .fco(\u2_Display/lt134_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_30|u2_Display/lt134_29  (
    .a({\u2_Display/n4210 ,\u2_Display/n4211 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c29 ),
    .fco(\u2_Display/lt134_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_4|u2_Display/lt134_3  (
    .a({\u2_Display/n4236 ,\u2_Display/n4237 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c3 ),
    .fco(\u2_Display/lt134_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_6|u2_Display/lt134_5  (
    .a({\u2_Display/n4234 ,\u2_Display/n4235 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c5 ),
    .fco(\u2_Display/lt134_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_8|u2_Display/lt134_7  (
    .a({\u2_Display/n4232 ,\u2_Display/n4233 }),
    .b(2'b00),
    .fci(\u2_Display/lt134_c7 ),
    .fco(\u2_Display/lt134_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt134_0|u2_Display/lt134_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt134_cout|u2_Display/lt134_31  (
    .a({1'b0,\u2_Display/n4209 }),
    .b(2'b10),
    .fci(\u2_Display/lt134_c31 ),
    .f({\u2_Display/n4241 ,open_n33353}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_0|u2_Display/lt135_cin  (
    .a({\u2_Display/n4275 ,1'b0}),
    .b({1'b0,open_n33359}),
    .fco(\u2_Display/lt135_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_10|u2_Display/lt135_9  (
    .a({\u2_Display/n4265 ,\u2_Display/n4266 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c9 ),
    .fco(\u2_Display/lt135_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_12|u2_Display/lt135_11  (
    .a({\u2_Display/n4263 ,\u2_Display/n4264 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c11 ),
    .fco(\u2_Display/lt135_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_14|u2_Display/lt135_13  (
    .a({\u2_Display/n4261 ,\u2_Display/n4262 }),
    .b(2'b01),
    .fci(\u2_Display/lt135_c13 ),
    .fco(\u2_Display/lt135_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_16|u2_Display/lt135_15  (
    .a({\u2_Display/n4259 ,\u2_Display/n4260 }),
    .b(2'b10),
    .fci(\u2_Display/lt135_c15 ),
    .fco(\u2_Display/lt135_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_18|u2_Display/lt135_17  (
    .a({\u2_Display/n4257 ,\u2_Display/n4258 }),
    .b(2'b01),
    .fci(\u2_Display/lt135_c17 ),
    .fco(\u2_Display/lt135_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_20|u2_Display/lt135_19  (
    .a({\u2_Display/n4255 ,\u2_Display/n4256 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c19 ),
    .fco(\u2_Display/lt135_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_22|u2_Display/lt135_21  (
    .a({\u2_Display/n4253 ,\u2_Display/n4254 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c21 ),
    .fco(\u2_Display/lt135_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_24|u2_Display/lt135_23  (
    .a({\u2_Display/n4251 ,\u2_Display/n4252 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c23 ),
    .fco(\u2_Display/lt135_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_26|u2_Display/lt135_25  (
    .a({\u2_Display/n4249 ,\u2_Display/n4250 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c25 ),
    .fco(\u2_Display/lt135_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_28|u2_Display/lt135_27  (
    .a({\u2_Display/n4247 ,\u2_Display/n4248 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c27 ),
    .fco(\u2_Display/lt135_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_2|u2_Display/lt135_1  (
    .a({\u2_Display/n4273 ,\u2_Display/n4274 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c1 ),
    .fco(\u2_Display/lt135_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_30|u2_Display/lt135_29  (
    .a({\u2_Display/n4245 ,\u2_Display/n4246 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c29 ),
    .fco(\u2_Display/lt135_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_4|u2_Display/lt135_3  (
    .a({\u2_Display/n4271 ,\u2_Display/n4272 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c3 ),
    .fco(\u2_Display/lt135_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_6|u2_Display/lt135_5  (
    .a({\u2_Display/n4269 ,\u2_Display/n4270 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c5 ),
    .fco(\u2_Display/lt135_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_8|u2_Display/lt135_7  (
    .a({\u2_Display/n4267 ,\u2_Display/n4268 }),
    .b(2'b00),
    .fci(\u2_Display/lt135_c7 ),
    .fco(\u2_Display/lt135_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt135_0|u2_Display/lt135_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt135_cout|u2_Display/lt135_31  (
    .a({1'b0,\u2_Display/n4244 }),
    .b(2'b10),
    .fci(\u2_Display/lt135_c31 ),
    .f({\u2_Display/n4276 ,open_n33763}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_0|u2_Display/lt136_cin  (
    .a({\u2_Display/n4310 ,1'b0}),
    .b({1'b0,open_n33769}),
    .fco(\u2_Display/lt136_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_10|u2_Display/lt136_9  (
    .a({\u2_Display/n4300 ,\u2_Display/n4301 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c9 ),
    .fco(\u2_Display/lt136_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_12|u2_Display/lt136_11  (
    .a({\u2_Display/n4298 ,\u2_Display/n4299 }),
    .b(2'b10),
    .fci(\u2_Display/lt136_c11 ),
    .fco(\u2_Display/lt136_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_14|u2_Display/lt136_13  (
    .a({\u2_Display/n4296 ,\u2_Display/n4297 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c13 ),
    .fco(\u2_Display/lt136_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_16|u2_Display/lt136_15  (
    .a({\u2_Display/n4294 ,\u2_Display/n4295 }),
    .b(2'b11),
    .fci(\u2_Display/lt136_c15 ),
    .fco(\u2_Display/lt136_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_18|u2_Display/lt136_17  (
    .a({\u2_Display/n4292 ,\u2_Display/n4293 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c17 ),
    .fco(\u2_Display/lt136_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_20|u2_Display/lt136_19  (
    .a({\u2_Display/n4290 ,\u2_Display/n4291 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c19 ),
    .fco(\u2_Display/lt136_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_22|u2_Display/lt136_21  (
    .a({\u2_Display/n4288 ,\u2_Display/n4289 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c21 ),
    .fco(\u2_Display/lt136_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_24|u2_Display/lt136_23  (
    .a({\u2_Display/n4286 ,\u2_Display/n4287 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c23 ),
    .fco(\u2_Display/lt136_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_26|u2_Display/lt136_25  (
    .a({\u2_Display/n4284 ,\u2_Display/n4285 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c25 ),
    .fco(\u2_Display/lt136_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_28|u2_Display/lt136_27  (
    .a({\u2_Display/n4282 ,\u2_Display/n4283 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c27 ),
    .fco(\u2_Display/lt136_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_2|u2_Display/lt136_1  (
    .a({\u2_Display/n4308 ,\u2_Display/n4309 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c1 ),
    .fco(\u2_Display/lt136_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_30|u2_Display/lt136_29  (
    .a({\u2_Display/n4280 ,\u2_Display/n4281 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c29 ),
    .fco(\u2_Display/lt136_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_4|u2_Display/lt136_3  (
    .a({\u2_Display/n4306 ,\u2_Display/n4307 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c3 ),
    .fco(\u2_Display/lt136_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_6|u2_Display/lt136_5  (
    .a({\u2_Display/n4304 ,\u2_Display/n4305 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c5 ),
    .fco(\u2_Display/lt136_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_8|u2_Display/lt136_7  (
    .a({\u2_Display/n4302 ,\u2_Display/n4303 }),
    .b(2'b00),
    .fci(\u2_Display/lt136_c7 ),
    .fco(\u2_Display/lt136_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt136_0|u2_Display/lt136_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt136_cout|u2_Display/lt136_31  (
    .a({1'b0,\u2_Display/n4279 }),
    .b(2'b10),
    .fci(\u2_Display/lt136_c31 ),
    .f({\u2_Display/n4311 ,open_n34173}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_0|u2_Display/lt137_cin  (
    .a({\u2_Display/n4345 ,1'b0}),
    .b({1'b0,open_n34179}),
    .fco(\u2_Display/lt137_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_10|u2_Display/lt137_9  (
    .a({\u2_Display/n4335 ,\u2_Display/n4336 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c9 ),
    .fco(\u2_Display/lt137_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_12|u2_Display/lt137_11  (
    .a({\u2_Display/n4333 ,\u2_Display/n4334 }),
    .b(2'b01),
    .fci(\u2_Display/lt137_c11 ),
    .fco(\u2_Display/lt137_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_14|u2_Display/lt137_13  (
    .a({\u2_Display/n4331 ,\u2_Display/n4332 }),
    .b(2'b10),
    .fci(\u2_Display/lt137_c13 ),
    .fco(\u2_Display/lt137_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_16|u2_Display/lt137_15  (
    .a({\u2_Display/n4329 ,\u2_Display/n4330 }),
    .b(2'b01),
    .fci(\u2_Display/lt137_c15 ),
    .fco(\u2_Display/lt137_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_18|u2_Display/lt137_17  (
    .a({\u2_Display/n4327 ,\u2_Display/n4328 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c17 ),
    .fco(\u2_Display/lt137_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_20|u2_Display/lt137_19  (
    .a({\u2_Display/n4325 ,\u2_Display/n4326 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c19 ),
    .fco(\u2_Display/lt137_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_22|u2_Display/lt137_21  (
    .a({\u2_Display/n4323 ,\u2_Display/n4324 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c21 ),
    .fco(\u2_Display/lt137_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_24|u2_Display/lt137_23  (
    .a({\u2_Display/n4321 ,\u2_Display/n4322 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c23 ),
    .fco(\u2_Display/lt137_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_26|u2_Display/lt137_25  (
    .a({\u2_Display/n4319 ,\u2_Display/n4320 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c25 ),
    .fco(\u2_Display/lt137_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_28|u2_Display/lt137_27  (
    .a({\u2_Display/n4317 ,\u2_Display/n4318 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c27 ),
    .fco(\u2_Display/lt137_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_2|u2_Display/lt137_1  (
    .a({\u2_Display/n4343 ,\u2_Display/n4344 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c1 ),
    .fco(\u2_Display/lt137_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_30|u2_Display/lt137_29  (
    .a({\u2_Display/n4315 ,\u2_Display/n4316 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c29 ),
    .fco(\u2_Display/lt137_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_4|u2_Display/lt137_3  (
    .a({\u2_Display/n4341 ,\u2_Display/n4342 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c3 ),
    .fco(\u2_Display/lt137_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_6|u2_Display/lt137_5  (
    .a({\u2_Display/n4339 ,\u2_Display/n4340 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c5 ),
    .fco(\u2_Display/lt137_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_8|u2_Display/lt137_7  (
    .a({\u2_Display/n4337 ,\u2_Display/n4338 }),
    .b(2'b00),
    .fci(\u2_Display/lt137_c7 ),
    .fco(\u2_Display/lt137_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt137_0|u2_Display/lt137_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt137_cout|u2_Display/lt137_31  (
    .a({1'b0,\u2_Display/n4314 }),
    .b(2'b10),
    .fci(\u2_Display/lt137_c31 ),
    .f({\u2_Display/n4346 ,open_n34583}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_0|u2_Display/lt138_cin  (
    .a({\u2_Display/n4380 ,1'b0}),
    .b({1'b0,open_n34589}),
    .fco(\u2_Display/lt138_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_10|u2_Display/lt138_9  (
    .a({\u2_Display/n4370 ,\u2_Display/n4371 }),
    .b(2'b10),
    .fci(\u2_Display/lt138_c9 ),
    .fco(\u2_Display/lt138_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_12|u2_Display/lt138_11  (
    .a({\u2_Display/n4368 ,\u2_Display/n4369 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c11 ),
    .fco(\u2_Display/lt138_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_14|u2_Display/lt138_13  (
    .a({\u2_Display/n4366 ,\u2_Display/n4367 }),
    .b(2'b11),
    .fci(\u2_Display/lt138_c13 ),
    .fco(\u2_Display/lt138_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_16|u2_Display/lt138_15  (
    .a({\u2_Display/n4364 ,\u2_Display/n4365 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c15 ),
    .fco(\u2_Display/lt138_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_18|u2_Display/lt138_17  (
    .a({\u2_Display/n4362 ,\u2_Display/n4363 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c17 ),
    .fco(\u2_Display/lt138_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_20|u2_Display/lt138_19  (
    .a({\u2_Display/n4360 ,\u2_Display/n4361 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c19 ),
    .fco(\u2_Display/lt138_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_22|u2_Display/lt138_21  (
    .a({\u2_Display/n4358 ,\u2_Display/n4359 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c21 ),
    .fco(\u2_Display/lt138_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_24|u2_Display/lt138_23  (
    .a({\u2_Display/n4356 ,\u2_Display/n4357 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c23 ),
    .fco(\u2_Display/lt138_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_26|u2_Display/lt138_25  (
    .a({\u2_Display/n4354 ,\u2_Display/n4355 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c25 ),
    .fco(\u2_Display/lt138_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_28|u2_Display/lt138_27  (
    .a({\u2_Display/n4352 ,\u2_Display/n4353 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c27 ),
    .fco(\u2_Display/lt138_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_2|u2_Display/lt138_1  (
    .a({\u2_Display/n4378 ,\u2_Display/n4379 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c1 ),
    .fco(\u2_Display/lt138_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_30|u2_Display/lt138_29  (
    .a({\u2_Display/n4350 ,\u2_Display/n4351 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c29 ),
    .fco(\u2_Display/lt138_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_4|u2_Display/lt138_3  (
    .a({\u2_Display/n4376 ,\u2_Display/n4377 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c3 ),
    .fco(\u2_Display/lt138_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_6|u2_Display/lt138_5  (
    .a({\u2_Display/n4374 ,\u2_Display/n4375 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c5 ),
    .fco(\u2_Display/lt138_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_8|u2_Display/lt138_7  (
    .a({\u2_Display/n4372 ,\u2_Display/n4373 }),
    .b(2'b00),
    .fci(\u2_Display/lt138_c7 ),
    .fco(\u2_Display/lt138_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt138_0|u2_Display/lt138_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt138_cout|u2_Display/lt138_31  (
    .a({1'b0,\u2_Display/n4349 }),
    .b(2'b10),
    .fci(\u2_Display/lt138_c31 ),
    .f({\u2_Display/n4381 ,open_n34993}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_0|u2_Display/lt139_cin  (
    .a({\u2_Display/n4415 ,1'b0}),
    .b({1'b0,open_n34999}),
    .fco(\u2_Display/lt139_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_10|u2_Display/lt139_9  (
    .a({\u2_Display/n4405 ,\u2_Display/n4406 }),
    .b(2'b01),
    .fci(\u2_Display/lt139_c9 ),
    .fco(\u2_Display/lt139_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_12|u2_Display/lt139_11  (
    .a({\u2_Display/n4403 ,\u2_Display/n4404 }),
    .b(2'b10),
    .fci(\u2_Display/lt139_c11 ),
    .fco(\u2_Display/lt139_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_14|u2_Display/lt139_13  (
    .a({\u2_Display/n4401 ,\u2_Display/n4402 }),
    .b(2'b01),
    .fci(\u2_Display/lt139_c13 ),
    .fco(\u2_Display/lt139_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_16|u2_Display/lt139_15  (
    .a({\u2_Display/n4399 ,\u2_Display/n4400 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c15 ),
    .fco(\u2_Display/lt139_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_18|u2_Display/lt139_17  (
    .a({\u2_Display/n4397 ,\u2_Display/n4398 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c17 ),
    .fco(\u2_Display/lt139_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_20|u2_Display/lt139_19  (
    .a({\u2_Display/n4395 ,\u2_Display/n4396 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c19 ),
    .fco(\u2_Display/lt139_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_22|u2_Display/lt139_21  (
    .a({\u2_Display/n4393 ,\u2_Display/n4394 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c21 ),
    .fco(\u2_Display/lt139_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_24|u2_Display/lt139_23  (
    .a({\u2_Display/n4391 ,\u2_Display/n4392 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c23 ),
    .fco(\u2_Display/lt139_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_26|u2_Display/lt139_25  (
    .a({\u2_Display/n4389 ,\u2_Display/n4390 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c25 ),
    .fco(\u2_Display/lt139_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_28|u2_Display/lt139_27  (
    .a({\u2_Display/n4387 ,\u2_Display/n4388 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c27 ),
    .fco(\u2_Display/lt139_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_2|u2_Display/lt139_1  (
    .a({\u2_Display/n4413 ,\u2_Display/n4414 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c1 ),
    .fco(\u2_Display/lt139_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_30|u2_Display/lt139_29  (
    .a({\u2_Display/n4385 ,\u2_Display/n4386 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c29 ),
    .fco(\u2_Display/lt139_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_4|u2_Display/lt139_3  (
    .a({\u2_Display/n4411 ,\u2_Display/n4412 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c3 ),
    .fco(\u2_Display/lt139_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_6|u2_Display/lt139_5  (
    .a({\u2_Display/n4409 ,\u2_Display/n4410 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c5 ),
    .fco(\u2_Display/lt139_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_8|u2_Display/lt139_7  (
    .a({\u2_Display/n4407 ,\u2_Display/n4408 }),
    .b(2'b00),
    .fci(\u2_Display/lt139_c7 ),
    .fco(\u2_Display/lt139_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt139_0|u2_Display/lt139_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt139_cout|u2_Display/lt139_31  (
    .a({1'b0,\u2_Display/n4384 }),
    .b(2'b10),
    .fci(\u2_Display/lt139_c31 ),
    .f({\u2_Display/n4416 ,open_n35403}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_0|u2_Display/lt140_cin  (
    .a({\u2_Display/n4450 ,1'b0}),
    .b({1'b0,open_n35409}),
    .fco(\u2_Display/lt140_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_10|u2_Display/lt140_9  (
    .a({\u2_Display/n4440 ,\u2_Display/n4441 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c9 ),
    .fco(\u2_Display/lt140_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_12|u2_Display/lt140_11  (
    .a({\u2_Display/n4438 ,\u2_Display/n4439 }),
    .b(2'b11),
    .fci(\u2_Display/lt140_c11 ),
    .fco(\u2_Display/lt140_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_14|u2_Display/lt140_13  (
    .a({\u2_Display/n4436 ,\u2_Display/n4437 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c13 ),
    .fco(\u2_Display/lt140_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_16|u2_Display/lt140_15  (
    .a({\u2_Display/n4434 ,\u2_Display/n4435 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c15 ),
    .fco(\u2_Display/lt140_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_18|u2_Display/lt140_17  (
    .a({\u2_Display/n4432 ,\u2_Display/n4433 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c17 ),
    .fco(\u2_Display/lt140_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_20|u2_Display/lt140_19  (
    .a({\u2_Display/n4430 ,\u2_Display/n4431 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c19 ),
    .fco(\u2_Display/lt140_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_22|u2_Display/lt140_21  (
    .a({\u2_Display/n4428 ,\u2_Display/n4429 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c21 ),
    .fco(\u2_Display/lt140_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_24|u2_Display/lt140_23  (
    .a({\u2_Display/n4426 ,\u2_Display/n4427 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c23 ),
    .fco(\u2_Display/lt140_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_26|u2_Display/lt140_25  (
    .a({\u2_Display/n4424 ,\u2_Display/n4425 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c25 ),
    .fco(\u2_Display/lt140_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_28|u2_Display/lt140_27  (
    .a({\u2_Display/n4422 ,\u2_Display/n4423 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c27 ),
    .fco(\u2_Display/lt140_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_2|u2_Display/lt140_1  (
    .a({\u2_Display/n4448 ,\u2_Display/n4449 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c1 ),
    .fco(\u2_Display/lt140_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_30|u2_Display/lt140_29  (
    .a({\u2_Display/n4420 ,\u2_Display/n4421 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c29 ),
    .fco(\u2_Display/lt140_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_4|u2_Display/lt140_3  (
    .a({\u2_Display/n4446 ,\u2_Display/n4447 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c3 ),
    .fco(\u2_Display/lt140_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_6|u2_Display/lt140_5  (
    .a({\u2_Display/n4444 ,\u2_Display/n4445 }),
    .b(2'b00),
    .fci(\u2_Display/lt140_c5 ),
    .fco(\u2_Display/lt140_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_8|u2_Display/lt140_7  (
    .a({\u2_Display/n4442 ,\u2_Display/n4443 }),
    .b(2'b10),
    .fci(\u2_Display/lt140_c7 ),
    .fco(\u2_Display/lt140_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt140_0|u2_Display/lt140_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt140_cout|u2_Display/lt140_31  (
    .a({1'b0,\u2_Display/n4419 }),
    .b(2'b10),
    .fci(\u2_Display/lt140_c31 ),
    .f({\u2_Display/n4451 ,open_n35813}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_0|u2_Display/lt141_cin  (
    .a({\u2_Display/n4485 ,1'b0}),
    .b({1'b0,open_n35819}),
    .fco(\u2_Display/lt141_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_10|u2_Display/lt141_9  (
    .a({\u2_Display/n4475 ,\u2_Display/n4476 }),
    .b(2'b10),
    .fci(\u2_Display/lt141_c9 ),
    .fco(\u2_Display/lt141_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_12|u2_Display/lt141_11  (
    .a({\u2_Display/n4473 ,\u2_Display/n4474 }),
    .b(2'b01),
    .fci(\u2_Display/lt141_c11 ),
    .fco(\u2_Display/lt141_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_14|u2_Display/lt141_13  (
    .a({\u2_Display/n4471 ,\u2_Display/n4472 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c13 ),
    .fco(\u2_Display/lt141_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_16|u2_Display/lt141_15  (
    .a({\u2_Display/n4469 ,\u2_Display/n4470 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c15 ),
    .fco(\u2_Display/lt141_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_18|u2_Display/lt141_17  (
    .a({\u2_Display/n4467 ,\u2_Display/n4468 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c17 ),
    .fco(\u2_Display/lt141_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_20|u2_Display/lt141_19  (
    .a({\u2_Display/n4465 ,\u2_Display/n4466 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c19 ),
    .fco(\u2_Display/lt141_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_22|u2_Display/lt141_21  (
    .a({\u2_Display/n4463 ,\u2_Display/n4464 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c21 ),
    .fco(\u2_Display/lt141_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_24|u2_Display/lt141_23  (
    .a({\u2_Display/n4461 ,\u2_Display/n4462 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c23 ),
    .fco(\u2_Display/lt141_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_26|u2_Display/lt141_25  (
    .a({\u2_Display/n4459 ,\u2_Display/n4460 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c25 ),
    .fco(\u2_Display/lt141_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_28|u2_Display/lt141_27  (
    .a({\u2_Display/n4457 ,\u2_Display/n4458 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c27 ),
    .fco(\u2_Display/lt141_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_2|u2_Display/lt141_1  (
    .a({\u2_Display/n4483 ,\u2_Display/n4484 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c1 ),
    .fco(\u2_Display/lt141_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_30|u2_Display/lt141_29  (
    .a({\u2_Display/n4455 ,\u2_Display/n4456 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c29 ),
    .fco(\u2_Display/lt141_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_4|u2_Display/lt141_3  (
    .a({\u2_Display/n4481 ,\u2_Display/n4482 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c3 ),
    .fco(\u2_Display/lt141_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_6|u2_Display/lt141_5  (
    .a({\u2_Display/n4479 ,\u2_Display/n4480 }),
    .b(2'b00),
    .fci(\u2_Display/lt141_c5 ),
    .fco(\u2_Display/lt141_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_8|u2_Display/lt141_7  (
    .a({\u2_Display/n4477 ,\u2_Display/n4478 }),
    .b(2'b01),
    .fci(\u2_Display/lt141_c7 ),
    .fco(\u2_Display/lt141_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt141_0|u2_Display/lt141_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt141_cout|u2_Display/lt141_31  (
    .a({1'b0,\u2_Display/n4454 }),
    .b(2'b10),
    .fci(\u2_Display/lt141_c31 ),
    .f({\u2_Display/n4486 ,open_n36223}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_0|u2_Display/lt142_cin  (
    .a({\u2_Display/n4520 ,1'b0}),
    .b({1'b0,open_n36229}),
    .fco(\u2_Display/lt142_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_10|u2_Display/lt142_9  (
    .a({\u2_Display/n4510 ,\u2_Display/n4511 }),
    .b(2'b11),
    .fci(\u2_Display/lt142_c9 ),
    .fco(\u2_Display/lt142_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_12|u2_Display/lt142_11  (
    .a({\u2_Display/n4508 ,\u2_Display/n4509 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c11 ),
    .fco(\u2_Display/lt142_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_14|u2_Display/lt142_13  (
    .a({\u2_Display/n4506 ,\u2_Display/n4507 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c13 ),
    .fco(\u2_Display/lt142_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_16|u2_Display/lt142_15  (
    .a({\u2_Display/n4504 ,\u2_Display/n4505 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c15 ),
    .fco(\u2_Display/lt142_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_18|u2_Display/lt142_17  (
    .a({\u2_Display/n4502 ,\u2_Display/n4503 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c17 ),
    .fco(\u2_Display/lt142_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_20|u2_Display/lt142_19  (
    .a({\u2_Display/n4500 ,\u2_Display/n4501 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c19 ),
    .fco(\u2_Display/lt142_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_22|u2_Display/lt142_21  (
    .a({\u2_Display/n4498 ,\u2_Display/n4499 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c21 ),
    .fco(\u2_Display/lt142_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_24|u2_Display/lt142_23  (
    .a({\u2_Display/n4496 ,\u2_Display/n4497 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c23 ),
    .fco(\u2_Display/lt142_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_26|u2_Display/lt142_25  (
    .a({\u2_Display/n4494 ,\u2_Display/n4495 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c25 ),
    .fco(\u2_Display/lt142_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_28|u2_Display/lt142_27  (
    .a({\u2_Display/n4492 ,\u2_Display/n4493 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c27 ),
    .fco(\u2_Display/lt142_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_2|u2_Display/lt142_1  (
    .a({\u2_Display/n4518 ,\u2_Display/n4519 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c1 ),
    .fco(\u2_Display/lt142_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_30|u2_Display/lt142_29  (
    .a({\u2_Display/n4490 ,\u2_Display/n4491 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c29 ),
    .fco(\u2_Display/lt142_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_4|u2_Display/lt142_3  (
    .a({\u2_Display/n4516 ,\u2_Display/n4517 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c3 ),
    .fco(\u2_Display/lt142_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_6|u2_Display/lt142_5  (
    .a({\u2_Display/n4514 ,\u2_Display/n4515 }),
    .b(2'b10),
    .fci(\u2_Display/lt142_c5 ),
    .fco(\u2_Display/lt142_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_8|u2_Display/lt142_7  (
    .a({\u2_Display/n4512 ,\u2_Display/n4513 }),
    .b(2'b00),
    .fci(\u2_Display/lt142_c7 ),
    .fco(\u2_Display/lt142_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt142_0|u2_Display/lt142_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt142_cout|u2_Display/lt142_31  (
    .a({1'b0,\u2_Display/n4489 }),
    .b(2'b10),
    .fci(\u2_Display/lt142_c31 ),
    .f({\u2_Display/n4521 ,open_n36633}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_0|u2_Display/lt143_cin  (
    .a({\u2_Display/n4555 ,1'b0}),
    .b({1'b0,open_n36639}),
    .fco(\u2_Display/lt143_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_10|u2_Display/lt143_9  (
    .a({\u2_Display/n4545 ,\u2_Display/n4546 }),
    .b(2'b01),
    .fci(\u2_Display/lt143_c9 ),
    .fco(\u2_Display/lt143_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_12|u2_Display/lt143_11  (
    .a({\u2_Display/n4543 ,\u2_Display/n4544 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c11 ),
    .fco(\u2_Display/lt143_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_14|u2_Display/lt143_13  (
    .a({\u2_Display/n4541 ,\u2_Display/n4542 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c13 ),
    .fco(\u2_Display/lt143_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_16|u2_Display/lt143_15  (
    .a({\u2_Display/n4539 ,\u2_Display/n4540 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c15 ),
    .fco(\u2_Display/lt143_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_18|u2_Display/lt143_17  (
    .a({\u2_Display/n4537 ,\u2_Display/n4538 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c17 ),
    .fco(\u2_Display/lt143_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_20|u2_Display/lt143_19  (
    .a({\u2_Display/n4535 ,\u2_Display/n4536 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c19 ),
    .fco(\u2_Display/lt143_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_22|u2_Display/lt143_21  (
    .a({\u2_Display/n4533 ,\u2_Display/n4534 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c21 ),
    .fco(\u2_Display/lt143_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_24|u2_Display/lt143_23  (
    .a({\u2_Display/n4531 ,\u2_Display/n4532 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c23 ),
    .fco(\u2_Display/lt143_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_26|u2_Display/lt143_25  (
    .a({\u2_Display/n4529 ,\u2_Display/n4530 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c25 ),
    .fco(\u2_Display/lt143_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_28|u2_Display/lt143_27  (
    .a({\u2_Display/n4527 ,\u2_Display/n4528 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c27 ),
    .fco(\u2_Display/lt143_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_2|u2_Display/lt143_1  (
    .a({\u2_Display/n4553 ,\u2_Display/n4554 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c1 ),
    .fco(\u2_Display/lt143_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_30|u2_Display/lt143_29  (
    .a({\u2_Display/n4525 ,\u2_Display/n4526 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c29 ),
    .fco(\u2_Display/lt143_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_4|u2_Display/lt143_3  (
    .a({\u2_Display/n4551 ,\u2_Display/n4552 }),
    .b(2'b00),
    .fci(\u2_Display/lt143_c3 ),
    .fco(\u2_Display/lt143_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_6|u2_Display/lt143_5  (
    .a({\u2_Display/n4549 ,\u2_Display/n4550 }),
    .b(2'b01),
    .fci(\u2_Display/lt143_c5 ),
    .fco(\u2_Display/lt143_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_8|u2_Display/lt143_7  (
    .a({\u2_Display/n4547 ,\u2_Display/n4548 }),
    .b(2'b10),
    .fci(\u2_Display/lt143_c7 ),
    .fco(\u2_Display/lt143_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt143_0|u2_Display/lt143_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt143_cout|u2_Display/lt143_31  (
    .a({1'b0,\u2_Display/n4524 }),
    .b(2'b10),
    .fci(\u2_Display/lt143_c31 ),
    .f({\u2_Display/n4556 ,open_n37043}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_0|u2_Display/lt154_cin  (
    .a({\u2_Display/counta [0],1'b0}),
    .b({1'b0,open_n37049}),
    .fco(\u2_Display/lt154_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_10|u2_Display/lt154_9  (
    .a(\u2_Display/counta [10:9]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c9 ),
    .fco(\u2_Display/lt154_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_12|u2_Display/lt154_11  (
    .a(\u2_Display/counta [12:11]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c11 ),
    .fco(\u2_Display/lt154_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_14|u2_Display/lt154_13  (
    .a(\u2_Display/counta [14:13]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c13 ),
    .fco(\u2_Display/lt154_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_16|u2_Display/lt154_15  (
    .a(\u2_Display/counta [16:15]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c15 ),
    .fco(\u2_Display/lt154_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_18|u2_Display/lt154_17  (
    .a(\u2_Display/counta [18:17]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c17 ),
    .fco(\u2_Display/lt154_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_20|u2_Display/lt154_19  (
    .a(\u2_Display/counta [20:19]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c19 ),
    .fco(\u2_Display/lt154_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_22|u2_Display/lt154_21  (
    .a(\u2_Display/counta [22:21]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c21 ),
    .fco(\u2_Display/lt154_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_24|u2_Display/lt154_23  (
    .a(\u2_Display/counta [24:23]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c23 ),
    .fco(\u2_Display/lt154_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_26|u2_Display/lt154_25  (
    .a(\u2_Display/counta [26:25]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c25 ),
    .fco(\u2_Display/lt154_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_28|u2_Display/lt154_27  (
    .a(\u2_Display/counta [28:27]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c27 ),
    .fco(\u2_Display/lt154_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_2|u2_Display/lt154_1  (
    .a(\u2_Display/counta [2:1]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c1 ),
    .fco(\u2_Display/lt154_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_30|u2_Display/lt154_29  (
    .a(\u2_Display/counta [30:29]),
    .b(2'b01),
    .fci(\u2_Display/lt154_c29 ),
    .fco(\u2_Display/lt154_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_4|u2_Display/lt154_3  (
    .a(\u2_Display/counta [4:3]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c3 ),
    .fco(\u2_Display/lt154_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_6|u2_Display/lt154_5  (
    .a(\u2_Display/counta [6:5]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c5 ),
    .fco(\u2_Display/lt154_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_8|u2_Display/lt154_7  (
    .a(\u2_Display/counta [8:7]),
    .b(2'b00),
    .fci(\u2_Display/lt154_c7 ),
    .fco(\u2_Display/lt154_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt154_0|u2_Display/lt154_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt154_cout|u2_Display/lt154_31  (
    .a({1'b0,\u2_Display/counta [31]}),
    .b(2'b11),
    .fci(\u2_Display/lt154_c31 ),
    .f({\u2_Display/n4909 ,open_n37453}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_0|u2_Display/lt155_cin  (
    .a({\u2_Display/n6101 ,1'b0}),
    .b({1'b0,open_n37459}),
    .fco(\u2_Display/lt155_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_10|u2_Display/lt155_9  (
    .a({\u2_Display/n6091 ,\u2_Display/n6092 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c9 ),
    .fco(\u2_Display/lt155_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_12|u2_Display/lt155_11  (
    .a({\u2_Display/n6089 ,\u2_Display/n6090 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c11 ),
    .fco(\u2_Display/lt155_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_14|u2_Display/lt155_13  (
    .a({\u2_Display/n6087 ,\u2_Display/n6088 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c13 ),
    .fco(\u2_Display/lt155_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_16|u2_Display/lt155_15  (
    .a({\u2_Display/n6085 ,\u2_Display/n6086 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c15 ),
    .fco(\u2_Display/lt155_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_18|u2_Display/lt155_17  (
    .a({\u2_Display/n6083 ,\u2_Display/n6084 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c17 ),
    .fco(\u2_Display/lt155_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_20|u2_Display/lt155_19  (
    .a({\u2_Display/n6081 ,\u2_Display/n6082 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c19 ),
    .fco(\u2_Display/lt155_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_22|u2_Display/lt155_21  (
    .a({\u2_Display/n6079 ,\u2_Display/n6080 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c21 ),
    .fco(\u2_Display/lt155_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_24|u2_Display/lt155_23  (
    .a({\u2_Display/n6077 ,\u2_Display/n6078 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c23 ),
    .fco(\u2_Display/lt155_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_26|u2_Display/lt155_25  (
    .a({\u2_Display/n6075 ,\u2_Display/n6076 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c25 ),
    .fco(\u2_Display/lt155_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_28|u2_Display/lt155_27  (
    .a({\u2_Display/n6073 ,\u2_Display/n6074 }),
    .b(2'b10),
    .fci(\u2_Display/lt155_c27 ),
    .fco(\u2_Display/lt155_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_2|u2_Display/lt155_1  (
    .a({\u2_Display/n6099 ,\u2_Display/n6100 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c1 ),
    .fco(\u2_Display/lt155_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_30|u2_Display/lt155_29  (
    .a({\u2_Display/n6071 ,\u2_Display/n6072 }),
    .b(2'b10),
    .fci(\u2_Display/lt155_c29 ),
    .fco(\u2_Display/lt155_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_4|u2_Display/lt155_3  (
    .a({\u2_Display/n6097 ,\u2_Display/n6098 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c3 ),
    .fco(\u2_Display/lt155_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_6|u2_Display/lt155_5  (
    .a({\u2_Display/n6095 ,\u2_Display/n6096 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c5 ),
    .fco(\u2_Display/lt155_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_8|u2_Display/lt155_7  (
    .a({\u2_Display/n6093 ,\u2_Display/n6094 }),
    .b(2'b00),
    .fci(\u2_Display/lt155_c7 ),
    .fco(\u2_Display/lt155_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt155_0|u2_Display/lt155_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt155_cout|u2_Display/lt155_31  (
    .a({1'b0,\u2_Display/n6070 }),
    .b(2'b10),
    .fci(\u2_Display/lt155_c31 ),
    .f({\u2_Display/n4944 ,open_n37863}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_0|u2_Display/lt156_cin  (
    .a({\u2_Display/n6136 ,1'b0}),
    .b({1'b0,open_n37869}),
    .fco(\u2_Display/lt156_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_10|u2_Display/lt156_9  (
    .a({\u2_Display/n6126 ,\u2_Display/n6127 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c9 ),
    .fco(\u2_Display/lt156_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_12|u2_Display/lt156_11  (
    .a({\u2_Display/n6124 ,\u2_Display/n6125 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c11 ),
    .fco(\u2_Display/lt156_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_14|u2_Display/lt156_13  (
    .a({\u2_Display/n6122 ,\u2_Display/n6123 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c13 ),
    .fco(\u2_Display/lt156_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_16|u2_Display/lt156_15  (
    .a({\u2_Display/n6120 ,\u2_Display/n6121 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c15 ),
    .fco(\u2_Display/lt156_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_18|u2_Display/lt156_17  (
    .a({\u2_Display/n6118 ,\u2_Display/n6119 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c17 ),
    .fco(\u2_Display/lt156_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_20|u2_Display/lt156_19  (
    .a({\u2_Display/n6116 ,\u2_Display/n6117 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c19 ),
    .fco(\u2_Display/lt156_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_22|u2_Display/lt156_21  (
    .a({\u2_Display/n6114 ,\u2_Display/n6115 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c21 ),
    .fco(\u2_Display/lt156_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_24|u2_Display/lt156_23  (
    .a({\u2_Display/n6112 ,\u2_Display/n6113 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c23 ),
    .fco(\u2_Display/lt156_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_26|u2_Display/lt156_25  (
    .a({\u2_Display/n6110 ,\u2_Display/n6111 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c25 ),
    .fco(\u2_Display/lt156_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_28|u2_Display/lt156_27  (
    .a({\u2_Display/n6108 ,\u2_Display/n6109 }),
    .b(2'b01),
    .fci(\u2_Display/lt156_c27 ),
    .fco(\u2_Display/lt156_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_2|u2_Display/lt156_1  (
    .a({\u2_Display/n6134 ,\u2_Display/n6135 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c1 ),
    .fco(\u2_Display/lt156_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_30|u2_Display/lt156_29  (
    .a({\u2_Display/n6106 ,\u2_Display/n6107 }),
    .b(2'b01),
    .fci(\u2_Display/lt156_c29 ),
    .fco(\u2_Display/lt156_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_4|u2_Display/lt156_3  (
    .a({\u2_Display/n6132 ,\u2_Display/n6133 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c3 ),
    .fco(\u2_Display/lt156_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_6|u2_Display/lt156_5  (
    .a({\u2_Display/n6130 ,\u2_Display/n6131 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c5 ),
    .fco(\u2_Display/lt156_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_8|u2_Display/lt156_7  (
    .a({\u2_Display/n6128 ,\u2_Display/n6129 }),
    .b(2'b00),
    .fci(\u2_Display/lt156_c7 ),
    .fco(\u2_Display/lt156_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt156_0|u2_Display/lt156_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt156_cout|u2_Display/lt156_31  (
    .a({1'b0,\u2_Display/n6105 }),
    .b(2'b10),
    .fci(\u2_Display/lt156_c31 ),
    .f({\u2_Display/n4979 ,open_n38273}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_0|u2_Display/lt157_cin  (
    .a({\u2_Display/n6171 ,1'b0}),
    .b({1'b0,open_n38279}),
    .fco(\u2_Display/lt157_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_10|u2_Display/lt157_9  (
    .a({\u2_Display/n6161 ,\u2_Display/n6162 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c9 ),
    .fco(\u2_Display/lt157_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_12|u2_Display/lt157_11  (
    .a({\u2_Display/n6159 ,\u2_Display/n6160 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c11 ),
    .fco(\u2_Display/lt157_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_14|u2_Display/lt157_13  (
    .a({\u2_Display/n6157 ,\u2_Display/n6158 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c13 ),
    .fco(\u2_Display/lt157_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_16|u2_Display/lt157_15  (
    .a({\u2_Display/n6155 ,\u2_Display/n6156 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c15 ),
    .fco(\u2_Display/lt157_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_18|u2_Display/lt157_17  (
    .a({\u2_Display/n6153 ,\u2_Display/n6154 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c17 ),
    .fco(\u2_Display/lt157_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_20|u2_Display/lt157_19  (
    .a({\u2_Display/n6151 ,\u2_Display/n6152 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c19 ),
    .fco(\u2_Display/lt157_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_22|u2_Display/lt157_21  (
    .a({\u2_Display/n6149 ,\u2_Display/n6150 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c21 ),
    .fco(\u2_Display/lt157_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_24|u2_Display/lt157_23  (
    .a({\u2_Display/n6147 ,\u2_Display/n6148 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c23 ),
    .fco(\u2_Display/lt157_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_26|u2_Display/lt157_25  (
    .a({\u2_Display/n6145 ,\u2_Display/n6146 }),
    .b(2'b10),
    .fci(\u2_Display/lt157_c25 ),
    .fco(\u2_Display/lt157_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_28|u2_Display/lt157_27  (
    .a({\u2_Display/n6143 ,\u2_Display/n6144 }),
    .b(2'b10),
    .fci(\u2_Display/lt157_c27 ),
    .fco(\u2_Display/lt157_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_2|u2_Display/lt157_1  (
    .a({\u2_Display/n6169 ,\u2_Display/n6170 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c1 ),
    .fco(\u2_Display/lt157_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_30|u2_Display/lt157_29  (
    .a({\u2_Display/n6141 ,\u2_Display/n6142 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c29 ),
    .fco(\u2_Display/lt157_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_4|u2_Display/lt157_3  (
    .a({\u2_Display/n6167 ,\u2_Display/n6168 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c3 ),
    .fco(\u2_Display/lt157_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_6|u2_Display/lt157_5  (
    .a({\u2_Display/n6165 ,\u2_Display/n6166 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c5 ),
    .fco(\u2_Display/lt157_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_8|u2_Display/lt157_7  (
    .a({\u2_Display/n6163 ,\u2_Display/n6164 }),
    .b(2'b00),
    .fci(\u2_Display/lt157_c7 ),
    .fco(\u2_Display/lt157_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt157_0|u2_Display/lt157_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt157_cout|u2_Display/lt157_31  (
    .a({1'b0,\u2_Display/n6140 }),
    .b(2'b10),
    .fci(\u2_Display/lt157_c31 ),
    .f({\u2_Display/n5014 ,open_n38683}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_0|u2_Display/lt158_cin  (
    .a({\u2_Display/n6206 ,1'b0}),
    .b({1'b0,open_n38689}),
    .fco(\u2_Display/lt158_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_10|u2_Display/lt158_9  (
    .a({\u2_Display/n6196 ,\u2_Display/n6197 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c9 ),
    .fco(\u2_Display/lt158_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_12|u2_Display/lt158_11  (
    .a({\u2_Display/n6194 ,\u2_Display/n6195 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c11 ),
    .fco(\u2_Display/lt158_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_14|u2_Display/lt158_13  (
    .a({\u2_Display/n6192 ,\u2_Display/n6193 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c13 ),
    .fco(\u2_Display/lt158_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_16|u2_Display/lt158_15  (
    .a({\u2_Display/n6190 ,\u2_Display/n6191 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c15 ),
    .fco(\u2_Display/lt158_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_18|u2_Display/lt158_17  (
    .a({\u2_Display/n6188 ,\u2_Display/n6189 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c17 ),
    .fco(\u2_Display/lt158_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_20|u2_Display/lt158_19  (
    .a({\u2_Display/n6186 ,\u2_Display/n6187 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c19 ),
    .fco(\u2_Display/lt158_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_22|u2_Display/lt158_21  (
    .a({\u2_Display/n6184 ,\u2_Display/n6185 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c21 ),
    .fco(\u2_Display/lt158_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_24|u2_Display/lt158_23  (
    .a({\u2_Display/n6182 ,\u2_Display/n6183 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c23 ),
    .fco(\u2_Display/lt158_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_26|u2_Display/lt158_25  (
    .a({\u2_Display/n6180 ,\u2_Display/n6181 }),
    .b(2'b01),
    .fci(\u2_Display/lt158_c25 ),
    .fco(\u2_Display/lt158_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_28|u2_Display/lt158_27  (
    .a({\u2_Display/n6178 ,\u2_Display/n6179 }),
    .b(2'b01),
    .fci(\u2_Display/lt158_c27 ),
    .fco(\u2_Display/lt158_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_2|u2_Display/lt158_1  (
    .a({\u2_Display/n6204 ,\u2_Display/n6205 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c1 ),
    .fco(\u2_Display/lt158_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_30|u2_Display/lt158_29  (
    .a({\u2_Display/n6176 ,\u2_Display/n6177 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c29 ),
    .fco(\u2_Display/lt158_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_4|u2_Display/lt158_3  (
    .a({\u2_Display/n6202 ,\u2_Display/n6203 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c3 ),
    .fco(\u2_Display/lt158_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_6|u2_Display/lt158_5  (
    .a({\u2_Display/n6200 ,\u2_Display/n6201 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c5 ),
    .fco(\u2_Display/lt158_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_8|u2_Display/lt158_7  (
    .a({\u2_Display/n6198 ,\u2_Display/n6199 }),
    .b(2'b00),
    .fci(\u2_Display/lt158_c7 ),
    .fco(\u2_Display/lt158_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt158_0|u2_Display/lt158_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt158_cout|u2_Display/lt158_31  (
    .a({1'b0,\u2_Display/n6175 }),
    .b(2'b10),
    .fci(\u2_Display/lt158_c31 ),
    .f({\u2_Display/n5049 ,open_n39093}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_0|u2_Display/lt159_cin  (
    .a({\u2_Display/n6241 ,1'b0}),
    .b({1'b0,open_n39099}),
    .fco(\u2_Display/lt159_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_10|u2_Display/lt159_9  (
    .a({\u2_Display/n6231 ,\u2_Display/n6232 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c9 ),
    .fco(\u2_Display/lt159_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_12|u2_Display/lt159_11  (
    .a({\u2_Display/n6229 ,\u2_Display/n6230 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c11 ),
    .fco(\u2_Display/lt159_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_14|u2_Display/lt159_13  (
    .a({\u2_Display/n6227 ,\u2_Display/n6228 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c13 ),
    .fco(\u2_Display/lt159_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_16|u2_Display/lt159_15  (
    .a({\u2_Display/n6225 ,\u2_Display/n6226 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c15 ),
    .fco(\u2_Display/lt159_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_18|u2_Display/lt159_17  (
    .a({\u2_Display/n6223 ,\u2_Display/n6224 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c17 ),
    .fco(\u2_Display/lt159_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_20|u2_Display/lt159_19  (
    .a({\u2_Display/n6221 ,\u2_Display/n6222 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c19 ),
    .fco(\u2_Display/lt159_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_22|u2_Display/lt159_21  (
    .a({\u2_Display/n6219 ,\u2_Display/n6220 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c21 ),
    .fco(\u2_Display/lt159_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_24|u2_Display/lt159_23  (
    .a({\u2_Display/n6217 ,\u2_Display/n6218 }),
    .b(2'b10),
    .fci(\u2_Display/lt159_c23 ),
    .fco(\u2_Display/lt159_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_26|u2_Display/lt159_25  (
    .a({\u2_Display/n6215 ,\u2_Display/n6216 }),
    .b(2'b10),
    .fci(\u2_Display/lt159_c25 ),
    .fco(\u2_Display/lt159_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_28|u2_Display/lt159_27  (
    .a({\u2_Display/n6213 ,\u2_Display/n6214 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c27 ),
    .fco(\u2_Display/lt159_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_2|u2_Display/lt159_1  (
    .a({\u2_Display/n6239 ,\u2_Display/n6240 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c1 ),
    .fco(\u2_Display/lt159_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_30|u2_Display/lt159_29  (
    .a({\u2_Display/n6211 ,\u2_Display/n6212 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c29 ),
    .fco(\u2_Display/lt159_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_4|u2_Display/lt159_3  (
    .a({\u2_Display/n6237 ,\u2_Display/n6238 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c3 ),
    .fco(\u2_Display/lt159_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_6|u2_Display/lt159_5  (
    .a({\u2_Display/n6235 ,\u2_Display/n6236 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c5 ),
    .fco(\u2_Display/lt159_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_8|u2_Display/lt159_7  (
    .a({\u2_Display/n6233 ,\u2_Display/n6234 }),
    .b(2'b00),
    .fci(\u2_Display/lt159_c7 ),
    .fco(\u2_Display/lt159_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt159_0|u2_Display/lt159_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt159_cout|u2_Display/lt159_31  (
    .a({1'b0,\u2_Display/n6210 }),
    .b(2'b10),
    .fci(\u2_Display/lt159_c31 ),
    .f({\u2_Display/n5084 ,open_n39503}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_0|u2_Display/lt160_cin  (
    .a({\u2_Display/n6276 ,1'b0}),
    .b({1'b0,open_n39509}),
    .fco(\u2_Display/lt160_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_10|u2_Display/lt160_9  (
    .a({\u2_Display/n6266 ,\u2_Display/n6267 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c9 ),
    .fco(\u2_Display/lt160_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_12|u2_Display/lt160_11  (
    .a({\u2_Display/n6264 ,\u2_Display/n6265 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c11 ),
    .fco(\u2_Display/lt160_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_14|u2_Display/lt160_13  (
    .a({\u2_Display/n6262 ,\u2_Display/n6263 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c13 ),
    .fco(\u2_Display/lt160_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_16|u2_Display/lt160_15  (
    .a({\u2_Display/n6260 ,\u2_Display/n6261 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c15 ),
    .fco(\u2_Display/lt160_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_18|u2_Display/lt160_17  (
    .a({\u2_Display/n6258 ,\u2_Display/n6259 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c17 ),
    .fco(\u2_Display/lt160_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_20|u2_Display/lt160_19  (
    .a({\u2_Display/n6256 ,\u2_Display/n6257 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c19 ),
    .fco(\u2_Display/lt160_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_22|u2_Display/lt160_21  (
    .a({\u2_Display/n6254 ,\u2_Display/n6255 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c21 ),
    .fco(\u2_Display/lt160_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_24|u2_Display/lt160_23  (
    .a({\u2_Display/n6252 ,\u2_Display/n6253 }),
    .b(2'b01),
    .fci(\u2_Display/lt160_c23 ),
    .fco(\u2_Display/lt160_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_26|u2_Display/lt160_25  (
    .a({\u2_Display/n6250 ,\u2_Display/n6251 }),
    .b(2'b01),
    .fci(\u2_Display/lt160_c25 ),
    .fco(\u2_Display/lt160_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_28|u2_Display/lt160_27  (
    .a({\u2_Display/n6248 ,\u2_Display/n6249 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c27 ),
    .fco(\u2_Display/lt160_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_2|u2_Display/lt160_1  (
    .a({\u2_Display/n6274 ,\u2_Display/n6275 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c1 ),
    .fco(\u2_Display/lt160_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_30|u2_Display/lt160_29  (
    .a({\u2_Display/n6246 ,\u2_Display/n6247 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c29 ),
    .fco(\u2_Display/lt160_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_4|u2_Display/lt160_3  (
    .a({\u2_Display/n6272 ,\u2_Display/n6273 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c3 ),
    .fco(\u2_Display/lt160_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_6|u2_Display/lt160_5  (
    .a({\u2_Display/n6270 ,\u2_Display/n6271 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c5 ),
    .fco(\u2_Display/lt160_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_8|u2_Display/lt160_7  (
    .a({\u2_Display/n6268 ,\u2_Display/n6269 }),
    .b(2'b00),
    .fci(\u2_Display/lt160_c7 ),
    .fco(\u2_Display/lt160_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt160_0|u2_Display/lt160_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt160_cout|u2_Display/lt160_31  (
    .a({1'b0,\u2_Display/n6245 }),
    .b(2'b10),
    .fci(\u2_Display/lt160_c31 ),
    .f({\u2_Display/n5119 ,open_n39913}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_0|u2_Display/lt161_cin  (
    .a({\u2_Display/n6311 ,1'b0}),
    .b({1'b0,open_n39919}),
    .fco(\u2_Display/lt161_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_10|u2_Display/lt161_9  (
    .a({\u2_Display/n6301 ,\u2_Display/n6302 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c9 ),
    .fco(\u2_Display/lt161_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_12|u2_Display/lt161_11  (
    .a({\u2_Display/n6299 ,\u2_Display/n6300 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c11 ),
    .fco(\u2_Display/lt161_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_14|u2_Display/lt161_13  (
    .a({\u2_Display/n6297 ,\u2_Display/n6298 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c13 ),
    .fco(\u2_Display/lt161_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_16|u2_Display/lt161_15  (
    .a({\u2_Display/n6295 ,\u2_Display/n6296 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c15 ),
    .fco(\u2_Display/lt161_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_18|u2_Display/lt161_17  (
    .a({\u2_Display/n6293 ,\u2_Display/n6294 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c17 ),
    .fco(\u2_Display/lt161_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_20|u2_Display/lt161_19  (
    .a({\u2_Display/n6291 ,\u2_Display/n6292 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c19 ),
    .fco(\u2_Display/lt161_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_22|u2_Display/lt161_21  (
    .a({\u2_Display/n6289 ,\u2_Display/n6290 }),
    .b(2'b10),
    .fci(\u2_Display/lt161_c21 ),
    .fco(\u2_Display/lt161_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_24|u2_Display/lt161_23  (
    .a({\u2_Display/n6287 ,\u2_Display/n6288 }),
    .b(2'b10),
    .fci(\u2_Display/lt161_c23 ),
    .fco(\u2_Display/lt161_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_26|u2_Display/lt161_25  (
    .a({\u2_Display/n6285 ,\u2_Display/n6286 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c25 ),
    .fco(\u2_Display/lt161_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_28|u2_Display/lt161_27  (
    .a({\u2_Display/n6283 ,\u2_Display/n6284 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c27 ),
    .fco(\u2_Display/lt161_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_2|u2_Display/lt161_1  (
    .a({\u2_Display/n6309 ,\u2_Display/n6310 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c1 ),
    .fco(\u2_Display/lt161_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_30|u2_Display/lt161_29  (
    .a({\u2_Display/n6281 ,\u2_Display/n6282 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c29 ),
    .fco(\u2_Display/lt161_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_4|u2_Display/lt161_3  (
    .a({\u2_Display/n6307 ,\u2_Display/n6308 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c3 ),
    .fco(\u2_Display/lt161_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_6|u2_Display/lt161_5  (
    .a({\u2_Display/n6305 ,\u2_Display/n6306 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c5 ),
    .fco(\u2_Display/lt161_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_8|u2_Display/lt161_7  (
    .a({\u2_Display/n6303 ,\u2_Display/n6304 }),
    .b(2'b00),
    .fci(\u2_Display/lt161_c7 ),
    .fco(\u2_Display/lt161_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt161_0|u2_Display/lt161_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt161_cout|u2_Display/lt161_31  (
    .a({1'b0,\u2_Display/n6280 }),
    .b(2'b10),
    .fci(\u2_Display/lt161_c31 ),
    .f({\u2_Display/n5154 ,open_n40323}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_0|u2_Display/lt162_cin  (
    .a({\u2_Display/n6346 ,1'b0}),
    .b({1'b0,open_n40329}),
    .fco(\u2_Display/lt162_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_10|u2_Display/lt162_9  (
    .a({\u2_Display/n6336 ,\u2_Display/n6337 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c9 ),
    .fco(\u2_Display/lt162_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_12|u2_Display/lt162_11  (
    .a({\u2_Display/n6334 ,\u2_Display/n6335 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c11 ),
    .fco(\u2_Display/lt162_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_14|u2_Display/lt162_13  (
    .a({\u2_Display/n6332 ,\u2_Display/n6333 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c13 ),
    .fco(\u2_Display/lt162_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_16|u2_Display/lt162_15  (
    .a({\u2_Display/n6330 ,\u2_Display/n6331 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c15 ),
    .fco(\u2_Display/lt162_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_18|u2_Display/lt162_17  (
    .a({\u2_Display/n6328 ,\u2_Display/n6329 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c17 ),
    .fco(\u2_Display/lt162_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_20|u2_Display/lt162_19  (
    .a({\u2_Display/n6326 ,\u2_Display/n6327 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c19 ),
    .fco(\u2_Display/lt162_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_22|u2_Display/lt162_21  (
    .a({\u2_Display/n6324 ,\u2_Display/n6325 }),
    .b(2'b01),
    .fci(\u2_Display/lt162_c21 ),
    .fco(\u2_Display/lt162_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_24|u2_Display/lt162_23  (
    .a({\u2_Display/n6322 ,\u2_Display/n6323 }),
    .b(2'b01),
    .fci(\u2_Display/lt162_c23 ),
    .fco(\u2_Display/lt162_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_26|u2_Display/lt162_25  (
    .a({\u2_Display/n6320 ,\u2_Display/n6321 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c25 ),
    .fco(\u2_Display/lt162_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_28|u2_Display/lt162_27  (
    .a({\u2_Display/n6318 ,\u2_Display/n6319 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c27 ),
    .fco(\u2_Display/lt162_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_2|u2_Display/lt162_1  (
    .a({\u2_Display/n6344 ,\u2_Display/n6345 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c1 ),
    .fco(\u2_Display/lt162_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_30|u2_Display/lt162_29  (
    .a({\u2_Display/n6316 ,\u2_Display/n6317 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c29 ),
    .fco(\u2_Display/lt162_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_4|u2_Display/lt162_3  (
    .a({\u2_Display/n6342 ,\u2_Display/n6343 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c3 ),
    .fco(\u2_Display/lt162_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_6|u2_Display/lt162_5  (
    .a({\u2_Display/n6340 ,\u2_Display/n6341 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c5 ),
    .fco(\u2_Display/lt162_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_8|u2_Display/lt162_7  (
    .a({\u2_Display/n6338 ,\u2_Display/n6339 }),
    .b(2'b00),
    .fci(\u2_Display/lt162_c7 ),
    .fco(\u2_Display/lt162_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt162_0|u2_Display/lt162_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt162_cout|u2_Display/lt162_31  (
    .a({1'b0,\u2_Display/n6315 }),
    .b(2'b10),
    .fci(\u2_Display/lt162_c31 ),
    .f({\u2_Display/n5189 ,open_n40733}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_0|u2_Display/lt163_cin  (
    .a({\u2_Display/n5223 ,1'b0}),
    .b({1'b0,open_n40739}),
    .fco(\u2_Display/lt163_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_10|u2_Display/lt163_9  (
    .a({\u2_Display/n5213 ,\u2_Display/n5214 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c9 ),
    .fco(\u2_Display/lt163_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_12|u2_Display/lt163_11  (
    .a({\u2_Display/n5211 ,\u2_Display/n5212 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c11 ),
    .fco(\u2_Display/lt163_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_14|u2_Display/lt163_13  (
    .a({\u2_Display/n5209 ,\u2_Display/n5210 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c13 ),
    .fco(\u2_Display/lt163_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_16|u2_Display/lt163_15  (
    .a({\u2_Display/n5207 ,\u2_Display/n5208 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c15 ),
    .fco(\u2_Display/lt163_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_18|u2_Display/lt163_17  (
    .a({\u2_Display/n5205 ,\u2_Display/n5206 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c17 ),
    .fco(\u2_Display/lt163_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_20|u2_Display/lt163_19  (
    .a({\u2_Display/n5203 ,\u2_Display/n5204 }),
    .b(2'b10),
    .fci(\u2_Display/lt163_c19 ),
    .fco(\u2_Display/lt163_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_22|u2_Display/lt163_21  (
    .a({\u2_Display/n5201 ,\u2_Display/n5202 }),
    .b(2'b10),
    .fci(\u2_Display/lt163_c21 ),
    .fco(\u2_Display/lt163_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_24|u2_Display/lt163_23  (
    .a({\u2_Display/n5199 ,\u2_Display/n5200 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c23 ),
    .fco(\u2_Display/lt163_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_26|u2_Display/lt163_25  (
    .a({\u2_Display/n5197 ,\u2_Display/n5198 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c25 ),
    .fco(\u2_Display/lt163_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_28|u2_Display/lt163_27  (
    .a({\u2_Display/n6353 ,\u2_Display/n5196 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c27 ),
    .fco(\u2_Display/lt163_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_2|u2_Display/lt163_1  (
    .a({\u2_Display/n5221 ,\u2_Display/n5222 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c1 ),
    .fco(\u2_Display/lt163_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_30|u2_Display/lt163_29  (
    .a({\u2_Display/n6351 ,\u2_Display/n6352 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c29 ),
    .fco(\u2_Display/lt163_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_4|u2_Display/lt163_3  (
    .a({\u2_Display/n5219 ,\u2_Display/n5220 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c3 ),
    .fco(\u2_Display/lt163_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_6|u2_Display/lt163_5  (
    .a({\u2_Display/n5217 ,\u2_Display/n5218 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c5 ),
    .fco(\u2_Display/lt163_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_8|u2_Display/lt163_7  (
    .a({\u2_Display/n5215 ,\u2_Display/n5216 }),
    .b(2'b00),
    .fci(\u2_Display/lt163_c7 ),
    .fco(\u2_Display/lt163_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt163_0|u2_Display/lt163_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt163_cout|u2_Display/lt163_31  (
    .a({1'b0,\u2_Display/n6350 }),
    .b(2'b10),
    .fci(\u2_Display/lt163_c31 ),
    .f({\u2_Display/n5224 ,open_n41143}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_0|u2_Display/lt164_cin  (
    .a({\u2_Display/n5258 ,1'b0}),
    .b({1'b0,open_n41149}),
    .fco(\u2_Display/lt164_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_10|u2_Display/lt164_9  (
    .a({\u2_Display/n5248 ,\u2_Display/n5249 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c9 ),
    .fco(\u2_Display/lt164_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_12|u2_Display/lt164_11  (
    .a({\u2_Display/n5246 ,\u2_Display/n5247 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c11 ),
    .fco(\u2_Display/lt164_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_14|u2_Display/lt164_13  (
    .a({\u2_Display/n5244 ,\u2_Display/n5245 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c13 ),
    .fco(\u2_Display/lt164_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_16|u2_Display/lt164_15  (
    .a({\u2_Display/n5242 ,\u2_Display/n5243 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c15 ),
    .fco(\u2_Display/lt164_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_18|u2_Display/lt164_17  (
    .a({\u2_Display/n5240 ,\u2_Display/n5241 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c17 ),
    .fco(\u2_Display/lt164_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_20|u2_Display/lt164_19  (
    .a({\u2_Display/n5238 ,\u2_Display/n5239 }),
    .b(2'b01),
    .fci(\u2_Display/lt164_c19 ),
    .fco(\u2_Display/lt164_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_22|u2_Display/lt164_21  (
    .a({\u2_Display/n5236 ,\u2_Display/n5237 }),
    .b(2'b01),
    .fci(\u2_Display/lt164_c21 ),
    .fco(\u2_Display/lt164_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_24|u2_Display/lt164_23  (
    .a({\u2_Display/n5234 ,\u2_Display/n5235 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c23 ),
    .fco(\u2_Display/lt164_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_26|u2_Display/lt164_25  (
    .a({\u2_Display/n5232 ,\u2_Display/n5233 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c25 ),
    .fco(\u2_Display/lt164_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_28|u2_Display/lt164_27  (
    .a({\u2_Display/n5230 ,\u2_Display/n5231 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c27 ),
    .fco(\u2_Display/lt164_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_2|u2_Display/lt164_1  (
    .a({\u2_Display/n5256 ,\u2_Display/n5257 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c1 ),
    .fco(\u2_Display/lt164_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_30|u2_Display/lt164_29  (
    .a({\u2_Display/n5228 ,\u2_Display/n5229 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c29 ),
    .fco(\u2_Display/lt164_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_4|u2_Display/lt164_3  (
    .a({\u2_Display/n5254 ,\u2_Display/n5255 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c3 ),
    .fco(\u2_Display/lt164_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_6|u2_Display/lt164_5  (
    .a({\u2_Display/n5252 ,\u2_Display/n5253 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c5 ),
    .fco(\u2_Display/lt164_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_8|u2_Display/lt164_7  (
    .a({\u2_Display/n5250 ,\u2_Display/n5251 }),
    .b(2'b00),
    .fci(\u2_Display/lt164_c7 ),
    .fco(\u2_Display/lt164_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt164_0|u2_Display/lt164_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt164_cout|u2_Display/lt164_31  (
    .a({1'b0,\u2_Display/n5227 }),
    .b(2'b10),
    .fci(\u2_Display/lt164_c31 ),
    .f({\u2_Display/n5259 ,open_n41553}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_0|u2_Display/lt165_cin  (
    .a({\u2_Display/n5293 ,1'b0}),
    .b({1'b0,open_n41559}),
    .fco(\u2_Display/lt165_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_10|u2_Display/lt165_9  (
    .a({\u2_Display/n5283 ,\u2_Display/n5284 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c9 ),
    .fco(\u2_Display/lt165_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_12|u2_Display/lt165_11  (
    .a({\u2_Display/n5281 ,\u2_Display/n5282 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c11 ),
    .fco(\u2_Display/lt165_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_14|u2_Display/lt165_13  (
    .a({\u2_Display/n5279 ,\u2_Display/n5280 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c13 ),
    .fco(\u2_Display/lt165_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_16|u2_Display/lt165_15  (
    .a({\u2_Display/n5277 ,\u2_Display/n5278 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c15 ),
    .fco(\u2_Display/lt165_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_18|u2_Display/lt165_17  (
    .a({\u2_Display/n5275 ,\u2_Display/n5276 }),
    .b(2'b10),
    .fci(\u2_Display/lt165_c17 ),
    .fco(\u2_Display/lt165_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_20|u2_Display/lt165_19  (
    .a({\u2_Display/n5273 ,\u2_Display/n5274 }),
    .b(2'b10),
    .fci(\u2_Display/lt165_c19 ),
    .fco(\u2_Display/lt165_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_22|u2_Display/lt165_21  (
    .a({\u2_Display/n5271 ,\u2_Display/n5272 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c21 ),
    .fco(\u2_Display/lt165_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_24|u2_Display/lt165_23  (
    .a({\u2_Display/n5269 ,\u2_Display/n5270 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c23 ),
    .fco(\u2_Display/lt165_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_26|u2_Display/lt165_25  (
    .a({\u2_Display/n5267 ,\u2_Display/n5268 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c25 ),
    .fco(\u2_Display/lt165_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_28|u2_Display/lt165_27  (
    .a({\u2_Display/n5265 ,\u2_Display/n5266 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c27 ),
    .fco(\u2_Display/lt165_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_2|u2_Display/lt165_1  (
    .a({\u2_Display/n5291 ,\u2_Display/n5292 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c1 ),
    .fco(\u2_Display/lt165_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_30|u2_Display/lt165_29  (
    .a({\u2_Display/n5263 ,\u2_Display/n5264 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c29 ),
    .fco(\u2_Display/lt165_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_4|u2_Display/lt165_3  (
    .a({\u2_Display/n5289 ,\u2_Display/n5290 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c3 ),
    .fco(\u2_Display/lt165_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_6|u2_Display/lt165_5  (
    .a({\u2_Display/n5287 ,\u2_Display/n5288 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c5 ),
    .fco(\u2_Display/lt165_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_8|u2_Display/lt165_7  (
    .a({\u2_Display/n5285 ,\u2_Display/n5286 }),
    .b(2'b00),
    .fci(\u2_Display/lt165_c7 ),
    .fco(\u2_Display/lt165_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt165_0|u2_Display/lt165_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt165_cout|u2_Display/lt165_31  (
    .a({1'b0,\u2_Display/n5262 }),
    .b(2'b10),
    .fci(\u2_Display/lt165_c31 ),
    .f({\u2_Display/n5294 ,open_n41963}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_0|u2_Display/lt166_cin  (
    .a({\u2_Display/n5328 ,1'b0}),
    .b({1'b0,open_n41969}),
    .fco(\u2_Display/lt166_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_10|u2_Display/lt166_9  (
    .a({\u2_Display/n5318 ,\u2_Display/n5319 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c9 ),
    .fco(\u2_Display/lt166_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_12|u2_Display/lt166_11  (
    .a({\u2_Display/n5316 ,\u2_Display/n5317 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c11 ),
    .fco(\u2_Display/lt166_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_14|u2_Display/lt166_13  (
    .a({\u2_Display/n5314 ,\u2_Display/n5315 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c13 ),
    .fco(\u2_Display/lt166_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_16|u2_Display/lt166_15  (
    .a({\u2_Display/n5312 ,\u2_Display/n5313 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c15 ),
    .fco(\u2_Display/lt166_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_18|u2_Display/lt166_17  (
    .a({\u2_Display/n5310 ,\u2_Display/n5311 }),
    .b(2'b01),
    .fci(\u2_Display/lt166_c17 ),
    .fco(\u2_Display/lt166_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_20|u2_Display/lt166_19  (
    .a({\u2_Display/n5308 ,\u2_Display/n5309 }),
    .b(2'b01),
    .fci(\u2_Display/lt166_c19 ),
    .fco(\u2_Display/lt166_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_22|u2_Display/lt166_21  (
    .a({\u2_Display/n5306 ,\u2_Display/n5307 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c21 ),
    .fco(\u2_Display/lt166_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_24|u2_Display/lt166_23  (
    .a({\u2_Display/n5304 ,\u2_Display/n5305 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c23 ),
    .fco(\u2_Display/lt166_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_26|u2_Display/lt166_25  (
    .a({\u2_Display/n5302 ,\u2_Display/n5303 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c25 ),
    .fco(\u2_Display/lt166_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_28|u2_Display/lt166_27  (
    .a({\u2_Display/n5300 ,\u2_Display/n5301 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c27 ),
    .fco(\u2_Display/lt166_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_2|u2_Display/lt166_1  (
    .a({\u2_Display/n5326 ,\u2_Display/n5327 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c1 ),
    .fco(\u2_Display/lt166_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_30|u2_Display/lt166_29  (
    .a({\u2_Display/n5298 ,\u2_Display/n5299 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c29 ),
    .fco(\u2_Display/lt166_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_4|u2_Display/lt166_3  (
    .a({\u2_Display/n5324 ,\u2_Display/n5325 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c3 ),
    .fco(\u2_Display/lt166_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_6|u2_Display/lt166_5  (
    .a({\u2_Display/n5322 ,\u2_Display/n5323 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c5 ),
    .fco(\u2_Display/lt166_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_8|u2_Display/lt166_7  (
    .a({\u2_Display/n5320 ,\u2_Display/n5321 }),
    .b(2'b00),
    .fci(\u2_Display/lt166_c7 ),
    .fco(\u2_Display/lt166_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt166_0|u2_Display/lt166_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt166_cout|u2_Display/lt166_31  (
    .a({1'b0,\u2_Display/n5297 }),
    .b(2'b10),
    .fci(\u2_Display/lt166_c31 ),
    .f({\u2_Display/n5329 ,open_n42373}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_0|u2_Display/lt167_cin  (
    .a({\u2_Display/n5363 ,1'b0}),
    .b({1'b0,open_n42379}),
    .fco(\u2_Display/lt167_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_10|u2_Display/lt167_9  (
    .a({\u2_Display/n5353 ,\u2_Display/n5354 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c9 ),
    .fco(\u2_Display/lt167_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_12|u2_Display/lt167_11  (
    .a({\u2_Display/n5351 ,\u2_Display/n5352 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c11 ),
    .fco(\u2_Display/lt167_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_14|u2_Display/lt167_13  (
    .a({\u2_Display/n5349 ,\u2_Display/n5350 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c13 ),
    .fco(\u2_Display/lt167_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_16|u2_Display/lt167_15  (
    .a({\u2_Display/n5347 ,\u2_Display/n5348 }),
    .b(2'b10),
    .fci(\u2_Display/lt167_c15 ),
    .fco(\u2_Display/lt167_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_18|u2_Display/lt167_17  (
    .a({\u2_Display/n5345 ,\u2_Display/n5346 }),
    .b(2'b10),
    .fci(\u2_Display/lt167_c17 ),
    .fco(\u2_Display/lt167_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_20|u2_Display/lt167_19  (
    .a({\u2_Display/n5343 ,\u2_Display/n5344 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c19 ),
    .fco(\u2_Display/lt167_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_22|u2_Display/lt167_21  (
    .a({\u2_Display/n5341 ,\u2_Display/n5342 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c21 ),
    .fco(\u2_Display/lt167_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_24|u2_Display/lt167_23  (
    .a({\u2_Display/n5339 ,\u2_Display/n5340 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c23 ),
    .fco(\u2_Display/lt167_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_26|u2_Display/lt167_25  (
    .a({\u2_Display/n5337 ,\u2_Display/n5338 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c25 ),
    .fco(\u2_Display/lt167_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_28|u2_Display/lt167_27  (
    .a({\u2_Display/n5335 ,\u2_Display/n5336 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c27 ),
    .fco(\u2_Display/lt167_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_2|u2_Display/lt167_1  (
    .a({\u2_Display/n5361 ,\u2_Display/n5362 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c1 ),
    .fco(\u2_Display/lt167_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_30|u2_Display/lt167_29  (
    .a({\u2_Display/n5333 ,\u2_Display/n5334 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c29 ),
    .fco(\u2_Display/lt167_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_4|u2_Display/lt167_3  (
    .a({\u2_Display/n5359 ,\u2_Display/n5360 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c3 ),
    .fco(\u2_Display/lt167_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_6|u2_Display/lt167_5  (
    .a({\u2_Display/n5357 ,\u2_Display/n5358 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c5 ),
    .fco(\u2_Display/lt167_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_8|u2_Display/lt167_7  (
    .a({\u2_Display/n5355 ,\u2_Display/n5356 }),
    .b(2'b00),
    .fci(\u2_Display/lt167_c7 ),
    .fco(\u2_Display/lt167_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt167_0|u2_Display/lt167_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt167_cout|u2_Display/lt167_31  (
    .a({1'b0,\u2_Display/n5332 }),
    .b(2'b10),
    .fci(\u2_Display/lt167_c31 ),
    .f({\u2_Display/n5364 ,open_n42783}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_0|u2_Display/lt168_cin  (
    .a({\u2_Display/n5398 ,1'b0}),
    .b({1'b0,open_n42789}),
    .fco(\u2_Display/lt168_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_10|u2_Display/lt168_9  (
    .a({\u2_Display/n5388 ,\u2_Display/n5389 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c9 ),
    .fco(\u2_Display/lt168_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_12|u2_Display/lt168_11  (
    .a({\u2_Display/n5386 ,\u2_Display/n5387 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c11 ),
    .fco(\u2_Display/lt168_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_14|u2_Display/lt168_13  (
    .a({\u2_Display/n5384 ,\u2_Display/n5385 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c13 ),
    .fco(\u2_Display/lt168_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_16|u2_Display/lt168_15  (
    .a({\u2_Display/n5382 ,\u2_Display/n5383 }),
    .b(2'b01),
    .fci(\u2_Display/lt168_c15 ),
    .fco(\u2_Display/lt168_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_18|u2_Display/lt168_17  (
    .a({\u2_Display/n5380 ,\u2_Display/n5381 }),
    .b(2'b01),
    .fci(\u2_Display/lt168_c17 ),
    .fco(\u2_Display/lt168_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_20|u2_Display/lt168_19  (
    .a({\u2_Display/n5378 ,\u2_Display/n5379 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c19 ),
    .fco(\u2_Display/lt168_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_22|u2_Display/lt168_21  (
    .a({\u2_Display/n5376 ,\u2_Display/n5377 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c21 ),
    .fco(\u2_Display/lt168_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_24|u2_Display/lt168_23  (
    .a({\u2_Display/n5374 ,\u2_Display/n5375 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c23 ),
    .fco(\u2_Display/lt168_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_26|u2_Display/lt168_25  (
    .a({\u2_Display/n5372 ,\u2_Display/n5373 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c25 ),
    .fco(\u2_Display/lt168_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_28|u2_Display/lt168_27  (
    .a({\u2_Display/n5370 ,\u2_Display/n5371 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c27 ),
    .fco(\u2_Display/lt168_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_2|u2_Display/lt168_1  (
    .a({\u2_Display/n5396 ,\u2_Display/n5397 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c1 ),
    .fco(\u2_Display/lt168_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_30|u2_Display/lt168_29  (
    .a({\u2_Display/n5368 ,\u2_Display/n5369 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c29 ),
    .fco(\u2_Display/lt168_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_4|u2_Display/lt168_3  (
    .a({\u2_Display/n5394 ,\u2_Display/n5395 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c3 ),
    .fco(\u2_Display/lt168_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_6|u2_Display/lt168_5  (
    .a({\u2_Display/n5392 ,\u2_Display/n5393 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c5 ),
    .fco(\u2_Display/lt168_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_8|u2_Display/lt168_7  (
    .a({\u2_Display/n5390 ,\u2_Display/n5391 }),
    .b(2'b00),
    .fci(\u2_Display/lt168_c7 ),
    .fco(\u2_Display/lt168_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt168_0|u2_Display/lt168_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt168_cout|u2_Display/lt168_31  (
    .a({1'b0,\u2_Display/n5367 }),
    .b(2'b10),
    .fci(\u2_Display/lt168_c31 ),
    .f({\u2_Display/n5399 ,open_n43193}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_0|u2_Display/lt169_cin  (
    .a({\u2_Display/n5433 ,1'b0}),
    .b({1'b0,open_n43199}),
    .fco(\u2_Display/lt169_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_10|u2_Display/lt169_9  (
    .a({\u2_Display/n5423 ,\u2_Display/n5424 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c9 ),
    .fco(\u2_Display/lt169_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_12|u2_Display/lt169_11  (
    .a({\u2_Display/n5421 ,\u2_Display/n5422 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c11 ),
    .fco(\u2_Display/lt169_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_14|u2_Display/lt169_13  (
    .a({\u2_Display/n5419 ,\u2_Display/n5420 }),
    .b(2'b10),
    .fci(\u2_Display/lt169_c13 ),
    .fco(\u2_Display/lt169_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_16|u2_Display/lt169_15  (
    .a({\u2_Display/n5417 ,\u2_Display/n5418 }),
    .b(2'b10),
    .fci(\u2_Display/lt169_c15 ),
    .fco(\u2_Display/lt169_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_18|u2_Display/lt169_17  (
    .a({\u2_Display/n5415 ,\u2_Display/n5416 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c17 ),
    .fco(\u2_Display/lt169_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_20|u2_Display/lt169_19  (
    .a({\u2_Display/n5413 ,\u2_Display/n5414 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c19 ),
    .fco(\u2_Display/lt169_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_22|u2_Display/lt169_21  (
    .a({\u2_Display/n5411 ,\u2_Display/n5412 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c21 ),
    .fco(\u2_Display/lt169_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_24|u2_Display/lt169_23  (
    .a({\u2_Display/n5409 ,\u2_Display/n5410 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c23 ),
    .fco(\u2_Display/lt169_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_26|u2_Display/lt169_25  (
    .a({\u2_Display/n5407 ,\u2_Display/n5408 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c25 ),
    .fco(\u2_Display/lt169_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_28|u2_Display/lt169_27  (
    .a({\u2_Display/n5405 ,\u2_Display/n5406 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c27 ),
    .fco(\u2_Display/lt169_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_2|u2_Display/lt169_1  (
    .a({\u2_Display/n5431 ,\u2_Display/n5432 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c1 ),
    .fco(\u2_Display/lt169_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_30|u2_Display/lt169_29  (
    .a({\u2_Display/n5403 ,\u2_Display/n5404 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c29 ),
    .fco(\u2_Display/lt169_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_4|u2_Display/lt169_3  (
    .a({\u2_Display/n5429 ,\u2_Display/n5430 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c3 ),
    .fco(\u2_Display/lt169_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_6|u2_Display/lt169_5  (
    .a({\u2_Display/n5427 ,\u2_Display/n5428 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c5 ),
    .fco(\u2_Display/lt169_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_8|u2_Display/lt169_7  (
    .a({\u2_Display/n5425 ,\u2_Display/n5426 }),
    .b(2'b00),
    .fci(\u2_Display/lt169_c7 ),
    .fco(\u2_Display/lt169_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt169_0|u2_Display/lt169_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt169_cout|u2_Display/lt169_31  (
    .a({1'b0,\u2_Display/n5402 }),
    .b(2'b10),
    .fci(\u2_Display/lt169_c31 ),
    .f({\u2_Display/n5434 ,open_n43603}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_0|u2_Display/lt170_cin  (
    .a({\u2_Display/n5468 ,1'b0}),
    .b({1'b0,open_n43609}),
    .fco(\u2_Display/lt170_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_10|u2_Display/lt170_9  (
    .a({\u2_Display/n5458 ,\u2_Display/n5459 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c9 ),
    .fco(\u2_Display/lt170_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_12|u2_Display/lt170_11  (
    .a({\u2_Display/n5456 ,\u2_Display/n5457 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c11 ),
    .fco(\u2_Display/lt170_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_14|u2_Display/lt170_13  (
    .a({\u2_Display/n5454 ,\u2_Display/n5455 }),
    .b(2'b01),
    .fci(\u2_Display/lt170_c13 ),
    .fco(\u2_Display/lt170_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_16|u2_Display/lt170_15  (
    .a({\u2_Display/n5452 ,\u2_Display/n5453 }),
    .b(2'b01),
    .fci(\u2_Display/lt170_c15 ),
    .fco(\u2_Display/lt170_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_18|u2_Display/lt170_17  (
    .a({\u2_Display/n5450 ,\u2_Display/n5451 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c17 ),
    .fco(\u2_Display/lt170_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_20|u2_Display/lt170_19  (
    .a({\u2_Display/n5448 ,\u2_Display/n5449 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c19 ),
    .fco(\u2_Display/lt170_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_22|u2_Display/lt170_21  (
    .a({\u2_Display/n5446 ,\u2_Display/n5447 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c21 ),
    .fco(\u2_Display/lt170_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_24|u2_Display/lt170_23  (
    .a({\u2_Display/n5444 ,\u2_Display/n5445 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c23 ),
    .fco(\u2_Display/lt170_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_26|u2_Display/lt170_25  (
    .a({\u2_Display/n5442 ,\u2_Display/n5443 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c25 ),
    .fco(\u2_Display/lt170_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_28|u2_Display/lt170_27  (
    .a({\u2_Display/n5440 ,\u2_Display/n5441 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c27 ),
    .fco(\u2_Display/lt170_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_2|u2_Display/lt170_1  (
    .a({\u2_Display/n5466 ,\u2_Display/n5467 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c1 ),
    .fco(\u2_Display/lt170_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_30|u2_Display/lt170_29  (
    .a({\u2_Display/n5438 ,\u2_Display/n5439 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c29 ),
    .fco(\u2_Display/lt170_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_4|u2_Display/lt170_3  (
    .a({\u2_Display/n5464 ,\u2_Display/n5465 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c3 ),
    .fco(\u2_Display/lt170_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_6|u2_Display/lt170_5  (
    .a({\u2_Display/n5462 ,\u2_Display/n5463 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c5 ),
    .fco(\u2_Display/lt170_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_8|u2_Display/lt170_7  (
    .a({\u2_Display/n5460 ,\u2_Display/n5461 }),
    .b(2'b00),
    .fci(\u2_Display/lt170_c7 ),
    .fco(\u2_Display/lt170_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt170_0|u2_Display/lt170_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt170_cout|u2_Display/lt170_31  (
    .a({1'b0,\u2_Display/n5437 }),
    .b(2'b10),
    .fci(\u2_Display/lt170_c31 ),
    .f({\u2_Display/n5469 ,open_n44013}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_0|u2_Display/lt171_cin  (
    .a({\u2_Display/n5503 ,1'b0}),
    .b({1'b0,open_n44019}),
    .fco(\u2_Display/lt171_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_10|u2_Display/lt171_9  (
    .a({\u2_Display/n5493 ,\u2_Display/n5494 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c9 ),
    .fco(\u2_Display/lt171_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_12|u2_Display/lt171_11  (
    .a({\u2_Display/n5491 ,\u2_Display/n5492 }),
    .b(2'b10),
    .fci(\u2_Display/lt171_c11 ),
    .fco(\u2_Display/lt171_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_14|u2_Display/lt171_13  (
    .a({\u2_Display/n5489 ,\u2_Display/n5490 }),
    .b(2'b10),
    .fci(\u2_Display/lt171_c13 ),
    .fco(\u2_Display/lt171_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_16|u2_Display/lt171_15  (
    .a({\u2_Display/n5487 ,\u2_Display/n5488 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c15 ),
    .fco(\u2_Display/lt171_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_18|u2_Display/lt171_17  (
    .a({\u2_Display/n5485 ,\u2_Display/n5486 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c17 ),
    .fco(\u2_Display/lt171_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_20|u2_Display/lt171_19  (
    .a({\u2_Display/n5483 ,\u2_Display/n5484 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c19 ),
    .fco(\u2_Display/lt171_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_22|u2_Display/lt171_21  (
    .a({\u2_Display/n5481 ,\u2_Display/n5482 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c21 ),
    .fco(\u2_Display/lt171_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_24|u2_Display/lt171_23  (
    .a({\u2_Display/n5479 ,\u2_Display/n5480 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c23 ),
    .fco(\u2_Display/lt171_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_26|u2_Display/lt171_25  (
    .a({\u2_Display/n5477 ,\u2_Display/n5478 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c25 ),
    .fco(\u2_Display/lt171_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_28|u2_Display/lt171_27  (
    .a({\u2_Display/n5475 ,\u2_Display/n5476 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c27 ),
    .fco(\u2_Display/lt171_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_2|u2_Display/lt171_1  (
    .a({\u2_Display/n5501 ,\u2_Display/n5502 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c1 ),
    .fco(\u2_Display/lt171_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_30|u2_Display/lt171_29  (
    .a({\u2_Display/n5473 ,\u2_Display/n5474 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c29 ),
    .fco(\u2_Display/lt171_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_4|u2_Display/lt171_3  (
    .a({\u2_Display/n5499 ,\u2_Display/n5500 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c3 ),
    .fco(\u2_Display/lt171_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_6|u2_Display/lt171_5  (
    .a({\u2_Display/n5497 ,\u2_Display/n5498 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c5 ),
    .fco(\u2_Display/lt171_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_8|u2_Display/lt171_7  (
    .a({\u2_Display/n5495 ,\u2_Display/n5496 }),
    .b(2'b00),
    .fci(\u2_Display/lt171_c7 ),
    .fco(\u2_Display/lt171_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt171_0|u2_Display/lt171_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt171_cout|u2_Display/lt171_31  (
    .a({1'b0,\u2_Display/n5472 }),
    .b(2'b10),
    .fci(\u2_Display/lt171_c31 ),
    .f({\u2_Display/n5504 ,open_n44423}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_0|u2_Display/lt172_cin  (
    .a({\u2_Display/n5538 ,1'b0}),
    .b({1'b0,open_n44429}),
    .fco(\u2_Display/lt172_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_10|u2_Display/lt172_9  (
    .a({\u2_Display/n5528 ,\u2_Display/n5529 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c9 ),
    .fco(\u2_Display/lt172_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_12|u2_Display/lt172_11  (
    .a({\u2_Display/n5526 ,\u2_Display/n5527 }),
    .b(2'b01),
    .fci(\u2_Display/lt172_c11 ),
    .fco(\u2_Display/lt172_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_14|u2_Display/lt172_13  (
    .a({\u2_Display/n5524 ,\u2_Display/n5525 }),
    .b(2'b01),
    .fci(\u2_Display/lt172_c13 ),
    .fco(\u2_Display/lt172_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_16|u2_Display/lt172_15  (
    .a({\u2_Display/n5522 ,\u2_Display/n5523 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c15 ),
    .fco(\u2_Display/lt172_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_18|u2_Display/lt172_17  (
    .a({\u2_Display/n5520 ,\u2_Display/n5521 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c17 ),
    .fco(\u2_Display/lt172_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_20|u2_Display/lt172_19  (
    .a({\u2_Display/n5518 ,\u2_Display/n5519 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c19 ),
    .fco(\u2_Display/lt172_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_22|u2_Display/lt172_21  (
    .a({\u2_Display/n5516 ,\u2_Display/n5517 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c21 ),
    .fco(\u2_Display/lt172_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_24|u2_Display/lt172_23  (
    .a({\u2_Display/n5514 ,\u2_Display/n5515 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c23 ),
    .fco(\u2_Display/lt172_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_26|u2_Display/lt172_25  (
    .a({\u2_Display/n5512 ,\u2_Display/n5513 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c25 ),
    .fco(\u2_Display/lt172_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_28|u2_Display/lt172_27  (
    .a({\u2_Display/n5510 ,\u2_Display/n5511 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c27 ),
    .fco(\u2_Display/lt172_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_2|u2_Display/lt172_1  (
    .a({\u2_Display/n5536 ,\u2_Display/n5537 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c1 ),
    .fco(\u2_Display/lt172_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_30|u2_Display/lt172_29  (
    .a({\u2_Display/n5508 ,\u2_Display/n5509 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c29 ),
    .fco(\u2_Display/lt172_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_4|u2_Display/lt172_3  (
    .a({\u2_Display/n5534 ,\u2_Display/n5535 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c3 ),
    .fco(\u2_Display/lt172_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_6|u2_Display/lt172_5  (
    .a({\u2_Display/n5532 ,\u2_Display/n5533 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c5 ),
    .fco(\u2_Display/lt172_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_8|u2_Display/lt172_7  (
    .a({\u2_Display/n5530 ,\u2_Display/n5531 }),
    .b(2'b00),
    .fci(\u2_Display/lt172_c7 ),
    .fco(\u2_Display/lt172_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt172_0|u2_Display/lt172_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt172_cout|u2_Display/lt172_31  (
    .a({1'b0,\u2_Display/n5507 }),
    .b(2'b10),
    .fci(\u2_Display/lt172_c31 ),
    .f({\u2_Display/n5539 ,open_n44833}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_0|u2_Display/lt173_cin  (
    .a({\u2_Display/n5573 ,1'b0}),
    .b({1'b0,open_n44839}),
    .fco(\u2_Display/lt173_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_10|u2_Display/lt173_9  (
    .a({\u2_Display/n5563 ,\u2_Display/n5564 }),
    .b(2'b10),
    .fci(\u2_Display/lt173_c9 ),
    .fco(\u2_Display/lt173_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_12|u2_Display/lt173_11  (
    .a({\u2_Display/n5561 ,\u2_Display/n5562 }),
    .b(2'b10),
    .fci(\u2_Display/lt173_c11 ),
    .fco(\u2_Display/lt173_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_14|u2_Display/lt173_13  (
    .a({\u2_Display/n5559 ,\u2_Display/n5560 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c13 ),
    .fco(\u2_Display/lt173_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_16|u2_Display/lt173_15  (
    .a({\u2_Display/n5557 ,\u2_Display/n5558 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c15 ),
    .fco(\u2_Display/lt173_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_18|u2_Display/lt173_17  (
    .a({\u2_Display/n5555 ,\u2_Display/n5556 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c17 ),
    .fco(\u2_Display/lt173_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_20|u2_Display/lt173_19  (
    .a({\u2_Display/n5553 ,\u2_Display/n5554 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c19 ),
    .fco(\u2_Display/lt173_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_22|u2_Display/lt173_21  (
    .a({\u2_Display/n5551 ,\u2_Display/n5552 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c21 ),
    .fco(\u2_Display/lt173_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_24|u2_Display/lt173_23  (
    .a({\u2_Display/n5549 ,\u2_Display/n5550 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c23 ),
    .fco(\u2_Display/lt173_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_26|u2_Display/lt173_25  (
    .a({\u2_Display/n5547 ,\u2_Display/n5548 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c25 ),
    .fco(\u2_Display/lt173_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_28|u2_Display/lt173_27  (
    .a({\u2_Display/n5545 ,\u2_Display/n5546 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c27 ),
    .fco(\u2_Display/lt173_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_2|u2_Display/lt173_1  (
    .a({\u2_Display/n5571 ,\u2_Display/n5572 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c1 ),
    .fco(\u2_Display/lt173_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_30|u2_Display/lt173_29  (
    .a({\u2_Display/n5543 ,\u2_Display/n5544 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c29 ),
    .fco(\u2_Display/lt173_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_4|u2_Display/lt173_3  (
    .a({\u2_Display/n5569 ,\u2_Display/n5570 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c3 ),
    .fco(\u2_Display/lt173_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_6|u2_Display/lt173_5  (
    .a({\u2_Display/n5567 ,\u2_Display/n5568 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c5 ),
    .fco(\u2_Display/lt173_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_8|u2_Display/lt173_7  (
    .a({\u2_Display/n5565 ,\u2_Display/n5566 }),
    .b(2'b00),
    .fci(\u2_Display/lt173_c7 ),
    .fco(\u2_Display/lt173_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt173_0|u2_Display/lt173_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt173_cout|u2_Display/lt173_31  (
    .a({1'b0,\u2_Display/n5542 }),
    .b(2'b10),
    .fci(\u2_Display/lt173_c31 ),
    .f({\u2_Display/n5574 ,open_n45243}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_0|u2_Display/lt174_cin  (
    .a({\u2_Display/n5608 ,1'b0}),
    .b({1'b0,open_n45249}),
    .fco(\u2_Display/lt174_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_10|u2_Display/lt174_9  (
    .a({\u2_Display/n5598 ,\u2_Display/n5599 }),
    .b(2'b01),
    .fci(\u2_Display/lt174_c9 ),
    .fco(\u2_Display/lt174_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_12|u2_Display/lt174_11  (
    .a({\u2_Display/n5596 ,\u2_Display/n5597 }),
    .b(2'b01),
    .fci(\u2_Display/lt174_c11 ),
    .fco(\u2_Display/lt174_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_14|u2_Display/lt174_13  (
    .a({\u2_Display/n5594 ,\u2_Display/n5595 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c13 ),
    .fco(\u2_Display/lt174_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_16|u2_Display/lt174_15  (
    .a({\u2_Display/n5592 ,\u2_Display/n5593 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c15 ),
    .fco(\u2_Display/lt174_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_18|u2_Display/lt174_17  (
    .a({\u2_Display/n5590 ,\u2_Display/n5591 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c17 ),
    .fco(\u2_Display/lt174_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_20|u2_Display/lt174_19  (
    .a({\u2_Display/n5588 ,\u2_Display/n5589 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c19 ),
    .fco(\u2_Display/lt174_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_22|u2_Display/lt174_21  (
    .a({\u2_Display/n5586 ,\u2_Display/n5587 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c21 ),
    .fco(\u2_Display/lt174_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_24|u2_Display/lt174_23  (
    .a({\u2_Display/n5584 ,\u2_Display/n5585 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c23 ),
    .fco(\u2_Display/lt174_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_26|u2_Display/lt174_25  (
    .a({\u2_Display/n5582 ,\u2_Display/n5583 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c25 ),
    .fco(\u2_Display/lt174_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_28|u2_Display/lt174_27  (
    .a({\u2_Display/n5580 ,\u2_Display/n5581 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c27 ),
    .fco(\u2_Display/lt174_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_2|u2_Display/lt174_1  (
    .a({\u2_Display/n5606 ,\u2_Display/n5607 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c1 ),
    .fco(\u2_Display/lt174_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_30|u2_Display/lt174_29  (
    .a({\u2_Display/n5578 ,\u2_Display/n5579 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c29 ),
    .fco(\u2_Display/lt174_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_4|u2_Display/lt174_3  (
    .a({\u2_Display/n5604 ,\u2_Display/n5605 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c3 ),
    .fco(\u2_Display/lt174_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_6|u2_Display/lt174_5  (
    .a({\u2_Display/n5602 ,\u2_Display/n5603 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c5 ),
    .fco(\u2_Display/lt174_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_8|u2_Display/lt174_7  (
    .a({\u2_Display/n5600 ,\u2_Display/n5601 }),
    .b(2'b00),
    .fci(\u2_Display/lt174_c7 ),
    .fco(\u2_Display/lt174_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt174_0|u2_Display/lt174_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt174_cout|u2_Display/lt174_31  (
    .a({1'b0,\u2_Display/n5577 }),
    .b(2'b10),
    .fci(\u2_Display/lt174_c31 ),
    .f({\u2_Display/n5609 ,open_n45653}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_0|u2_Display/lt175_cin  (
    .a({\u2_Display/n5643 ,1'b0}),
    .b({1'b0,open_n45659}),
    .fco(\u2_Display/lt175_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_10|u2_Display/lt175_9  (
    .a({\u2_Display/n5633 ,\u2_Display/n5634 }),
    .b(2'b10),
    .fci(\u2_Display/lt175_c9 ),
    .fco(\u2_Display/lt175_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_12|u2_Display/lt175_11  (
    .a({\u2_Display/n5631 ,\u2_Display/n5632 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c11 ),
    .fco(\u2_Display/lt175_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_14|u2_Display/lt175_13  (
    .a({\u2_Display/n5629 ,\u2_Display/n5630 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c13 ),
    .fco(\u2_Display/lt175_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_16|u2_Display/lt175_15  (
    .a({\u2_Display/n5627 ,\u2_Display/n5628 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c15 ),
    .fco(\u2_Display/lt175_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_18|u2_Display/lt175_17  (
    .a({\u2_Display/n5625 ,\u2_Display/n5626 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c17 ),
    .fco(\u2_Display/lt175_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_20|u2_Display/lt175_19  (
    .a({\u2_Display/n5623 ,\u2_Display/n5624 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c19 ),
    .fco(\u2_Display/lt175_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_22|u2_Display/lt175_21  (
    .a({\u2_Display/n5621 ,\u2_Display/n5622 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c21 ),
    .fco(\u2_Display/lt175_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_24|u2_Display/lt175_23  (
    .a({\u2_Display/n5619 ,\u2_Display/n5620 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c23 ),
    .fco(\u2_Display/lt175_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_26|u2_Display/lt175_25  (
    .a({\u2_Display/n5617 ,\u2_Display/n5618 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c25 ),
    .fco(\u2_Display/lt175_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_28|u2_Display/lt175_27  (
    .a({\u2_Display/n5615 ,\u2_Display/n5616 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c27 ),
    .fco(\u2_Display/lt175_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_2|u2_Display/lt175_1  (
    .a({\u2_Display/n5641 ,\u2_Display/n5642 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c1 ),
    .fco(\u2_Display/lt175_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_30|u2_Display/lt175_29  (
    .a({\u2_Display/n5613 ,\u2_Display/n5614 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c29 ),
    .fco(\u2_Display/lt175_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_4|u2_Display/lt175_3  (
    .a({\u2_Display/n5639 ,\u2_Display/n5640 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c3 ),
    .fco(\u2_Display/lt175_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_6|u2_Display/lt175_5  (
    .a({\u2_Display/n5637 ,\u2_Display/n5638 }),
    .b(2'b00),
    .fci(\u2_Display/lt175_c5 ),
    .fco(\u2_Display/lt175_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_8|u2_Display/lt175_7  (
    .a({\u2_Display/n5635 ,\u2_Display/n5636 }),
    .b(2'b10),
    .fci(\u2_Display/lt175_c7 ),
    .fco(\u2_Display/lt175_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt175_0|u2_Display/lt175_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt175_cout|u2_Display/lt175_31  (
    .a({1'b0,\u2_Display/n5612 }),
    .b(2'b10),
    .fci(\u2_Display/lt175_c31 ),
    .f({\u2_Display/n5644 ,open_n46063}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_0|u2_Display/lt176_cin  (
    .a({\u2_Display/n5678 ,1'b0}),
    .b({1'b0,open_n46069}),
    .fco(\u2_Display/lt176_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_10|u2_Display/lt176_9  (
    .a({\u2_Display/n5668 ,\u2_Display/n5669 }),
    .b(2'b01),
    .fci(\u2_Display/lt176_c9 ),
    .fco(\u2_Display/lt176_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_12|u2_Display/lt176_11  (
    .a({\u2_Display/n5666 ,\u2_Display/n5667 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c11 ),
    .fco(\u2_Display/lt176_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_14|u2_Display/lt176_13  (
    .a({\u2_Display/n5664 ,\u2_Display/n5665 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c13 ),
    .fco(\u2_Display/lt176_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_16|u2_Display/lt176_15  (
    .a({\u2_Display/n5662 ,\u2_Display/n5663 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c15 ),
    .fco(\u2_Display/lt176_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_18|u2_Display/lt176_17  (
    .a({\u2_Display/n5660 ,\u2_Display/n5661 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c17 ),
    .fco(\u2_Display/lt176_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_20|u2_Display/lt176_19  (
    .a({\u2_Display/n5658 ,\u2_Display/n5659 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c19 ),
    .fco(\u2_Display/lt176_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_22|u2_Display/lt176_21  (
    .a({\u2_Display/n5656 ,\u2_Display/n5657 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c21 ),
    .fco(\u2_Display/lt176_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_24|u2_Display/lt176_23  (
    .a({\u2_Display/n5654 ,\u2_Display/n5655 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c23 ),
    .fco(\u2_Display/lt176_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_26|u2_Display/lt176_25  (
    .a({\u2_Display/n5652 ,\u2_Display/n5653 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c25 ),
    .fco(\u2_Display/lt176_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_28|u2_Display/lt176_27  (
    .a({\u2_Display/n5650 ,\u2_Display/n5651 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c27 ),
    .fco(\u2_Display/lt176_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_2|u2_Display/lt176_1  (
    .a({\u2_Display/n5676 ,\u2_Display/n5677 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c1 ),
    .fco(\u2_Display/lt176_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_30|u2_Display/lt176_29  (
    .a({\u2_Display/n5648 ,\u2_Display/n5649 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c29 ),
    .fco(\u2_Display/lt176_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_4|u2_Display/lt176_3  (
    .a({\u2_Display/n5674 ,\u2_Display/n5675 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c3 ),
    .fco(\u2_Display/lt176_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_6|u2_Display/lt176_5  (
    .a({\u2_Display/n5672 ,\u2_Display/n5673 }),
    .b(2'b00),
    .fci(\u2_Display/lt176_c5 ),
    .fco(\u2_Display/lt176_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_8|u2_Display/lt176_7  (
    .a({\u2_Display/n5670 ,\u2_Display/n5671 }),
    .b(2'b01),
    .fci(\u2_Display/lt176_c7 ),
    .fco(\u2_Display/lt176_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt176_0|u2_Display/lt176_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt176_cout|u2_Display/lt176_31  (
    .a({1'b0,\u2_Display/n5647 }),
    .b(2'b10),
    .fci(\u2_Display/lt176_c31 ),
    .f({\u2_Display/n5679 ,open_n46473}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_0|u2_Display/lt1_cin  (
    .a({\u2_Display/i [0],1'b0}),
    .b({lcd_xpos[0],open_n46479}),
    .fco(\u2_Display/lt1_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_10|u2_Display/lt1_9  (
    .a(\u2_Display/i [10:9]),
    .b(lcd_xpos[10:9]),
    .fci(\u2_Display/lt1_c9 ),
    .fco(\u2_Display/lt1_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_2|u2_Display/lt1_1  (
    .a(\u2_Display/i [2:1]),
    .b(lcd_xpos[2:1]),
    .fci(\u2_Display/lt1_c1 ),
    .fco(\u2_Display/lt1_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_4|u2_Display/lt1_3  (
    .a(\u2_Display/i [4:3]),
    .b(lcd_xpos[4:3]),
    .fci(\u2_Display/lt1_c3 ),
    .fco(\u2_Display/lt1_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_6|u2_Display/lt1_5  (
    .a(\u2_Display/i [6:5]),
    .b(lcd_xpos[6:5]),
    .fci(\u2_Display/lt1_c5 ),
    .fco(\u2_Display/lt1_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_8|u2_Display/lt1_7  (
    .a(\u2_Display/i [8:7]),
    .b(lcd_xpos[8:7]),
    .fci(\u2_Display/lt1_c7 ),
    .fco(\u2_Display/lt1_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt1_0|u2_Display/lt1_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt1_cout|u2_Display/lt1_11  (
    .a(2'b00),
    .b({1'b1,lcd_xpos[11]}),
    .fci(\u2_Display/lt1_c11 ),
    .f({\u2_Display/n45 ,open_n46643}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_0|u2_Display/lt22_cin  (
    .a({\u2_Display/counta [0],1'b0}),
    .b({1'b0,open_n46649}),
    .fco(\u2_Display/lt22_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_10|u2_Display/lt22_9  (
    .a(\u2_Display/counta [10:9]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c9 ),
    .fco(\u2_Display/lt22_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_12|u2_Display/lt22_11  (
    .a(\u2_Display/counta [12:11]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c11 ),
    .fco(\u2_Display/lt22_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_14|u2_Display/lt22_13  (
    .a(\u2_Display/counta [14:13]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c13 ),
    .fco(\u2_Display/lt22_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_16|u2_Display/lt22_15  (
    .a(\u2_Display/counta [16:15]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c15 ),
    .fco(\u2_Display/lt22_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_18|u2_Display/lt22_17  (
    .a(\u2_Display/counta [18:17]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c17 ),
    .fco(\u2_Display/lt22_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_20|u2_Display/lt22_19  (
    .a(\u2_Display/counta [20:19]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c19 ),
    .fco(\u2_Display/lt22_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_22|u2_Display/lt22_21  (
    .a(\u2_Display/counta [22:21]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c21 ),
    .fco(\u2_Display/lt22_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_24|u2_Display/lt22_23  (
    .a(\u2_Display/counta [24:23]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c23 ),
    .fco(\u2_Display/lt22_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_26|u2_Display/lt22_25  (
    .a(\u2_Display/counta [26:25]),
    .b(2'b01),
    .fci(\u2_Display/lt22_c25 ),
    .fco(\u2_Display/lt22_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_28|u2_Display/lt22_27  (
    .a(\u2_Display/counta [28:27]),
    .b(2'b11),
    .fci(\u2_Display/lt22_c27 ),
    .fco(\u2_Display/lt22_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_2|u2_Display/lt22_1  (
    .a(\u2_Display/counta [2:1]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c1 ),
    .fco(\u2_Display/lt22_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_30|u2_Display/lt22_29  (
    .a(\u2_Display/counta [30:29]),
    .b(2'b11),
    .fci(\u2_Display/lt22_c29 ),
    .fco(\u2_Display/lt22_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_4|u2_Display/lt22_3  (
    .a(\u2_Display/counta [4:3]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c3 ),
    .fco(\u2_Display/lt22_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_6|u2_Display/lt22_5  (
    .a(\u2_Display/counta [6:5]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c5 ),
    .fco(\u2_Display/lt22_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_8|u2_Display/lt22_7  (
    .a(\u2_Display/counta [8:7]),
    .b(2'b00),
    .fci(\u2_Display/lt22_c7 ),
    .fco(\u2_Display/lt22_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt22_0|u2_Display/lt22_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt22_cout|u2_Display/lt22_31  (
    .a({1'b0,\u2_Display/counta [31]}),
    .b(2'b11),
    .fci(\u2_Display/lt22_c31 ),
    .f({\u2_Display/n417 ,open_n47053}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_0|u2_Display/lt23_cin  (
    .a({\u2_Display/n451 ,1'b0}),
    .b({1'b0,open_n47059}),
    .fco(\u2_Display/lt23_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_10|u2_Display/lt23_9  (
    .a({\u2_Display/n441 ,\u2_Display/n442 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c9 ),
    .fco(\u2_Display/lt23_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_12|u2_Display/lt23_11  (
    .a({\u2_Display/n439 ,\u2_Display/n440 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c11 ),
    .fco(\u2_Display/lt23_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_14|u2_Display/lt23_13  (
    .a({\u2_Display/n437 ,\u2_Display/n438 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c13 ),
    .fco(\u2_Display/lt23_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_16|u2_Display/lt23_15  (
    .a({\u2_Display/n435 ,\u2_Display/n436 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c15 ),
    .fco(\u2_Display/lt23_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_18|u2_Display/lt23_17  (
    .a({\u2_Display/n433 ,\u2_Display/n434 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c17 ),
    .fco(\u2_Display/lt23_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_20|u2_Display/lt23_19  (
    .a({\u2_Display/n431 ,\u2_Display/n432 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c19 ),
    .fco(\u2_Display/lt23_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_22|u2_Display/lt23_21  (
    .a({\u2_Display/n429 ,\u2_Display/n430 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c21 ),
    .fco(\u2_Display/lt23_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_24|u2_Display/lt23_23  (
    .a({\u2_Display/n427 ,\u2_Display/n428 }),
    .b(2'b10),
    .fci(\u2_Display/lt23_c23 ),
    .fco(\u2_Display/lt23_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_26|u2_Display/lt23_25  (
    .a({\u2_Display/n425 ,\u2_Display/n426 }),
    .b(2'b10),
    .fci(\u2_Display/lt23_c25 ),
    .fco(\u2_Display/lt23_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_28|u2_Display/lt23_27  (
    .a({\u2_Display/n423 ,\u2_Display/n424 }),
    .b(2'b11),
    .fci(\u2_Display/lt23_c27 ),
    .fco(\u2_Display/lt23_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_2|u2_Display/lt23_1  (
    .a({\u2_Display/n449 ,\u2_Display/n450 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c1 ),
    .fco(\u2_Display/lt23_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_30|u2_Display/lt23_29  (
    .a({\u2_Display/n421 ,\u2_Display/n422 }),
    .b(2'b11),
    .fci(\u2_Display/lt23_c29 ),
    .fco(\u2_Display/lt23_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_4|u2_Display/lt23_3  (
    .a({\u2_Display/n447 ,\u2_Display/n448 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c3 ),
    .fco(\u2_Display/lt23_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_6|u2_Display/lt23_5  (
    .a({\u2_Display/n445 ,\u2_Display/n446 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c5 ),
    .fco(\u2_Display/lt23_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_8|u2_Display/lt23_7  (
    .a({\u2_Display/n443 ,\u2_Display/n444 }),
    .b(2'b00),
    .fci(\u2_Display/lt23_c7 ),
    .fco(\u2_Display/lt23_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt23_0|u2_Display/lt23_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt23_cout|u2_Display/lt23_31  (
    .a({1'b0,\u2_Display/n420 }),
    .b(2'b10),
    .fci(\u2_Display/lt23_c31 ),
    .f({\u2_Display/n452 ,open_n47463}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_0|u2_Display/lt24_cin  (
    .a({\u2_Display/n486 ,1'b0}),
    .b({1'b0,open_n47469}),
    .fco(\u2_Display/lt24_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_10|u2_Display/lt24_9  (
    .a({\u2_Display/n476 ,\u2_Display/n477 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c9 ),
    .fco(\u2_Display/lt24_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_12|u2_Display/lt24_11  (
    .a({\u2_Display/n474 ,\u2_Display/n475 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c11 ),
    .fco(\u2_Display/lt24_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_14|u2_Display/lt24_13  (
    .a({\u2_Display/n472 ,\u2_Display/n473 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c13 ),
    .fco(\u2_Display/lt24_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_16|u2_Display/lt24_15  (
    .a({\u2_Display/n470 ,\u2_Display/n471 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c15 ),
    .fco(\u2_Display/lt24_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_18|u2_Display/lt24_17  (
    .a({\u2_Display/n468 ,\u2_Display/n469 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c17 ),
    .fco(\u2_Display/lt24_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_20|u2_Display/lt24_19  (
    .a({\u2_Display/n466 ,\u2_Display/n467 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c19 ),
    .fco(\u2_Display/lt24_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_22|u2_Display/lt24_21  (
    .a({\u2_Display/n464 ,\u2_Display/n465 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c21 ),
    .fco(\u2_Display/lt24_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_24|u2_Display/lt24_23  (
    .a({\u2_Display/n462 ,\u2_Display/n463 }),
    .b(2'b01),
    .fci(\u2_Display/lt24_c23 ),
    .fco(\u2_Display/lt24_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_26|u2_Display/lt24_25  (
    .a({\u2_Display/n460 ,\u2_Display/n461 }),
    .b(2'b11),
    .fci(\u2_Display/lt24_c25 ),
    .fco(\u2_Display/lt24_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_28|u2_Display/lt24_27  (
    .a({\u2_Display/n458 ,\u2_Display/n459 }),
    .b(2'b11),
    .fci(\u2_Display/lt24_c27 ),
    .fco(\u2_Display/lt24_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_2|u2_Display/lt24_1  (
    .a({\u2_Display/n484 ,\u2_Display/n485 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c1 ),
    .fco(\u2_Display/lt24_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_30|u2_Display/lt24_29  (
    .a({\u2_Display/n456 ,\u2_Display/n457 }),
    .b(2'b01),
    .fci(\u2_Display/lt24_c29 ),
    .fco(\u2_Display/lt24_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_4|u2_Display/lt24_3  (
    .a({\u2_Display/n482 ,\u2_Display/n483 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c3 ),
    .fco(\u2_Display/lt24_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_6|u2_Display/lt24_5  (
    .a({\u2_Display/n480 ,\u2_Display/n481 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c5 ),
    .fco(\u2_Display/lt24_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_8|u2_Display/lt24_7  (
    .a({\u2_Display/n478 ,\u2_Display/n479 }),
    .b(2'b00),
    .fci(\u2_Display/lt24_c7 ),
    .fco(\u2_Display/lt24_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt24_0|u2_Display/lt24_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt24_cout|u2_Display/lt24_31  (
    .a({1'b0,\u2_Display/n455 }),
    .b(2'b10),
    .fci(\u2_Display/lt24_c31 ),
    .f({\u2_Display/n487 ,open_n47873}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_0|u2_Display/lt25_cin  (
    .a({\u2_Display/n521 ,1'b0}),
    .b({1'b0,open_n47879}),
    .fco(\u2_Display/lt25_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_10|u2_Display/lt25_9  (
    .a({\u2_Display/n511 ,\u2_Display/n512 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c9 ),
    .fco(\u2_Display/lt25_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_12|u2_Display/lt25_11  (
    .a({\u2_Display/n509 ,\u2_Display/n510 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c11 ),
    .fco(\u2_Display/lt25_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_14|u2_Display/lt25_13  (
    .a({\u2_Display/n507 ,\u2_Display/n508 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c13 ),
    .fco(\u2_Display/lt25_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_16|u2_Display/lt25_15  (
    .a({\u2_Display/n505 ,\u2_Display/n506 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c15 ),
    .fco(\u2_Display/lt25_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_18|u2_Display/lt25_17  (
    .a({\u2_Display/n503 ,\u2_Display/n504 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c17 ),
    .fco(\u2_Display/lt25_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_20|u2_Display/lt25_19  (
    .a({\u2_Display/n501 ,\u2_Display/n502 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c19 ),
    .fco(\u2_Display/lt25_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_22|u2_Display/lt25_21  (
    .a({\u2_Display/n499 ,\u2_Display/n500 }),
    .b(2'b10),
    .fci(\u2_Display/lt25_c21 ),
    .fco(\u2_Display/lt25_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_24|u2_Display/lt25_23  (
    .a({\u2_Display/n497 ,\u2_Display/n498 }),
    .b(2'b10),
    .fci(\u2_Display/lt25_c23 ),
    .fco(\u2_Display/lt25_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_26|u2_Display/lt25_25  (
    .a({\u2_Display/n495 ,\u2_Display/n496 }),
    .b(2'b11),
    .fci(\u2_Display/lt25_c25 ),
    .fco(\u2_Display/lt25_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_28|u2_Display/lt25_27  (
    .a({\u2_Display/n493 ,\u2_Display/n494 }),
    .b(2'b11),
    .fci(\u2_Display/lt25_c27 ),
    .fco(\u2_Display/lt25_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_2|u2_Display/lt25_1  (
    .a({\u2_Display/n519 ,\u2_Display/n520 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c1 ),
    .fco(\u2_Display/lt25_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_30|u2_Display/lt25_29  (
    .a({\u2_Display/n491 ,\u2_Display/n492 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c29 ),
    .fco(\u2_Display/lt25_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_4|u2_Display/lt25_3  (
    .a({\u2_Display/n517 ,\u2_Display/n518 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c3 ),
    .fco(\u2_Display/lt25_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_6|u2_Display/lt25_5  (
    .a({\u2_Display/n515 ,\u2_Display/n516 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c5 ),
    .fco(\u2_Display/lt25_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_8|u2_Display/lt25_7  (
    .a({\u2_Display/n513 ,\u2_Display/n514 }),
    .b(2'b00),
    .fci(\u2_Display/lt25_c7 ),
    .fco(\u2_Display/lt25_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt25_0|u2_Display/lt25_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt25_cout|u2_Display/lt25_31  (
    .a({1'b0,\u2_Display/n490 }),
    .b(2'b10),
    .fci(\u2_Display/lt25_c31 ),
    .f({\u2_Display/n522 ,open_n48283}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_0|u2_Display/lt26_cin  (
    .a({\u2_Display/n556 ,1'b0}),
    .b({1'b0,open_n48289}),
    .fco(\u2_Display/lt26_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_10|u2_Display/lt26_9  (
    .a({\u2_Display/n546 ,\u2_Display/n547 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c9 ),
    .fco(\u2_Display/lt26_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_12|u2_Display/lt26_11  (
    .a({\u2_Display/n544 ,\u2_Display/n545 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c11 ),
    .fco(\u2_Display/lt26_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_14|u2_Display/lt26_13  (
    .a({\u2_Display/n542 ,\u2_Display/n543 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c13 ),
    .fco(\u2_Display/lt26_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_16|u2_Display/lt26_15  (
    .a({\u2_Display/n540 ,\u2_Display/n541 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c15 ),
    .fco(\u2_Display/lt26_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_18|u2_Display/lt26_17  (
    .a({\u2_Display/n538 ,\u2_Display/n539 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c17 ),
    .fco(\u2_Display/lt26_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_20|u2_Display/lt26_19  (
    .a({\u2_Display/n536 ,\u2_Display/n537 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c19 ),
    .fco(\u2_Display/lt26_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_22|u2_Display/lt26_21  (
    .a({\u2_Display/n534 ,\u2_Display/n535 }),
    .b(2'b01),
    .fci(\u2_Display/lt26_c21 ),
    .fco(\u2_Display/lt26_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_24|u2_Display/lt26_23  (
    .a({\u2_Display/n532 ,\u2_Display/n533 }),
    .b(2'b11),
    .fci(\u2_Display/lt26_c23 ),
    .fco(\u2_Display/lt26_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_26|u2_Display/lt26_25  (
    .a({\u2_Display/n530 ,\u2_Display/n531 }),
    .b(2'b11),
    .fci(\u2_Display/lt26_c25 ),
    .fco(\u2_Display/lt26_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_28|u2_Display/lt26_27  (
    .a({\u2_Display/n528 ,\u2_Display/n529 }),
    .b(2'b01),
    .fci(\u2_Display/lt26_c27 ),
    .fco(\u2_Display/lt26_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_2|u2_Display/lt26_1  (
    .a({\u2_Display/n554 ,\u2_Display/n555 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c1 ),
    .fco(\u2_Display/lt26_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_30|u2_Display/lt26_29  (
    .a({\u2_Display/n526 ,\u2_Display/n527 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c29 ),
    .fco(\u2_Display/lt26_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_4|u2_Display/lt26_3  (
    .a({\u2_Display/n552 ,\u2_Display/n553 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c3 ),
    .fco(\u2_Display/lt26_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_6|u2_Display/lt26_5  (
    .a({\u2_Display/n550 ,\u2_Display/n551 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c5 ),
    .fco(\u2_Display/lt26_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_8|u2_Display/lt26_7  (
    .a({\u2_Display/n548 ,\u2_Display/n549 }),
    .b(2'b00),
    .fci(\u2_Display/lt26_c7 ),
    .fco(\u2_Display/lt26_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt26_0|u2_Display/lt26_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt26_cout|u2_Display/lt26_31  (
    .a({1'b0,\u2_Display/n525 }),
    .b(2'b10),
    .fci(\u2_Display/lt26_c31 ),
    .f({\u2_Display/n557 ,open_n48693}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_0|u2_Display/lt27_cin  (
    .a({\u2_Display/n591 ,1'b0}),
    .b({1'b0,open_n48699}),
    .fco(\u2_Display/lt27_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_10|u2_Display/lt27_9  (
    .a({\u2_Display/n581 ,\u2_Display/n582 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c9 ),
    .fco(\u2_Display/lt27_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_12|u2_Display/lt27_11  (
    .a({\u2_Display/n579 ,\u2_Display/n580 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c11 ),
    .fco(\u2_Display/lt27_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_14|u2_Display/lt27_13  (
    .a({\u2_Display/n577 ,\u2_Display/n578 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c13 ),
    .fco(\u2_Display/lt27_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_16|u2_Display/lt27_15  (
    .a({\u2_Display/n575 ,\u2_Display/n576 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c15 ),
    .fco(\u2_Display/lt27_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_18|u2_Display/lt27_17  (
    .a({\u2_Display/n573 ,\u2_Display/n574 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c17 ),
    .fco(\u2_Display/lt27_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_20|u2_Display/lt27_19  (
    .a({\u2_Display/n571 ,\u2_Display/n572 }),
    .b(2'b10),
    .fci(\u2_Display/lt27_c19 ),
    .fco(\u2_Display/lt27_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_22|u2_Display/lt27_21  (
    .a({\u2_Display/n569 ,\u2_Display/n570 }),
    .b(2'b10),
    .fci(\u2_Display/lt27_c21 ),
    .fco(\u2_Display/lt27_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_24|u2_Display/lt27_23  (
    .a({\u2_Display/n567 ,\u2_Display/n568 }),
    .b(2'b11),
    .fci(\u2_Display/lt27_c23 ),
    .fco(\u2_Display/lt27_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_26|u2_Display/lt27_25  (
    .a({\u2_Display/n565 ,\u2_Display/n566 }),
    .b(2'b11),
    .fci(\u2_Display/lt27_c25 ),
    .fco(\u2_Display/lt27_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_28|u2_Display/lt27_27  (
    .a({\u2_Display/n563 ,\u2_Display/n564 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c27 ),
    .fco(\u2_Display/lt27_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_2|u2_Display/lt27_1  (
    .a({\u2_Display/n589 ,\u2_Display/n590 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c1 ),
    .fco(\u2_Display/lt27_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_30|u2_Display/lt27_29  (
    .a({\u2_Display/n561 ,\u2_Display/n562 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c29 ),
    .fco(\u2_Display/lt27_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_4|u2_Display/lt27_3  (
    .a({\u2_Display/n587 ,\u2_Display/n588 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c3 ),
    .fco(\u2_Display/lt27_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_6|u2_Display/lt27_5  (
    .a({\u2_Display/n585 ,\u2_Display/n586 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c5 ),
    .fco(\u2_Display/lt27_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_8|u2_Display/lt27_7  (
    .a({\u2_Display/n583 ,\u2_Display/n584 }),
    .b(2'b00),
    .fci(\u2_Display/lt27_c7 ),
    .fco(\u2_Display/lt27_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt27_0|u2_Display/lt27_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt27_cout|u2_Display/lt27_31  (
    .a({1'b0,\u2_Display/n560 }),
    .b(2'b10),
    .fci(\u2_Display/lt27_c31 ),
    .f({\u2_Display/n592 ,open_n49103}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_0|u2_Display/lt28_cin  (
    .a({\u2_Display/n626 ,1'b0}),
    .b({1'b0,open_n49109}),
    .fco(\u2_Display/lt28_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_10|u2_Display/lt28_9  (
    .a({\u2_Display/n616 ,\u2_Display/n617 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c9 ),
    .fco(\u2_Display/lt28_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_12|u2_Display/lt28_11  (
    .a({\u2_Display/n614 ,\u2_Display/n615 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c11 ),
    .fco(\u2_Display/lt28_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_14|u2_Display/lt28_13  (
    .a({\u2_Display/n612 ,\u2_Display/n613 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c13 ),
    .fco(\u2_Display/lt28_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_16|u2_Display/lt28_15  (
    .a({\u2_Display/n610 ,\u2_Display/n611 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c15 ),
    .fco(\u2_Display/lt28_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_18|u2_Display/lt28_17  (
    .a({\u2_Display/n608 ,\u2_Display/n609 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c17 ),
    .fco(\u2_Display/lt28_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_20|u2_Display/lt28_19  (
    .a({\u2_Display/n606 ,\u2_Display/n607 }),
    .b(2'b01),
    .fci(\u2_Display/lt28_c19 ),
    .fco(\u2_Display/lt28_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_22|u2_Display/lt28_21  (
    .a({\u2_Display/n604 ,\u2_Display/n605 }),
    .b(2'b11),
    .fci(\u2_Display/lt28_c21 ),
    .fco(\u2_Display/lt28_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_24|u2_Display/lt28_23  (
    .a({\u2_Display/n602 ,\u2_Display/n603 }),
    .b(2'b11),
    .fci(\u2_Display/lt28_c23 ),
    .fco(\u2_Display/lt28_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_26|u2_Display/lt28_25  (
    .a({\u2_Display/n600 ,\u2_Display/n601 }),
    .b(2'b01),
    .fci(\u2_Display/lt28_c25 ),
    .fco(\u2_Display/lt28_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_28|u2_Display/lt28_27  (
    .a({\u2_Display/n598 ,\u2_Display/n599 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c27 ),
    .fco(\u2_Display/lt28_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_2|u2_Display/lt28_1  (
    .a({\u2_Display/n624 ,\u2_Display/n625 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c1 ),
    .fco(\u2_Display/lt28_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_30|u2_Display/lt28_29  (
    .a({\u2_Display/n596 ,\u2_Display/n597 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c29 ),
    .fco(\u2_Display/lt28_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_4|u2_Display/lt28_3  (
    .a({\u2_Display/n622 ,\u2_Display/n623 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c3 ),
    .fco(\u2_Display/lt28_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_6|u2_Display/lt28_5  (
    .a({\u2_Display/n620 ,\u2_Display/n621 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c5 ),
    .fco(\u2_Display/lt28_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_8|u2_Display/lt28_7  (
    .a({\u2_Display/n618 ,\u2_Display/n619 }),
    .b(2'b00),
    .fci(\u2_Display/lt28_c7 ),
    .fco(\u2_Display/lt28_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt28_0|u2_Display/lt28_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt28_cout|u2_Display/lt28_31  (
    .a({1'b0,\u2_Display/n595 }),
    .b(2'b10),
    .fci(\u2_Display/lt28_c31 ),
    .f({\u2_Display/n627 ,open_n49513}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_0|u2_Display/lt29_cin  (
    .a({\u2_Display/n661 ,1'b0}),
    .b({1'b0,open_n49519}),
    .fco(\u2_Display/lt29_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_10|u2_Display/lt29_9  (
    .a({\u2_Display/n651 ,\u2_Display/n652 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c9 ),
    .fco(\u2_Display/lt29_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_12|u2_Display/lt29_11  (
    .a({\u2_Display/n649 ,\u2_Display/n650 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c11 ),
    .fco(\u2_Display/lt29_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_14|u2_Display/lt29_13  (
    .a({\u2_Display/n647 ,\u2_Display/n648 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c13 ),
    .fco(\u2_Display/lt29_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_16|u2_Display/lt29_15  (
    .a({\u2_Display/n645 ,\u2_Display/n646 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c15 ),
    .fco(\u2_Display/lt29_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_18|u2_Display/lt29_17  (
    .a({\u2_Display/n643 ,\u2_Display/n644 }),
    .b(2'b10),
    .fci(\u2_Display/lt29_c17 ),
    .fco(\u2_Display/lt29_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_20|u2_Display/lt29_19  (
    .a({\u2_Display/n641 ,\u2_Display/n642 }),
    .b(2'b10),
    .fci(\u2_Display/lt29_c19 ),
    .fco(\u2_Display/lt29_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_22|u2_Display/lt29_21  (
    .a({\u2_Display/n639 ,\u2_Display/n640 }),
    .b(2'b11),
    .fci(\u2_Display/lt29_c21 ),
    .fco(\u2_Display/lt29_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_24|u2_Display/lt29_23  (
    .a({\u2_Display/n637 ,\u2_Display/n638 }),
    .b(2'b11),
    .fci(\u2_Display/lt29_c23 ),
    .fco(\u2_Display/lt29_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_26|u2_Display/lt29_25  (
    .a({\u2_Display/n635 ,\u2_Display/n636 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c25 ),
    .fco(\u2_Display/lt29_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_28|u2_Display/lt29_27  (
    .a({\u2_Display/n633 ,\u2_Display/n634 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c27 ),
    .fco(\u2_Display/lt29_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_2|u2_Display/lt29_1  (
    .a({\u2_Display/n659 ,\u2_Display/n660 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c1 ),
    .fco(\u2_Display/lt29_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_30|u2_Display/lt29_29  (
    .a({\u2_Display/n631 ,\u2_Display/n632 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c29 ),
    .fco(\u2_Display/lt29_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_4|u2_Display/lt29_3  (
    .a({\u2_Display/n657 ,\u2_Display/n658 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c3 ),
    .fco(\u2_Display/lt29_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_6|u2_Display/lt29_5  (
    .a({\u2_Display/n655 ,\u2_Display/n656 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c5 ),
    .fco(\u2_Display/lt29_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_8|u2_Display/lt29_7  (
    .a({\u2_Display/n653 ,\u2_Display/n654 }),
    .b(2'b00),
    .fci(\u2_Display/lt29_c7 ),
    .fco(\u2_Display/lt29_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt29_0|u2_Display/lt29_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt29_cout|u2_Display/lt29_31  (
    .a({1'b0,\u2_Display/n630 }),
    .b(2'b10),
    .fci(\u2_Display/lt29_c31 ),
    .f({\u2_Display/n662 ,open_n49923}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_0|u2_Display/lt2_2_cin  (
    .a({lcd_ypos[0],1'b0}),
    .b({\u2_Display/j [0],open_n49929}),
    .fco(\u2_Display/lt2_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_10|u2_Display/lt2_2_9  (
    .a(lcd_ypos[10:9]),
    .b({1'b1,\u2_Display/j [9]}),
    .fci(\u2_Display/lt2_2_c9 ),
    .fco(\u2_Display/lt2_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_2|u2_Display/lt2_2_1  (
    .a(lcd_ypos[2:1]),
    .b(\u2_Display/j [2:1]),
    .fci(\u2_Display/lt2_2_c1 ),
    .fco(\u2_Display/lt2_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_4|u2_Display/lt2_2_3  (
    .a(lcd_ypos[4:3]),
    .b(\u2_Display/j [4:3]),
    .fci(\u2_Display/lt2_2_c3 ),
    .fco(\u2_Display/lt2_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_6|u2_Display/lt2_2_5  (
    .a(lcd_ypos[6:5]),
    .b(\u2_Display/j [6:5]),
    .fci(\u2_Display/lt2_2_c5 ),
    .fco(\u2_Display/lt2_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_8|u2_Display/lt2_2_7  (
    .a(lcd_ypos[8:7]),
    .b(\u2_Display/j [8:7]),
    .fci(\u2_Display/lt2_2_c7 ),
    .fco(\u2_Display/lt2_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt2_2_0|u2_Display/lt2_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt2_2_cout|u2_Display/lt2_2_11  (
    .a({1'b0,lcd_ypos[11]}),
    .b(2'b10),
    .fci(\u2_Display/lt2_2_c11 ),
    .f({\u2_Display/n48 ,open_n50093}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_0|u2_Display/lt30_cin  (
    .a({\u2_Display/n696 ,1'b0}),
    .b({1'b0,open_n50099}),
    .fco(\u2_Display/lt30_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_10|u2_Display/lt30_9  (
    .a({\u2_Display/n686 ,\u2_Display/n687 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c9 ),
    .fco(\u2_Display/lt30_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_12|u2_Display/lt30_11  (
    .a({\u2_Display/n684 ,\u2_Display/n685 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c11 ),
    .fco(\u2_Display/lt30_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_14|u2_Display/lt30_13  (
    .a({\u2_Display/n682 ,\u2_Display/n683 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c13 ),
    .fco(\u2_Display/lt30_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_16|u2_Display/lt30_15  (
    .a({\u2_Display/n680 ,\u2_Display/n681 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c15 ),
    .fco(\u2_Display/lt30_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_18|u2_Display/lt30_17  (
    .a({\u2_Display/n678 ,\u2_Display/n679 }),
    .b(2'b01),
    .fci(\u2_Display/lt30_c17 ),
    .fco(\u2_Display/lt30_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_20|u2_Display/lt30_19  (
    .a({\u2_Display/n676 ,\u2_Display/n677 }),
    .b(2'b11),
    .fci(\u2_Display/lt30_c19 ),
    .fco(\u2_Display/lt30_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_22|u2_Display/lt30_21  (
    .a({\u2_Display/n674 ,\u2_Display/n675 }),
    .b(2'b11),
    .fci(\u2_Display/lt30_c21 ),
    .fco(\u2_Display/lt30_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_24|u2_Display/lt30_23  (
    .a({\u2_Display/n672 ,\u2_Display/n673 }),
    .b(2'b01),
    .fci(\u2_Display/lt30_c23 ),
    .fco(\u2_Display/lt30_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_26|u2_Display/lt30_25  (
    .a({\u2_Display/n670 ,\u2_Display/n671 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c25 ),
    .fco(\u2_Display/lt30_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_28|u2_Display/lt30_27  (
    .a({\u2_Display/n668 ,\u2_Display/n669 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c27 ),
    .fco(\u2_Display/lt30_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_2|u2_Display/lt30_1  (
    .a({\u2_Display/n694 ,\u2_Display/n695 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c1 ),
    .fco(\u2_Display/lt30_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_30|u2_Display/lt30_29  (
    .a({\u2_Display/n666 ,\u2_Display/n667 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c29 ),
    .fco(\u2_Display/lt30_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_4|u2_Display/lt30_3  (
    .a({\u2_Display/n692 ,\u2_Display/n693 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c3 ),
    .fco(\u2_Display/lt30_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_6|u2_Display/lt30_5  (
    .a({\u2_Display/n690 ,\u2_Display/n691 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c5 ),
    .fco(\u2_Display/lt30_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_8|u2_Display/lt30_7  (
    .a({\u2_Display/n688 ,\u2_Display/n689 }),
    .b(2'b00),
    .fci(\u2_Display/lt30_c7 ),
    .fco(\u2_Display/lt30_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt30_0|u2_Display/lt30_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt30_cout|u2_Display/lt30_31  (
    .a({1'b0,\u2_Display/n665 }),
    .b(2'b10),
    .fci(\u2_Display/lt30_c31 ),
    .f({\u2_Display/n697 ,open_n50503}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_0|u2_Display/lt31_cin  (
    .a({\u2_Display/n731 ,1'b0}),
    .b({1'b0,open_n50509}),
    .fco(\u2_Display/lt31_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_10|u2_Display/lt31_9  (
    .a({\u2_Display/n721 ,\u2_Display/n722 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c9 ),
    .fco(\u2_Display/lt31_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_12|u2_Display/lt31_11  (
    .a({\u2_Display/n719 ,\u2_Display/n720 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c11 ),
    .fco(\u2_Display/lt31_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_14|u2_Display/lt31_13  (
    .a({\u2_Display/n717 ,\u2_Display/n718 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c13 ),
    .fco(\u2_Display/lt31_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_16|u2_Display/lt31_15  (
    .a({\u2_Display/n715 ,\u2_Display/n716 }),
    .b(2'b10),
    .fci(\u2_Display/lt31_c15 ),
    .fco(\u2_Display/lt31_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_18|u2_Display/lt31_17  (
    .a({\u2_Display/n713 ,\u2_Display/n714 }),
    .b(2'b10),
    .fci(\u2_Display/lt31_c17 ),
    .fco(\u2_Display/lt31_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_20|u2_Display/lt31_19  (
    .a({\u2_Display/n711 ,\u2_Display/n712 }),
    .b(2'b11),
    .fci(\u2_Display/lt31_c19 ),
    .fco(\u2_Display/lt31_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_22|u2_Display/lt31_21  (
    .a({\u2_Display/n709 ,\u2_Display/n710 }),
    .b(2'b11),
    .fci(\u2_Display/lt31_c21 ),
    .fco(\u2_Display/lt31_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_24|u2_Display/lt31_23  (
    .a({\u2_Display/n707 ,\u2_Display/n708 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c23 ),
    .fco(\u2_Display/lt31_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_26|u2_Display/lt31_25  (
    .a({\u2_Display/n705 ,\u2_Display/n706 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c25 ),
    .fco(\u2_Display/lt31_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_28|u2_Display/lt31_27  (
    .a({\u2_Display/n703 ,\u2_Display/n704 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c27 ),
    .fco(\u2_Display/lt31_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_2|u2_Display/lt31_1  (
    .a({\u2_Display/n729 ,\u2_Display/n730 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c1 ),
    .fco(\u2_Display/lt31_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_30|u2_Display/lt31_29  (
    .a({\u2_Display/n701 ,\u2_Display/n702 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c29 ),
    .fco(\u2_Display/lt31_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_4|u2_Display/lt31_3  (
    .a({\u2_Display/n727 ,\u2_Display/n728 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c3 ),
    .fco(\u2_Display/lt31_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_6|u2_Display/lt31_5  (
    .a({\u2_Display/n725 ,\u2_Display/n726 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c5 ),
    .fco(\u2_Display/lt31_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_8|u2_Display/lt31_7  (
    .a({\u2_Display/n723 ,\u2_Display/n724 }),
    .b(2'b00),
    .fci(\u2_Display/lt31_c7 ),
    .fco(\u2_Display/lt31_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt31_0|u2_Display/lt31_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt31_cout|u2_Display/lt31_31  (
    .a({1'b0,\u2_Display/n700 }),
    .b(2'b10),
    .fci(\u2_Display/lt31_c31 ),
    .f({\u2_Display/n732 ,open_n50913}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_0|u2_Display/lt32_cin  (
    .a({\u2_Display/n766 ,1'b0}),
    .b({1'b0,open_n50919}),
    .fco(\u2_Display/lt32_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_10|u2_Display/lt32_9  (
    .a({\u2_Display/n756 ,\u2_Display/n757 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c9 ),
    .fco(\u2_Display/lt32_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_12|u2_Display/lt32_11  (
    .a({\u2_Display/n754 ,\u2_Display/n755 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c11 ),
    .fco(\u2_Display/lt32_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_14|u2_Display/lt32_13  (
    .a({\u2_Display/n752 ,\u2_Display/n753 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c13 ),
    .fco(\u2_Display/lt32_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_16|u2_Display/lt32_15  (
    .a({\u2_Display/n750 ,\u2_Display/n751 }),
    .b(2'b01),
    .fci(\u2_Display/lt32_c15 ),
    .fco(\u2_Display/lt32_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_18|u2_Display/lt32_17  (
    .a({\u2_Display/n748 ,\u2_Display/n749 }),
    .b(2'b11),
    .fci(\u2_Display/lt32_c17 ),
    .fco(\u2_Display/lt32_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_20|u2_Display/lt32_19  (
    .a({\u2_Display/n746 ,\u2_Display/n747 }),
    .b(2'b11),
    .fci(\u2_Display/lt32_c19 ),
    .fco(\u2_Display/lt32_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_22|u2_Display/lt32_21  (
    .a({\u2_Display/n744 ,\u2_Display/n745 }),
    .b(2'b01),
    .fci(\u2_Display/lt32_c21 ),
    .fco(\u2_Display/lt32_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_24|u2_Display/lt32_23  (
    .a({\u2_Display/n742 ,\u2_Display/n743 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c23 ),
    .fco(\u2_Display/lt32_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_26|u2_Display/lt32_25  (
    .a({\u2_Display/n740 ,\u2_Display/n741 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c25 ),
    .fco(\u2_Display/lt32_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_28|u2_Display/lt32_27  (
    .a({\u2_Display/n738 ,\u2_Display/n739 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c27 ),
    .fco(\u2_Display/lt32_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_2|u2_Display/lt32_1  (
    .a({\u2_Display/n764 ,\u2_Display/n765 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c1 ),
    .fco(\u2_Display/lt32_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_30|u2_Display/lt32_29  (
    .a({\u2_Display/n736 ,\u2_Display/n737 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c29 ),
    .fco(\u2_Display/lt32_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_4|u2_Display/lt32_3  (
    .a({\u2_Display/n762 ,\u2_Display/n763 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c3 ),
    .fco(\u2_Display/lt32_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_6|u2_Display/lt32_5  (
    .a({\u2_Display/n760 ,\u2_Display/n761 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c5 ),
    .fco(\u2_Display/lt32_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_8|u2_Display/lt32_7  (
    .a({\u2_Display/n758 ,\u2_Display/n759 }),
    .b(2'b00),
    .fci(\u2_Display/lt32_c7 ),
    .fco(\u2_Display/lt32_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt32_0|u2_Display/lt32_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt32_cout|u2_Display/lt32_31  (
    .a({1'b0,\u2_Display/n735 }),
    .b(2'b10),
    .fci(\u2_Display/lt32_c31 ),
    .f({\u2_Display/n767 ,open_n51323}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_0|u2_Display/lt33_cin  (
    .a({\u2_Display/n801 ,1'b0}),
    .b({1'b0,open_n51329}),
    .fco(\u2_Display/lt33_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_10|u2_Display/lt33_9  (
    .a({\u2_Display/n791 ,\u2_Display/n792 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c9 ),
    .fco(\u2_Display/lt33_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_12|u2_Display/lt33_11  (
    .a({\u2_Display/n789 ,\u2_Display/n790 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c11 ),
    .fco(\u2_Display/lt33_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_14|u2_Display/lt33_13  (
    .a({\u2_Display/n787 ,\u2_Display/n788 }),
    .b(2'b10),
    .fci(\u2_Display/lt33_c13 ),
    .fco(\u2_Display/lt33_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_16|u2_Display/lt33_15  (
    .a({\u2_Display/n785 ,\u2_Display/n786 }),
    .b(2'b10),
    .fci(\u2_Display/lt33_c15 ),
    .fco(\u2_Display/lt33_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_18|u2_Display/lt33_17  (
    .a({\u2_Display/n783 ,\u2_Display/n784 }),
    .b(2'b11),
    .fci(\u2_Display/lt33_c17 ),
    .fco(\u2_Display/lt33_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_20|u2_Display/lt33_19  (
    .a({\u2_Display/n781 ,\u2_Display/n782 }),
    .b(2'b11),
    .fci(\u2_Display/lt33_c19 ),
    .fco(\u2_Display/lt33_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_22|u2_Display/lt33_21  (
    .a({\u2_Display/n779 ,\u2_Display/n780 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c21 ),
    .fco(\u2_Display/lt33_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_24|u2_Display/lt33_23  (
    .a({\u2_Display/n777 ,\u2_Display/n778 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c23 ),
    .fco(\u2_Display/lt33_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_26|u2_Display/lt33_25  (
    .a({\u2_Display/n775 ,\u2_Display/n776 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c25 ),
    .fco(\u2_Display/lt33_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_28|u2_Display/lt33_27  (
    .a({\u2_Display/n773 ,\u2_Display/n774 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c27 ),
    .fco(\u2_Display/lt33_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_2|u2_Display/lt33_1  (
    .a({\u2_Display/n799 ,\u2_Display/n800 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c1 ),
    .fco(\u2_Display/lt33_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_30|u2_Display/lt33_29  (
    .a({\u2_Display/n771 ,\u2_Display/n772 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c29 ),
    .fco(\u2_Display/lt33_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_4|u2_Display/lt33_3  (
    .a({\u2_Display/n797 ,\u2_Display/n798 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c3 ),
    .fco(\u2_Display/lt33_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_6|u2_Display/lt33_5  (
    .a({\u2_Display/n795 ,\u2_Display/n796 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c5 ),
    .fco(\u2_Display/lt33_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_8|u2_Display/lt33_7  (
    .a({\u2_Display/n793 ,\u2_Display/n794 }),
    .b(2'b00),
    .fci(\u2_Display/lt33_c7 ),
    .fco(\u2_Display/lt33_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt33_0|u2_Display/lt33_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt33_cout|u2_Display/lt33_31  (
    .a({1'b0,\u2_Display/n770 }),
    .b(2'b10),
    .fci(\u2_Display/lt33_c31 ),
    .f({\u2_Display/n802 ,open_n51733}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_0|u2_Display/lt34_cin  (
    .a({\u2_Display/n836 ,1'b0}),
    .b({1'b0,open_n51739}),
    .fco(\u2_Display/lt34_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_10|u2_Display/lt34_9  (
    .a({\u2_Display/n826 ,\u2_Display/n827 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c9 ),
    .fco(\u2_Display/lt34_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_12|u2_Display/lt34_11  (
    .a({\u2_Display/n824 ,\u2_Display/n825 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c11 ),
    .fco(\u2_Display/lt34_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_14|u2_Display/lt34_13  (
    .a({\u2_Display/n822 ,\u2_Display/n823 }),
    .b(2'b01),
    .fci(\u2_Display/lt34_c13 ),
    .fco(\u2_Display/lt34_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_16|u2_Display/lt34_15  (
    .a({\u2_Display/n820 ,\u2_Display/n821 }),
    .b(2'b11),
    .fci(\u2_Display/lt34_c15 ),
    .fco(\u2_Display/lt34_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_18|u2_Display/lt34_17  (
    .a({\u2_Display/n818 ,\u2_Display/n819 }),
    .b(2'b11),
    .fci(\u2_Display/lt34_c17 ),
    .fco(\u2_Display/lt34_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_20|u2_Display/lt34_19  (
    .a({\u2_Display/n816 ,\u2_Display/n817 }),
    .b(2'b01),
    .fci(\u2_Display/lt34_c19 ),
    .fco(\u2_Display/lt34_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_22|u2_Display/lt34_21  (
    .a({\u2_Display/n814 ,\u2_Display/n815 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c21 ),
    .fco(\u2_Display/lt34_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_24|u2_Display/lt34_23  (
    .a({\u2_Display/n812 ,\u2_Display/n813 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c23 ),
    .fco(\u2_Display/lt34_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_26|u2_Display/lt34_25  (
    .a({\u2_Display/n810 ,\u2_Display/n811 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c25 ),
    .fco(\u2_Display/lt34_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_28|u2_Display/lt34_27  (
    .a({\u2_Display/n808 ,\u2_Display/n809 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c27 ),
    .fco(\u2_Display/lt34_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_2|u2_Display/lt34_1  (
    .a({\u2_Display/n834 ,\u2_Display/n835 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c1 ),
    .fco(\u2_Display/lt34_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_30|u2_Display/lt34_29  (
    .a({\u2_Display/n806 ,\u2_Display/n807 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c29 ),
    .fco(\u2_Display/lt34_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_4|u2_Display/lt34_3  (
    .a({\u2_Display/n832 ,\u2_Display/n833 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c3 ),
    .fco(\u2_Display/lt34_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_6|u2_Display/lt34_5  (
    .a({\u2_Display/n830 ,\u2_Display/n831 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c5 ),
    .fco(\u2_Display/lt34_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_8|u2_Display/lt34_7  (
    .a({\u2_Display/n828 ,\u2_Display/n829 }),
    .b(2'b00),
    .fci(\u2_Display/lt34_c7 ),
    .fco(\u2_Display/lt34_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt34_0|u2_Display/lt34_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt34_cout|u2_Display/lt34_31  (
    .a({1'b0,\u2_Display/n805 }),
    .b(2'b10),
    .fci(\u2_Display/lt34_c31 ),
    .f({\u2_Display/n837 ,open_n52143}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_0|u2_Display/lt35_cin  (
    .a({\u2_Display/n871 ,1'b0}),
    .b({1'b0,open_n52149}),
    .fco(\u2_Display/lt35_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_10|u2_Display/lt35_9  (
    .a({\u2_Display/n861 ,\u2_Display/n862 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c9 ),
    .fco(\u2_Display/lt35_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_12|u2_Display/lt35_11  (
    .a({\u2_Display/n859 ,\u2_Display/n860 }),
    .b(2'b10),
    .fci(\u2_Display/lt35_c11 ),
    .fco(\u2_Display/lt35_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_14|u2_Display/lt35_13  (
    .a({\u2_Display/n857 ,\u2_Display/n858 }),
    .b(2'b10),
    .fci(\u2_Display/lt35_c13 ),
    .fco(\u2_Display/lt35_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_16|u2_Display/lt35_15  (
    .a({\u2_Display/n855 ,\u2_Display/n856 }),
    .b(2'b11),
    .fci(\u2_Display/lt35_c15 ),
    .fco(\u2_Display/lt35_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_18|u2_Display/lt35_17  (
    .a({\u2_Display/n853 ,\u2_Display/n854 }),
    .b(2'b11),
    .fci(\u2_Display/lt35_c17 ),
    .fco(\u2_Display/lt35_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_20|u2_Display/lt35_19  (
    .a({\u2_Display/n851 ,\u2_Display/n852 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c19 ),
    .fco(\u2_Display/lt35_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_22|u2_Display/lt35_21  (
    .a({\u2_Display/n849 ,\u2_Display/n850 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c21 ),
    .fco(\u2_Display/lt35_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_24|u2_Display/lt35_23  (
    .a({\u2_Display/n847 ,\u2_Display/n848 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c23 ),
    .fco(\u2_Display/lt35_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_26|u2_Display/lt35_25  (
    .a({\u2_Display/n845 ,\u2_Display/n846 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c25 ),
    .fco(\u2_Display/lt35_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_28|u2_Display/lt35_27  (
    .a({\u2_Display/n843 ,\u2_Display/n844 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c27 ),
    .fco(\u2_Display/lt35_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_2|u2_Display/lt35_1  (
    .a({\u2_Display/n869 ,\u2_Display/n870 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c1 ),
    .fco(\u2_Display/lt35_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_30|u2_Display/lt35_29  (
    .a({\u2_Display/n841 ,\u2_Display/n842 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c29 ),
    .fco(\u2_Display/lt35_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_4|u2_Display/lt35_3  (
    .a({\u2_Display/n867 ,\u2_Display/n868 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c3 ),
    .fco(\u2_Display/lt35_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_6|u2_Display/lt35_5  (
    .a({\u2_Display/n865 ,\u2_Display/n866 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c5 ),
    .fco(\u2_Display/lt35_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_8|u2_Display/lt35_7  (
    .a({\u2_Display/n863 ,\u2_Display/n864 }),
    .b(2'b00),
    .fci(\u2_Display/lt35_c7 ),
    .fco(\u2_Display/lt35_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt35_0|u2_Display/lt35_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt35_cout|u2_Display/lt35_31  (
    .a({1'b0,\u2_Display/n840 }),
    .b(2'b10),
    .fci(\u2_Display/lt35_c31 ),
    .f({\u2_Display/n872 ,open_n52553}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_0|u2_Display/lt36_cin  (
    .a({\u2_Display/n906 ,1'b0}),
    .b({1'b0,open_n52559}),
    .fco(\u2_Display/lt36_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_10|u2_Display/lt36_9  (
    .a({\u2_Display/n896 ,\u2_Display/n897 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c9 ),
    .fco(\u2_Display/lt36_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_12|u2_Display/lt36_11  (
    .a({\u2_Display/n894 ,\u2_Display/n895 }),
    .b(2'b01),
    .fci(\u2_Display/lt36_c11 ),
    .fco(\u2_Display/lt36_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_14|u2_Display/lt36_13  (
    .a({\u2_Display/n892 ,\u2_Display/n893 }),
    .b(2'b11),
    .fci(\u2_Display/lt36_c13 ),
    .fco(\u2_Display/lt36_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_16|u2_Display/lt36_15  (
    .a({\u2_Display/n890 ,\u2_Display/n891 }),
    .b(2'b11),
    .fci(\u2_Display/lt36_c15 ),
    .fco(\u2_Display/lt36_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_18|u2_Display/lt36_17  (
    .a({\u2_Display/n888 ,\u2_Display/n889 }),
    .b(2'b01),
    .fci(\u2_Display/lt36_c17 ),
    .fco(\u2_Display/lt36_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_20|u2_Display/lt36_19  (
    .a({\u2_Display/n886 ,\u2_Display/n887 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c19 ),
    .fco(\u2_Display/lt36_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_22|u2_Display/lt36_21  (
    .a({\u2_Display/n884 ,\u2_Display/n885 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c21 ),
    .fco(\u2_Display/lt36_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_24|u2_Display/lt36_23  (
    .a({\u2_Display/n882 ,\u2_Display/n883 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c23 ),
    .fco(\u2_Display/lt36_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_26|u2_Display/lt36_25  (
    .a({\u2_Display/n880 ,\u2_Display/n881 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c25 ),
    .fco(\u2_Display/lt36_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_28|u2_Display/lt36_27  (
    .a({\u2_Display/n878 ,\u2_Display/n879 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c27 ),
    .fco(\u2_Display/lt36_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_2|u2_Display/lt36_1  (
    .a({\u2_Display/n904 ,\u2_Display/n905 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c1 ),
    .fco(\u2_Display/lt36_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_30|u2_Display/lt36_29  (
    .a({\u2_Display/n876 ,\u2_Display/n877 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c29 ),
    .fco(\u2_Display/lt36_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_4|u2_Display/lt36_3  (
    .a({\u2_Display/n902 ,\u2_Display/n903 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c3 ),
    .fco(\u2_Display/lt36_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_6|u2_Display/lt36_5  (
    .a({\u2_Display/n900 ,\u2_Display/n901 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c5 ),
    .fco(\u2_Display/lt36_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_8|u2_Display/lt36_7  (
    .a({\u2_Display/n898 ,\u2_Display/n899 }),
    .b(2'b00),
    .fci(\u2_Display/lt36_c7 ),
    .fco(\u2_Display/lt36_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt36_0|u2_Display/lt36_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt36_cout|u2_Display/lt36_31  (
    .a({1'b0,\u2_Display/n875 }),
    .b(2'b10),
    .fci(\u2_Display/lt36_c31 ),
    .f({\u2_Display/n907 ,open_n52963}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_0|u2_Display/lt37_cin  (
    .a({\u2_Display/n941 ,1'b0}),
    .b({1'b0,open_n52969}),
    .fco(\u2_Display/lt37_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_10|u2_Display/lt37_9  (
    .a({\u2_Display/n931 ,\u2_Display/n932 }),
    .b(2'b10),
    .fci(\u2_Display/lt37_c9 ),
    .fco(\u2_Display/lt37_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_12|u2_Display/lt37_11  (
    .a({\u2_Display/n929 ,\u2_Display/n930 }),
    .b(2'b10),
    .fci(\u2_Display/lt37_c11 ),
    .fco(\u2_Display/lt37_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_14|u2_Display/lt37_13  (
    .a({\u2_Display/n927 ,\u2_Display/n928 }),
    .b(2'b11),
    .fci(\u2_Display/lt37_c13 ),
    .fco(\u2_Display/lt37_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_16|u2_Display/lt37_15  (
    .a({\u2_Display/n925 ,\u2_Display/n926 }),
    .b(2'b11),
    .fci(\u2_Display/lt37_c15 ),
    .fco(\u2_Display/lt37_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_18|u2_Display/lt37_17  (
    .a({\u2_Display/n923 ,\u2_Display/n924 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c17 ),
    .fco(\u2_Display/lt37_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_20|u2_Display/lt37_19  (
    .a({\u2_Display/n921 ,\u2_Display/n922 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c19 ),
    .fco(\u2_Display/lt37_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_22|u2_Display/lt37_21  (
    .a({\u2_Display/n919 ,\u2_Display/n920 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c21 ),
    .fco(\u2_Display/lt37_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_24|u2_Display/lt37_23  (
    .a({\u2_Display/n917 ,\u2_Display/n918 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c23 ),
    .fco(\u2_Display/lt37_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_26|u2_Display/lt37_25  (
    .a({\u2_Display/n915 ,\u2_Display/n916 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c25 ),
    .fco(\u2_Display/lt37_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_28|u2_Display/lt37_27  (
    .a({\u2_Display/n913 ,\u2_Display/n914 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c27 ),
    .fco(\u2_Display/lt37_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_2|u2_Display/lt37_1  (
    .a({\u2_Display/n939 ,\u2_Display/n940 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c1 ),
    .fco(\u2_Display/lt37_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_30|u2_Display/lt37_29  (
    .a({\u2_Display/n911 ,\u2_Display/n912 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c29 ),
    .fco(\u2_Display/lt37_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_4|u2_Display/lt37_3  (
    .a({\u2_Display/n937 ,\u2_Display/n938 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c3 ),
    .fco(\u2_Display/lt37_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_6|u2_Display/lt37_5  (
    .a({\u2_Display/n935 ,\u2_Display/n936 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c5 ),
    .fco(\u2_Display/lt37_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_8|u2_Display/lt37_7  (
    .a({\u2_Display/n933 ,\u2_Display/n934 }),
    .b(2'b00),
    .fci(\u2_Display/lt37_c7 ),
    .fco(\u2_Display/lt37_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt37_0|u2_Display/lt37_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt37_cout|u2_Display/lt37_31  (
    .a({1'b0,\u2_Display/n910 }),
    .b(2'b10),
    .fci(\u2_Display/lt37_c31 ),
    .f({\u2_Display/n942 ,open_n53373}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_0|u2_Display/lt38_cin  (
    .a({\u2_Display/n976 ,1'b0}),
    .b({1'b0,open_n53379}),
    .fco(\u2_Display/lt38_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_10|u2_Display/lt38_9  (
    .a({\u2_Display/n966 ,\u2_Display/n967 }),
    .b(2'b01),
    .fci(\u2_Display/lt38_c9 ),
    .fco(\u2_Display/lt38_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_12|u2_Display/lt38_11  (
    .a({\u2_Display/n964 ,\u2_Display/n965 }),
    .b(2'b11),
    .fci(\u2_Display/lt38_c11 ),
    .fco(\u2_Display/lt38_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_14|u2_Display/lt38_13  (
    .a({\u2_Display/n962 ,\u2_Display/n963 }),
    .b(2'b11),
    .fci(\u2_Display/lt38_c13 ),
    .fco(\u2_Display/lt38_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_16|u2_Display/lt38_15  (
    .a({\u2_Display/n960 ,\u2_Display/n961 }),
    .b(2'b01),
    .fci(\u2_Display/lt38_c15 ),
    .fco(\u2_Display/lt38_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_18|u2_Display/lt38_17  (
    .a({\u2_Display/n958 ,\u2_Display/n959 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c17 ),
    .fco(\u2_Display/lt38_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_20|u2_Display/lt38_19  (
    .a({\u2_Display/n956 ,\u2_Display/n957 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c19 ),
    .fco(\u2_Display/lt38_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_22|u2_Display/lt38_21  (
    .a({\u2_Display/n954 ,\u2_Display/n955 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c21 ),
    .fco(\u2_Display/lt38_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_24|u2_Display/lt38_23  (
    .a({\u2_Display/n952 ,\u2_Display/n953 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c23 ),
    .fco(\u2_Display/lt38_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_26|u2_Display/lt38_25  (
    .a({\u2_Display/n950 ,\u2_Display/n951 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c25 ),
    .fco(\u2_Display/lt38_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_28|u2_Display/lt38_27  (
    .a({\u2_Display/n948 ,\u2_Display/n949 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c27 ),
    .fco(\u2_Display/lt38_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_2|u2_Display/lt38_1  (
    .a({\u2_Display/n974 ,\u2_Display/n975 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c1 ),
    .fco(\u2_Display/lt38_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_30|u2_Display/lt38_29  (
    .a({\u2_Display/n946 ,\u2_Display/n947 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c29 ),
    .fco(\u2_Display/lt38_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_4|u2_Display/lt38_3  (
    .a({\u2_Display/n972 ,\u2_Display/n973 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c3 ),
    .fco(\u2_Display/lt38_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_6|u2_Display/lt38_5  (
    .a({\u2_Display/n970 ,\u2_Display/n971 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c5 ),
    .fco(\u2_Display/lt38_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_8|u2_Display/lt38_7  (
    .a({\u2_Display/n968 ,\u2_Display/n969 }),
    .b(2'b00),
    .fci(\u2_Display/lt38_c7 ),
    .fco(\u2_Display/lt38_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt38_0|u2_Display/lt38_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt38_cout|u2_Display/lt38_31  (
    .a({1'b0,\u2_Display/n945 }),
    .b(2'b10),
    .fci(\u2_Display/lt38_c31 ),
    .f({\u2_Display/n977 ,open_n53783}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_0|u2_Display/lt39_cin  (
    .a({\u2_Display/n1011 ,1'b0}),
    .b({1'b0,open_n53789}),
    .fco(\u2_Display/lt39_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_10|u2_Display/lt39_9  (
    .a({\u2_Display/n1001 ,\u2_Display/n1002 }),
    .b(2'b10),
    .fci(\u2_Display/lt39_c9 ),
    .fco(\u2_Display/lt39_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_12|u2_Display/lt39_11  (
    .a({\u2_Display/n999 ,\u2_Display/n1000 }),
    .b(2'b11),
    .fci(\u2_Display/lt39_c11 ),
    .fco(\u2_Display/lt39_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_14|u2_Display/lt39_13  (
    .a({\u2_Display/n997 ,\u2_Display/n998 }),
    .b(2'b11),
    .fci(\u2_Display/lt39_c13 ),
    .fco(\u2_Display/lt39_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_16|u2_Display/lt39_15  (
    .a({\u2_Display/n995 ,\u2_Display/n996 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c15 ),
    .fco(\u2_Display/lt39_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_18|u2_Display/lt39_17  (
    .a({\u2_Display/n993 ,\u2_Display/n994 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c17 ),
    .fco(\u2_Display/lt39_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_20|u2_Display/lt39_19  (
    .a({\u2_Display/n991 ,\u2_Display/n992 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c19 ),
    .fco(\u2_Display/lt39_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_22|u2_Display/lt39_21  (
    .a({\u2_Display/n989 ,\u2_Display/n990 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c21 ),
    .fco(\u2_Display/lt39_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_24|u2_Display/lt39_23  (
    .a({\u2_Display/n987 ,\u2_Display/n988 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c23 ),
    .fco(\u2_Display/lt39_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_26|u2_Display/lt39_25  (
    .a({\u2_Display/n985 ,\u2_Display/n986 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c25 ),
    .fco(\u2_Display/lt39_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_28|u2_Display/lt39_27  (
    .a({\u2_Display/n983 ,\u2_Display/n984 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c27 ),
    .fco(\u2_Display/lt39_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_2|u2_Display/lt39_1  (
    .a({\u2_Display/n1009 ,\u2_Display/n1010 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c1 ),
    .fco(\u2_Display/lt39_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_30|u2_Display/lt39_29  (
    .a({\u2_Display/n981 ,\u2_Display/n982 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c29 ),
    .fco(\u2_Display/lt39_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_4|u2_Display/lt39_3  (
    .a({\u2_Display/n1007 ,\u2_Display/n1008 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c3 ),
    .fco(\u2_Display/lt39_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_6|u2_Display/lt39_5  (
    .a({\u2_Display/n1005 ,\u2_Display/n1006 }),
    .b(2'b00),
    .fci(\u2_Display/lt39_c5 ),
    .fco(\u2_Display/lt39_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_8|u2_Display/lt39_7  (
    .a({\u2_Display/n1003 ,\u2_Display/n1004 }),
    .b(2'b10),
    .fci(\u2_Display/lt39_c7 ),
    .fco(\u2_Display/lt39_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt39_0|u2_Display/lt39_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt39_cout|u2_Display/lt39_31  (
    .a({1'b0,\u2_Display/n980 }),
    .b(2'b10),
    .fci(\u2_Display/lt39_c31 ),
    .f({\u2_Display/n1012 ,open_n54193}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_0|u2_Display/lt3_cin  (
    .a({\u2_Display/j [0],1'b0}),
    .b({lcd_ypos[0],open_n54199}),
    .fco(\u2_Display/lt3_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_10|u2_Display/lt3_9  (
    .a({1'b0,\u2_Display/j [9]}),
    .b(lcd_ypos[10:9]),
    .fci(\u2_Display/lt3_c9 ),
    .fco(\u2_Display/lt3_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_2|u2_Display/lt3_1  (
    .a(\u2_Display/j [2:1]),
    .b(lcd_ypos[2:1]),
    .fci(\u2_Display/lt3_c1 ),
    .fco(\u2_Display/lt3_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_4|u2_Display/lt3_3  (
    .a(\u2_Display/j [4:3]),
    .b(lcd_ypos[4:3]),
    .fci(\u2_Display/lt3_c3 ),
    .fco(\u2_Display/lt3_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_6|u2_Display/lt3_5  (
    .a(\u2_Display/j [6:5]),
    .b(lcd_ypos[6:5]),
    .fci(\u2_Display/lt3_c5 ),
    .fco(\u2_Display/lt3_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_8|u2_Display/lt3_7  (
    .a(\u2_Display/j [8:7]),
    .b(lcd_ypos[8:7]),
    .fci(\u2_Display/lt3_c7 ),
    .fco(\u2_Display/lt3_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt3_0|u2_Display/lt3_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt3_cout|u2_Display/lt3_11  (
    .a(2'b00),
    .b({1'b1,lcd_ypos[11]}),
    .fci(\u2_Display/lt3_c11 ),
    .f({\u2_Display/n50 ,open_n54363}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_0|u2_Display/lt40_cin  (
    .a({\u2_Display/n1046 ,1'b0}),
    .b({1'b0,open_n54369}),
    .fco(\u2_Display/lt40_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_10|u2_Display/lt40_9  (
    .a({\u2_Display/n1036 ,\u2_Display/n1037 }),
    .b(2'b11),
    .fci(\u2_Display/lt40_c9 ),
    .fco(\u2_Display/lt40_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_12|u2_Display/lt40_11  (
    .a({\u2_Display/n1034 ,\u2_Display/n1035 }),
    .b(2'b11),
    .fci(\u2_Display/lt40_c11 ),
    .fco(\u2_Display/lt40_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_14|u2_Display/lt40_13  (
    .a({\u2_Display/n1032 ,\u2_Display/n1033 }),
    .b(2'b01),
    .fci(\u2_Display/lt40_c13 ),
    .fco(\u2_Display/lt40_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_16|u2_Display/lt40_15  (
    .a({\u2_Display/n1030 ,\u2_Display/n1031 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c15 ),
    .fco(\u2_Display/lt40_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_18|u2_Display/lt40_17  (
    .a({\u2_Display/n1028 ,\u2_Display/n1029 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c17 ),
    .fco(\u2_Display/lt40_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_20|u2_Display/lt40_19  (
    .a({\u2_Display/n1026 ,\u2_Display/n1027 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c19 ),
    .fco(\u2_Display/lt40_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_22|u2_Display/lt40_21  (
    .a({\u2_Display/n1024 ,\u2_Display/n1025 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c21 ),
    .fco(\u2_Display/lt40_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_24|u2_Display/lt40_23  (
    .a({\u2_Display/n1022 ,\u2_Display/n1023 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c23 ),
    .fco(\u2_Display/lt40_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_26|u2_Display/lt40_25  (
    .a({\u2_Display/n1020 ,\u2_Display/n1021 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c25 ),
    .fco(\u2_Display/lt40_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_28|u2_Display/lt40_27  (
    .a({\u2_Display/n1018 ,\u2_Display/n1019 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c27 ),
    .fco(\u2_Display/lt40_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_2|u2_Display/lt40_1  (
    .a({\u2_Display/n1044 ,\u2_Display/n1045 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c1 ),
    .fco(\u2_Display/lt40_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_30|u2_Display/lt40_29  (
    .a({\u2_Display/n1016 ,\u2_Display/n1017 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c29 ),
    .fco(\u2_Display/lt40_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_4|u2_Display/lt40_3  (
    .a({\u2_Display/n1042 ,\u2_Display/n1043 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c3 ),
    .fco(\u2_Display/lt40_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_6|u2_Display/lt40_5  (
    .a({\u2_Display/n1040 ,\u2_Display/n1041 }),
    .b(2'b00),
    .fci(\u2_Display/lt40_c5 ),
    .fco(\u2_Display/lt40_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_8|u2_Display/lt40_7  (
    .a({\u2_Display/n1038 ,\u2_Display/n1039 }),
    .b(2'b01),
    .fci(\u2_Display/lt40_c7 ),
    .fco(\u2_Display/lt40_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt40_0|u2_Display/lt40_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt40_cout|u2_Display/lt40_31  (
    .a({1'b0,\u2_Display/n1015 }),
    .b(2'b10),
    .fci(\u2_Display/lt40_c31 ),
    .f({\u2_Display/n1047 ,open_n54773}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_0|u2_Display/lt41_cin  (
    .a({\u2_Display/n1081 ,1'b0}),
    .b({1'b0,open_n54779}),
    .fco(\u2_Display/lt41_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_10|u2_Display/lt41_9  (
    .a({\u2_Display/n1071 ,\u2_Display/n1072 }),
    .b(2'b11),
    .fci(\u2_Display/lt41_c9 ),
    .fco(\u2_Display/lt41_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_12|u2_Display/lt41_11  (
    .a({\u2_Display/n1069 ,\u2_Display/n1070 }),
    .b(2'b11),
    .fci(\u2_Display/lt41_c11 ),
    .fco(\u2_Display/lt41_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_14|u2_Display/lt41_13  (
    .a({\u2_Display/n1067 ,\u2_Display/n1068 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c13 ),
    .fco(\u2_Display/lt41_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_16|u2_Display/lt41_15  (
    .a({\u2_Display/n1065 ,\u2_Display/n1066 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c15 ),
    .fco(\u2_Display/lt41_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_18|u2_Display/lt41_17  (
    .a({\u2_Display/n1063 ,\u2_Display/n1064 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c17 ),
    .fco(\u2_Display/lt41_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_20|u2_Display/lt41_19  (
    .a({\u2_Display/n1061 ,\u2_Display/n1062 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c19 ),
    .fco(\u2_Display/lt41_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_22|u2_Display/lt41_21  (
    .a({\u2_Display/n1059 ,\u2_Display/n1060 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c21 ),
    .fco(\u2_Display/lt41_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_24|u2_Display/lt41_23  (
    .a({\u2_Display/n1057 ,\u2_Display/n1058 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c23 ),
    .fco(\u2_Display/lt41_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_26|u2_Display/lt41_25  (
    .a({\u2_Display/n1055 ,\u2_Display/n1056 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c25 ),
    .fco(\u2_Display/lt41_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_28|u2_Display/lt41_27  (
    .a({\u2_Display/n1053 ,\u2_Display/n1054 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c27 ),
    .fco(\u2_Display/lt41_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_2|u2_Display/lt41_1  (
    .a({\u2_Display/n1079 ,\u2_Display/n1080 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c1 ),
    .fco(\u2_Display/lt41_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_30|u2_Display/lt41_29  (
    .a({\u2_Display/n1051 ,\u2_Display/n1052 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c29 ),
    .fco(\u2_Display/lt41_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_4|u2_Display/lt41_3  (
    .a({\u2_Display/n1077 ,\u2_Display/n1078 }),
    .b(2'b00),
    .fci(\u2_Display/lt41_c3 ),
    .fco(\u2_Display/lt41_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_6|u2_Display/lt41_5  (
    .a({\u2_Display/n1075 ,\u2_Display/n1076 }),
    .b(2'b10),
    .fci(\u2_Display/lt41_c5 ),
    .fco(\u2_Display/lt41_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_8|u2_Display/lt41_7  (
    .a({\u2_Display/n1073 ,\u2_Display/n1074 }),
    .b(2'b10),
    .fci(\u2_Display/lt41_c7 ),
    .fco(\u2_Display/lt41_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt41_0|u2_Display/lt41_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt41_cout|u2_Display/lt41_31  (
    .a({1'b0,\u2_Display/n1050 }),
    .b(2'b10),
    .fci(\u2_Display/lt41_c31 ),
    .f({\u2_Display/n1082 ,open_n55183}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_0|u2_Display/lt42_cin  (
    .a({\u2_Display/n1116 ,1'b0}),
    .b({1'b0,open_n55189}),
    .fco(\u2_Display/lt42_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_10|u2_Display/lt42_9  (
    .a({\u2_Display/n1106 ,\u2_Display/n1107 }),
    .b(2'b11),
    .fci(\u2_Display/lt42_c9 ),
    .fco(\u2_Display/lt42_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_12|u2_Display/lt42_11  (
    .a({\u2_Display/n1104 ,\u2_Display/n1105 }),
    .b(2'b01),
    .fci(\u2_Display/lt42_c11 ),
    .fco(\u2_Display/lt42_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_14|u2_Display/lt42_13  (
    .a({\u2_Display/n1102 ,\u2_Display/n1103 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c13 ),
    .fco(\u2_Display/lt42_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_16|u2_Display/lt42_15  (
    .a({\u2_Display/n1100 ,\u2_Display/n1101 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c15 ),
    .fco(\u2_Display/lt42_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_18|u2_Display/lt42_17  (
    .a({\u2_Display/n1098 ,\u2_Display/n1099 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c17 ),
    .fco(\u2_Display/lt42_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_20|u2_Display/lt42_19  (
    .a({\u2_Display/n1096 ,\u2_Display/n1097 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c19 ),
    .fco(\u2_Display/lt42_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_22|u2_Display/lt42_21  (
    .a({\u2_Display/n1094 ,\u2_Display/n1095 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c21 ),
    .fco(\u2_Display/lt42_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_24|u2_Display/lt42_23  (
    .a({\u2_Display/n1092 ,\u2_Display/n1093 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c23 ),
    .fco(\u2_Display/lt42_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_26|u2_Display/lt42_25  (
    .a({\u2_Display/n1090 ,\u2_Display/n1091 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c25 ),
    .fco(\u2_Display/lt42_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_28|u2_Display/lt42_27  (
    .a({\u2_Display/n1088 ,\u2_Display/n1089 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c27 ),
    .fco(\u2_Display/lt42_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_2|u2_Display/lt42_1  (
    .a({\u2_Display/n1114 ,\u2_Display/n1115 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c1 ),
    .fco(\u2_Display/lt42_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_30|u2_Display/lt42_29  (
    .a({\u2_Display/n1086 ,\u2_Display/n1087 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c29 ),
    .fco(\u2_Display/lt42_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_4|u2_Display/lt42_3  (
    .a({\u2_Display/n1112 ,\u2_Display/n1113 }),
    .b(2'b00),
    .fci(\u2_Display/lt42_c3 ),
    .fco(\u2_Display/lt42_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_6|u2_Display/lt42_5  (
    .a({\u2_Display/n1110 ,\u2_Display/n1111 }),
    .b(2'b01),
    .fci(\u2_Display/lt42_c5 ),
    .fco(\u2_Display/lt42_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_8|u2_Display/lt42_7  (
    .a({\u2_Display/n1108 ,\u2_Display/n1109 }),
    .b(2'b11),
    .fci(\u2_Display/lt42_c7 ),
    .fco(\u2_Display/lt42_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt42_0|u2_Display/lt42_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt42_cout|u2_Display/lt42_31  (
    .a({1'b0,\u2_Display/n1085 }),
    .b(2'b10),
    .fci(\u2_Display/lt42_c31 ),
    .f({\u2_Display/n1117 ,open_n55593}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_0|u2_Display/lt43_cin  (
    .a({\u2_Display/n1151 ,1'b0}),
    .b({1'b0,open_n55599}),
    .fco(\u2_Display/lt43_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_10|u2_Display/lt43_9  (
    .a({\u2_Display/n1141 ,\u2_Display/n1142 }),
    .b(2'b11),
    .fci(\u2_Display/lt43_c9 ),
    .fco(\u2_Display/lt43_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_12|u2_Display/lt43_11  (
    .a({\u2_Display/n1139 ,\u2_Display/n1140 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c11 ),
    .fco(\u2_Display/lt43_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_14|u2_Display/lt43_13  (
    .a({\u2_Display/n1137 ,\u2_Display/n1138 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c13 ),
    .fco(\u2_Display/lt43_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_16|u2_Display/lt43_15  (
    .a({\u2_Display/n1135 ,\u2_Display/n1136 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c15 ),
    .fco(\u2_Display/lt43_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_18|u2_Display/lt43_17  (
    .a({\u2_Display/n1133 ,\u2_Display/n1134 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c17 ),
    .fco(\u2_Display/lt43_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_20|u2_Display/lt43_19  (
    .a({\u2_Display/n1131 ,\u2_Display/n1132 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c19 ),
    .fco(\u2_Display/lt43_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_22|u2_Display/lt43_21  (
    .a({\u2_Display/n1129 ,\u2_Display/n1130 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c21 ),
    .fco(\u2_Display/lt43_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_24|u2_Display/lt43_23  (
    .a({\u2_Display/n1127 ,\u2_Display/n1128 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c23 ),
    .fco(\u2_Display/lt43_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_26|u2_Display/lt43_25  (
    .a({\u2_Display/n1125 ,\u2_Display/n1126 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c25 ),
    .fco(\u2_Display/lt43_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_28|u2_Display/lt43_27  (
    .a({\u2_Display/n1123 ,\u2_Display/n1124 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c27 ),
    .fco(\u2_Display/lt43_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_2|u2_Display/lt43_1  (
    .a({\u2_Display/n1149 ,\u2_Display/n1150 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c1 ),
    .fco(\u2_Display/lt43_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_30|u2_Display/lt43_29  (
    .a({\u2_Display/n1121 ,\u2_Display/n1122 }),
    .b(2'b00),
    .fci(\u2_Display/lt43_c29 ),
    .fco(\u2_Display/lt43_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_4|u2_Display/lt43_3  (
    .a({\u2_Display/n1147 ,\u2_Display/n1148 }),
    .b(2'b10),
    .fci(\u2_Display/lt43_c3 ),
    .fco(\u2_Display/lt43_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_6|u2_Display/lt43_5  (
    .a({\u2_Display/n1145 ,\u2_Display/n1146 }),
    .b(2'b10),
    .fci(\u2_Display/lt43_c5 ),
    .fco(\u2_Display/lt43_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_8|u2_Display/lt43_7  (
    .a({\u2_Display/n1143 ,\u2_Display/n1144 }),
    .b(2'b11),
    .fci(\u2_Display/lt43_c7 ),
    .fco(\u2_Display/lt43_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt43_0|u2_Display/lt43_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt43_cout|u2_Display/lt43_31  (
    .a({1'b0,\u2_Display/n1120 }),
    .b(2'b10),
    .fci(\u2_Display/lt43_c31 ),
    .f({\u2_Display/n1152 ,open_n56003}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_0|u2_Display/lt44_cin  (
    .a({\u2_Display/n1186 ,1'b0}),
    .b({1'b0,open_n56009}),
    .fco(\u2_Display/lt44_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_10|u2_Display/lt44_9  (
    .a({\u2_Display/n1176 ,\u2_Display/n1177 }),
    .b(2'b01),
    .fci(\u2_Display/lt44_c9 ),
    .fco(\u2_Display/lt44_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_12|u2_Display/lt44_11  (
    .a({\u2_Display/n1174 ,\u2_Display/n1175 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c11 ),
    .fco(\u2_Display/lt44_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_14|u2_Display/lt44_13  (
    .a({\u2_Display/n1172 ,\u2_Display/n1173 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c13 ),
    .fco(\u2_Display/lt44_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_16|u2_Display/lt44_15  (
    .a({\u2_Display/n1170 ,\u2_Display/n1171 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c15 ),
    .fco(\u2_Display/lt44_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_18|u2_Display/lt44_17  (
    .a({\u2_Display/n1168 ,\u2_Display/n1169 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c17 ),
    .fco(\u2_Display/lt44_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_20|u2_Display/lt44_19  (
    .a({\u2_Display/n1166 ,\u2_Display/n1167 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c19 ),
    .fco(\u2_Display/lt44_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_22|u2_Display/lt44_21  (
    .a({\u2_Display/n1164 ,\u2_Display/n1165 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c21 ),
    .fco(\u2_Display/lt44_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_24|u2_Display/lt44_23  (
    .a({\u2_Display/n1162 ,\u2_Display/n1163 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c23 ),
    .fco(\u2_Display/lt44_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_26|u2_Display/lt44_25  (
    .a({\u2_Display/n1160 ,\u2_Display/n1161 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c25 ),
    .fco(\u2_Display/lt44_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_28|u2_Display/lt44_27  (
    .a({\u2_Display/n1158 ,\u2_Display/n1159 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c27 ),
    .fco(\u2_Display/lt44_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_2|u2_Display/lt44_1  (
    .a({\u2_Display/n1184 ,\u2_Display/n1185 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c1 ),
    .fco(\u2_Display/lt44_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_30|u2_Display/lt44_29  (
    .a({\u2_Display/n1156 ,\u2_Display/n1157 }),
    .b(2'b00),
    .fci(\u2_Display/lt44_c29 ),
    .fco(\u2_Display/lt44_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_4|u2_Display/lt44_3  (
    .a({\u2_Display/n1182 ,\u2_Display/n1183 }),
    .b(2'b01),
    .fci(\u2_Display/lt44_c3 ),
    .fco(\u2_Display/lt44_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_6|u2_Display/lt44_5  (
    .a({\u2_Display/n1180 ,\u2_Display/n1181 }),
    .b(2'b11),
    .fci(\u2_Display/lt44_c5 ),
    .fco(\u2_Display/lt44_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_8|u2_Display/lt44_7  (
    .a({\u2_Display/n1178 ,\u2_Display/n1179 }),
    .b(2'b11),
    .fci(\u2_Display/lt44_c7 ),
    .fco(\u2_Display/lt44_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt44_0|u2_Display/lt44_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt44_cout|u2_Display/lt44_31  (
    .a({1'b0,\u2_Display/n1155 }),
    .b(2'b10),
    .fci(\u2_Display/lt44_c31 ),
    .f({\u2_Display/n1187 ,open_n56413}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_0|u2_Display/lt4_2_cin  (
    .a({lcd_xpos[0],1'b0}),
    .b({\u2_Display/i [0],open_n56419}),
    .fco(\u2_Display/lt4_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_10|u2_Display/lt4_2_9  (
    .a(lcd_xpos[10:9]),
    .b(\u2_Display/n94 [3:2]),
    .fci(\u2_Display/lt4_2_c9 ),
    .fco(\u2_Display/lt4_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_2|u2_Display/lt4_2_1  (
    .a(lcd_xpos[2:1]),
    .b(\u2_Display/i [2:1]),
    .fci(\u2_Display/lt4_2_c1 ),
    .fco(\u2_Display/lt4_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_4|u2_Display/lt4_2_3  (
    .a(lcd_xpos[4:3]),
    .b(\u2_Display/i [4:3]),
    .fci(\u2_Display/lt4_2_c3 ),
    .fco(\u2_Display/lt4_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_6|u2_Display/lt4_2_5  (
    .a(lcd_xpos[6:5]),
    .b(\u2_Display/i [6:5]),
    .fci(\u2_Display/lt4_2_c5 ),
    .fco(\u2_Display/lt4_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_8|u2_Display/lt4_2_7  (
    .a(lcd_xpos[8:7]),
    .b(\u2_Display/n94 [1:0]),
    .fci(\u2_Display/lt4_2_c7 ),
    .fco(\u2_Display/lt4_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt4_2_0|u2_Display/lt4_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt4_2_cout|u2_Display/lt4_2_11  (
    .a({1'b0,lcd_xpos[11]}),
    .b({1'b1,\u2_Display/add4_2_co }),
    .fci(\u2_Display/lt4_2_c11 ),
    .f({\u2_Display/n95 ,open_n56583}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_0|u2_Display/lt55_cin  (
    .a({\u2_Display/counta [0],1'b0}),
    .b({1'b0,open_n56589}),
    .fco(\u2_Display/lt55_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_10|u2_Display/lt55_9  (
    .a(\u2_Display/counta [10:9]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c9 ),
    .fco(\u2_Display/lt55_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_12|u2_Display/lt55_11  (
    .a(\u2_Display/counta [12:11]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c11 ),
    .fco(\u2_Display/lt55_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_14|u2_Display/lt55_13  (
    .a(\u2_Display/counta [14:13]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c13 ),
    .fco(\u2_Display/lt55_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_16|u2_Display/lt55_15  (
    .a(\u2_Display/counta [16:15]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c15 ),
    .fco(\u2_Display/lt55_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_18|u2_Display/lt55_17  (
    .a(\u2_Display/counta [18:17]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c17 ),
    .fco(\u2_Display/lt55_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_20|u2_Display/lt55_19  (
    .a(\u2_Display/counta [20:19]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c19 ),
    .fco(\u2_Display/lt55_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_22|u2_Display/lt55_21  (
    .a(\u2_Display/counta [22:21]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c21 ),
    .fco(\u2_Display/lt55_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_24|u2_Display/lt55_23  (
    .a(\u2_Display/counta [24:23]),
    .b(2'b10),
    .fci(\u2_Display/lt55_c23 ),
    .fco(\u2_Display/lt55_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_26|u2_Display/lt55_25  (
    .a(\u2_Display/counta [26:25]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c25 ),
    .fco(\u2_Display/lt55_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_28|u2_Display/lt55_27  (
    .a(\u2_Display/counta [28:27]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c27 ),
    .fco(\u2_Display/lt55_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_2|u2_Display/lt55_1  (
    .a(\u2_Display/counta [2:1]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c1 ),
    .fco(\u2_Display/lt55_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_30|u2_Display/lt55_29  (
    .a(\u2_Display/counta [30:29]),
    .b(2'b11),
    .fci(\u2_Display/lt55_c29 ),
    .fco(\u2_Display/lt55_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_4|u2_Display/lt55_3  (
    .a(\u2_Display/counta [4:3]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c3 ),
    .fco(\u2_Display/lt55_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_6|u2_Display/lt55_5  (
    .a(\u2_Display/counta [6:5]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c5 ),
    .fco(\u2_Display/lt55_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_8|u2_Display/lt55_7  (
    .a(\u2_Display/counta [8:7]),
    .b(2'b00),
    .fci(\u2_Display/lt55_c7 ),
    .fco(\u2_Display/lt55_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt55_0|u2_Display/lt55_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt55_cout|u2_Display/lt55_31  (
    .a({1'b0,\u2_Display/counta [31]}),
    .b(2'b11),
    .fci(\u2_Display/lt55_c31 ),
    .f({\u2_Display/n1540 ,open_n56993}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_0|u2_Display/lt56_cin  (
    .a({\u2_Display/n1574 ,1'b0}),
    .b({1'b0,open_n56999}),
    .fco(\u2_Display/lt56_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_10|u2_Display/lt56_9  (
    .a({\u2_Display/n1564 ,\u2_Display/n1565 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c9 ),
    .fco(\u2_Display/lt56_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_12|u2_Display/lt56_11  (
    .a({\u2_Display/n1562 ,\u2_Display/n1563 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c11 ),
    .fco(\u2_Display/lt56_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_14|u2_Display/lt56_13  (
    .a({\u2_Display/n1560 ,\u2_Display/n1561 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c13 ),
    .fco(\u2_Display/lt56_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_16|u2_Display/lt56_15  (
    .a({\u2_Display/n1558 ,\u2_Display/n1559 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c15 ),
    .fco(\u2_Display/lt56_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_18|u2_Display/lt56_17  (
    .a({\u2_Display/n1556 ,\u2_Display/n1557 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c17 ),
    .fco(\u2_Display/lt56_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_20|u2_Display/lt56_19  (
    .a({\u2_Display/n1554 ,\u2_Display/n1555 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c19 ),
    .fco(\u2_Display/lt56_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_22|u2_Display/lt56_21  (
    .a({\u2_Display/n1552 ,\u2_Display/n1553 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c21 ),
    .fco(\u2_Display/lt56_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_24|u2_Display/lt56_23  (
    .a({\u2_Display/n1550 ,\u2_Display/n1551 }),
    .b(2'b01),
    .fci(\u2_Display/lt56_c23 ),
    .fco(\u2_Display/lt56_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_26|u2_Display/lt56_25  (
    .a({\u2_Display/n1548 ,\u2_Display/n1549 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c25 ),
    .fco(\u2_Display/lt56_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_28|u2_Display/lt56_27  (
    .a({\u2_Display/n1546 ,\u2_Display/n1547 }),
    .b(2'b10),
    .fci(\u2_Display/lt56_c27 ),
    .fco(\u2_Display/lt56_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_2|u2_Display/lt56_1  (
    .a({\u2_Display/n1572 ,\u2_Display/n1573 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c1 ),
    .fco(\u2_Display/lt56_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_30|u2_Display/lt56_29  (
    .a({\u2_Display/n1544 ,\u2_Display/n1545 }),
    .b(2'b11),
    .fci(\u2_Display/lt56_c29 ),
    .fco(\u2_Display/lt56_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_4|u2_Display/lt56_3  (
    .a({\u2_Display/n1570 ,\u2_Display/n1571 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c3 ),
    .fco(\u2_Display/lt56_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_6|u2_Display/lt56_5  (
    .a({\u2_Display/n1568 ,\u2_Display/n1569 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c5 ),
    .fco(\u2_Display/lt56_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_8|u2_Display/lt56_7  (
    .a({\u2_Display/n1566 ,\u2_Display/n1567 }),
    .b(2'b00),
    .fci(\u2_Display/lt56_c7 ),
    .fco(\u2_Display/lt56_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt56_0|u2_Display/lt56_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt56_cout|u2_Display/lt56_31  (
    .a({1'b0,\u2_Display/n1543 }),
    .b(2'b10),
    .fci(\u2_Display/lt56_c31 ),
    .f({\u2_Display/n1575 ,open_n57403}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_0|u2_Display/lt57_cin  (
    .a({\u2_Display/n1609 ,1'b0}),
    .b({1'b0,open_n57409}),
    .fco(\u2_Display/lt57_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_10|u2_Display/lt57_9  (
    .a({\u2_Display/n1599 ,\u2_Display/n1600 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c9 ),
    .fco(\u2_Display/lt57_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_12|u2_Display/lt57_11  (
    .a({\u2_Display/n1597 ,\u2_Display/n1598 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c11 ),
    .fco(\u2_Display/lt57_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_14|u2_Display/lt57_13  (
    .a({\u2_Display/n1595 ,\u2_Display/n1596 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c13 ),
    .fco(\u2_Display/lt57_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_16|u2_Display/lt57_15  (
    .a({\u2_Display/n1593 ,\u2_Display/n1594 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c15 ),
    .fco(\u2_Display/lt57_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_18|u2_Display/lt57_17  (
    .a({\u2_Display/n1591 ,\u2_Display/n1592 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c17 ),
    .fco(\u2_Display/lt57_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_20|u2_Display/lt57_19  (
    .a({\u2_Display/n1589 ,\u2_Display/n1590 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c19 ),
    .fco(\u2_Display/lt57_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_22|u2_Display/lt57_21  (
    .a({\u2_Display/n1587 ,\u2_Display/n1588 }),
    .b(2'b10),
    .fci(\u2_Display/lt57_c21 ),
    .fco(\u2_Display/lt57_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_24|u2_Display/lt57_23  (
    .a({\u2_Display/n1585 ,\u2_Display/n1586 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c23 ),
    .fco(\u2_Display/lt57_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_26|u2_Display/lt57_25  (
    .a({\u2_Display/n1583 ,\u2_Display/n1584 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c25 ),
    .fco(\u2_Display/lt57_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_28|u2_Display/lt57_27  (
    .a({\u2_Display/n1581 ,\u2_Display/n1582 }),
    .b(2'b11),
    .fci(\u2_Display/lt57_c27 ),
    .fco(\u2_Display/lt57_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_2|u2_Display/lt57_1  (
    .a({\u2_Display/n1607 ,\u2_Display/n1608 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c1 ),
    .fco(\u2_Display/lt57_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_30|u2_Display/lt57_29  (
    .a({\u2_Display/n1579 ,\u2_Display/n1580 }),
    .b(2'b01),
    .fci(\u2_Display/lt57_c29 ),
    .fco(\u2_Display/lt57_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_4|u2_Display/lt57_3  (
    .a({\u2_Display/n1605 ,\u2_Display/n1606 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c3 ),
    .fco(\u2_Display/lt57_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_6|u2_Display/lt57_5  (
    .a({\u2_Display/n1603 ,\u2_Display/n1604 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c5 ),
    .fco(\u2_Display/lt57_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_8|u2_Display/lt57_7  (
    .a({\u2_Display/n1601 ,\u2_Display/n1602 }),
    .b(2'b00),
    .fci(\u2_Display/lt57_c7 ),
    .fco(\u2_Display/lt57_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt57_0|u2_Display/lt57_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt57_cout|u2_Display/lt57_31  (
    .a({1'b0,\u2_Display/n1578 }),
    .b(2'b10),
    .fci(\u2_Display/lt57_c31 ),
    .f({\u2_Display/n1610 ,open_n57813}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_0|u2_Display/lt58_cin  (
    .a({\u2_Display/n1644 ,1'b0}),
    .b({1'b0,open_n57819}),
    .fco(\u2_Display/lt58_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_10|u2_Display/lt58_9  (
    .a({\u2_Display/n1634 ,\u2_Display/n1635 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c9 ),
    .fco(\u2_Display/lt58_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_12|u2_Display/lt58_11  (
    .a({\u2_Display/n1632 ,\u2_Display/n1633 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c11 ),
    .fco(\u2_Display/lt58_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_14|u2_Display/lt58_13  (
    .a({\u2_Display/n1630 ,\u2_Display/n1631 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c13 ),
    .fco(\u2_Display/lt58_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_16|u2_Display/lt58_15  (
    .a({\u2_Display/n1628 ,\u2_Display/n1629 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c15 ),
    .fco(\u2_Display/lt58_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_18|u2_Display/lt58_17  (
    .a({\u2_Display/n1626 ,\u2_Display/n1627 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c17 ),
    .fco(\u2_Display/lt58_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_20|u2_Display/lt58_19  (
    .a({\u2_Display/n1624 ,\u2_Display/n1625 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c19 ),
    .fco(\u2_Display/lt58_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_22|u2_Display/lt58_21  (
    .a({\u2_Display/n1622 ,\u2_Display/n1623 }),
    .b(2'b01),
    .fci(\u2_Display/lt58_c21 ),
    .fco(\u2_Display/lt58_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_24|u2_Display/lt58_23  (
    .a({\u2_Display/n1620 ,\u2_Display/n1621 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c23 ),
    .fco(\u2_Display/lt58_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_26|u2_Display/lt58_25  (
    .a({\u2_Display/n1618 ,\u2_Display/n1619 }),
    .b(2'b10),
    .fci(\u2_Display/lt58_c25 ),
    .fco(\u2_Display/lt58_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_28|u2_Display/lt58_27  (
    .a({\u2_Display/n1616 ,\u2_Display/n1617 }),
    .b(2'b11),
    .fci(\u2_Display/lt58_c27 ),
    .fco(\u2_Display/lt58_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_2|u2_Display/lt58_1  (
    .a({\u2_Display/n1642 ,\u2_Display/n1643 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c1 ),
    .fco(\u2_Display/lt58_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_30|u2_Display/lt58_29  (
    .a({\u2_Display/n1614 ,\u2_Display/n1615 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c29 ),
    .fco(\u2_Display/lt58_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_4|u2_Display/lt58_3  (
    .a({\u2_Display/n1640 ,\u2_Display/n1641 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c3 ),
    .fco(\u2_Display/lt58_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_6|u2_Display/lt58_5  (
    .a({\u2_Display/n1638 ,\u2_Display/n1639 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c5 ),
    .fco(\u2_Display/lt58_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_8|u2_Display/lt58_7  (
    .a({\u2_Display/n1636 ,\u2_Display/n1637 }),
    .b(2'b00),
    .fci(\u2_Display/lt58_c7 ),
    .fco(\u2_Display/lt58_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt58_0|u2_Display/lt58_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt58_cout|u2_Display/lt58_31  (
    .a({1'b0,\u2_Display/n1613 }),
    .b(2'b10),
    .fci(\u2_Display/lt58_c31 ),
    .f({\u2_Display/n1645 ,open_n58223}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_0|u2_Display/lt59_cin  (
    .a({\u2_Display/n1679 ,1'b0}),
    .b({1'b0,open_n58229}),
    .fco(\u2_Display/lt59_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_10|u2_Display/lt59_9  (
    .a({\u2_Display/n1669 ,\u2_Display/n1670 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c9 ),
    .fco(\u2_Display/lt59_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_12|u2_Display/lt59_11  (
    .a({\u2_Display/n1667 ,\u2_Display/n1668 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c11 ),
    .fco(\u2_Display/lt59_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_14|u2_Display/lt59_13  (
    .a({\u2_Display/n1665 ,\u2_Display/n1666 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c13 ),
    .fco(\u2_Display/lt59_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_16|u2_Display/lt59_15  (
    .a({\u2_Display/n1663 ,\u2_Display/n1664 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c15 ),
    .fco(\u2_Display/lt59_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_18|u2_Display/lt59_17  (
    .a({\u2_Display/n1661 ,\u2_Display/n1662 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c17 ),
    .fco(\u2_Display/lt59_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_20|u2_Display/lt59_19  (
    .a({\u2_Display/n1659 ,\u2_Display/n1660 }),
    .b(2'b10),
    .fci(\u2_Display/lt59_c19 ),
    .fco(\u2_Display/lt59_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_22|u2_Display/lt59_21  (
    .a({\u2_Display/n1657 ,\u2_Display/n1658 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c21 ),
    .fco(\u2_Display/lt59_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_24|u2_Display/lt59_23  (
    .a({\u2_Display/n1655 ,\u2_Display/n1656 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c23 ),
    .fco(\u2_Display/lt59_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_26|u2_Display/lt59_25  (
    .a({\u2_Display/n1653 ,\u2_Display/n1654 }),
    .b(2'b11),
    .fci(\u2_Display/lt59_c25 ),
    .fco(\u2_Display/lt59_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_28|u2_Display/lt59_27  (
    .a({\u2_Display/n1651 ,\u2_Display/n1652 }),
    .b(2'b01),
    .fci(\u2_Display/lt59_c27 ),
    .fco(\u2_Display/lt59_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_2|u2_Display/lt59_1  (
    .a({\u2_Display/n1677 ,\u2_Display/n1678 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c1 ),
    .fco(\u2_Display/lt59_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_30|u2_Display/lt59_29  (
    .a({\u2_Display/n1649 ,\u2_Display/n1650 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c29 ),
    .fco(\u2_Display/lt59_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_4|u2_Display/lt59_3  (
    .a({\u2_Display/n1675 ,\u2_Display/n1676 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c3 ),
    .fco(\u2_Display/lt59_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_6|u2_Display/lt59_5  (
    .a({\u2_Display/n1673 ,\u2_Display/n1674 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c5 ),
    .fco(\u2_Display/lt59_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_8|u2_Display/lt59_7  (
    .a({\u2_Display/n1671 ,\u2_Display/n1672 }),
    .b(2'b00),
    .fci(\u2_Display/lt59_c7 ),
    .fco(\u2_Display/lt59_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt59_0|u2_Display/lt59_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt59_cout|u2_Display/lt59_31  (
    .a({1'b0,\u2_Display/n1648 }),
    .b(2'b10),
    .fci(\u2_Display/lt59_c31 ),
    .f({\u2_Display/n1680 ,open_n58633}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_0|u2_Display/lt5_2_cin  (
    .a({\u2_Display/n96 [0],1'b0}),
    .b({lcd_xpos[0],open_n58639}),
    .fco(\u2_Display/lt5_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_10|u2_Display/lt5_2_9  (
    .a(\u2_Display/n96 [10:9]),
    .b(lcd_xpos[10:9]),
    .fci(\u2_Display/lt5_2_c9 ),
    .fco(\u2_Display/lt5_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_12|u2_Display/lt5_2_11  (
    .a({\u2_Display/n96 [31],\u2_Display/n96 [31]}),
    .b({1'b0,lcd_xpos[11]}),
    .fci(\u2_Display/lt5_2_c11 ),
    .fco(\u2_Display/lt5_2_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_2|u2_Display/lt5_2_1  (
    .a(\u2_Display/n96 [2:1]),
    .b(lcd_xpos[2:1]),
    .fci(\u2_Display/lt5_2_c1 ),
    .fco(\u2_Display/lt5_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_4|u2_Display/lt5_2_3  (
    .a(\u2_Display/n96 [4:3]),
    .b(lcd_xpos[4:3]),
    .fci(\u2_Display/lt5_2_c3 ),
    .fco(\u2_Display/lt5_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_6|u2_Display/lt5_2_5  (
    .a(\u2_Display/n96 [6:5]),
    .b(lcd_xpos[6:5]),
    .fci(\u2_Display/lt5_2_c5 ),
    .fco(\u2_Display/lt5_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_8|u2_Display/lt5_2_7  (
    .a(\u2_Display/n96 [8:7]),
    .b(lcd_xpos[8:7]),
    .fci(\u2_Display/lt5_2_c7 ),
    .fco(\u2_Display/lt5_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt5_2_0|u2_Display/lt5_2_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt5_2_cout_al_u5061  (
    .a({open_n58809,1'b0}),
    .b({open_n58810,1'b1}),
    .fci(\u2_Display/lt5_2_c13 ),
    .f({open_n58829,\u2_Display/n97 }));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_0|u2_Display/lt60_cin  (
    .a({\u2_Display/n1714 ,1'b0}),
    .b({1'b0,open_n58835}),
    .fco(\u2_Display/lt60_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_10|u2_Display/lt60_9  (
    .a({\u2_Display/n1704 ,\u2_Display/n1705 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c9 ),
    .fco(\u2_Display/lt60_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_12|u2_Display/lt60_11  (
    .a({\u2_Display/n1702 ,\u2_Display/n1703 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c11 ),
    .fco(\u2_Display/lt60_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_14|u2_Display/lt60_13  (
    .a({\u2_Display/n1700 ,\u2_Display/n1701 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c13 ),
    .fco(\u2_Display/lt60_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_16|u2_Display/lt60_15  (
    .a({\u2_Display/n1698 ,\u2_Display/n1699 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c15 ),
    .fco(\u2_Display/lt60_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_18|u2_Display/lt60_17  (
    .a({\u2_Display/n1696 ,\u2_Display/n1697 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c17 ),
    .fco(\u2_Display/lt60_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_20|u2_Display/lt60_19  (
    .a({\u2_Display/n1694 ,\u2_Display/n1695 }),
    .b(2'b01),
    .fci(\u2_Display/lt60_c19 ),
    .fco(\u2_Display/lt60_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_22|u2_Display/lt60_21  (
    .a({\u2_Display/n1692 ,\u2_Display/n1693 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c21 ),
    .fco(\u2_Display/lt60_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_24|u2_Display/lt60_23  (
    .a({\u2_Display/n1690 ,\u2_Display/n1691 }),
    .b(2'b10),
    .fci(\u2_Display/lt60_c23 ),
    .fco(\u2_Display/lt60_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_26|u2_Display/lt60_25  (
    .a({\u2_Display/n1688 ,\u2_Display/n1689 }),
    .b(2'b11),
    .fci(\u2_Display/lt60_c25 ),
    .fco(\u2_Display/lt60_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_28|u2_Display/lt60_27  (
    .a({\u2_Display/n1686 ,\u2_Display/n1687 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c27 ),
    .fco(\u2_Display/lt60_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_2|u2_Display/lt60_1  (
    .a({\u2_Display/n1712 ,\u2_Display/n1713 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c1 ),
    .fco(\u2_Display/lt60_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_30|u2_Display/lt60_29  (
    .a({\u2_Display/n1684 ,\u2_Display/n1685 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c29 ),
    .fco(\u2_Display/lt60_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_4|u2_Display/lt60_3  (
    .a({\u2_Display/n1710 ,\u2_Display/n1711 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c3 ),
    .fco(\u2_Display/lt60_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_6|u2_Display/lt60_5  (
    .a({\u2_Display/n1708 ,\u2_Display/n1709 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c5 ),
    .fco(\u2_Display/lt60_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_8|u2_Display/lt60_7  (
    .a({\u2_Display/n1706 ,\u2_Display/n1707 }),
    .b(2'b00),
    .fci(\u2_Display/lt60_c7 ),
    .fco(\u2_Display/lt60_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt60_0|u2_Display/lt60_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt60_cout|u2_Display/lt60_31  (
    .a({1'b0,\u2_Display/n1683 }),
    .b(2'b10),
    .fci(\u2_Display/lt60_c31 ),
    .f({\u2_Display/n1715 ,open_n59239}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_0|u2_Display/lt61_cin  (
    .a({\u2_Display/n1749 ,1'b0}),
    .b({1'b0,open_n59245}),
    .fco(\u2_Display/lt61_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_10|u2_Display/lt61_9  (
    .a({\u2_Display/n1739 ,\u2_Display/n1740 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c9 ),
    .fco(\u2_Display/lt61_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_12|u2_Display/lt61_11  (
    .a({\u2_Display/n1737 ,\u2_Display/n1738 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c11 ),
    .fco(\u2_Display/lt61_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_14|u2_Display/lt61_13  (
    .a({\u2_Display/n1735 ,\u2_Display/n1736 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c13 ),
    .fco(\u2_Display/lt61_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_16|u2_Display/lt61_15  (
    .a({\u2_Display/n1733 ,\u2_Display/n1734 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c15 ),
    .fco(\u2_Display/lt61_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_18|u2_Display/lt61_17  (
    .a({\u2_Display/n1731 ,\u2_Display/n1732 }),
    .b(2'b10),
    .fci(\u2_Display/lt61_c17 ),
    .fco(\u2_Display/lt61_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_20|u2_Display/lt61_19  (
    .a({\u2_Display/n1729 ,\u2_Display/n1730 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c19 ),
    .fco(\u2_Display/lt61_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_22|u2_Display/lt61_21  (
    .a({\u2_Display/n1727 ,\u2_Display/n1728 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c21 ),
    .fco(\u2_Display/lt61_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_24|u2_Display/lt61_23  (
    .a({\u2_Display/n1725 ,\u2_Display/n1726 }),
    .b(2'b11),
    .fci(\u2_Display/lt61_c23 ),
    .fco(\u2_Display/lt61_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_26|u2_Display/lt61_25  (
    .a({\u2_Display/n1723 ,\u2_Display/n1724 }),
    .b(2'b01),
    .fci(\u2_Display/lt61_c25 ),
    .fco(\u2_Display/lt61_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_28|u2_Display/lt61_27  (
    .a({\u2_Display/n1721 ,\u2_Display/n1722 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c27 ),
    .fco(\u2_Display/lt61_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_2|u2_Display/lt61_1  (
    .a({\u2_Display/n1747 ,\u2_Display/n1748 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c1 ),
    .fco(\u2_Display/lt61_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_30|u2_Display/lt61_29  (
    .a({\u2_Display/n1719 ,\u2_Display/n1720 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c29 ),
    .fco(\u2_Display/lt61_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_4|u2_Display/lt61_3  (
    .a({\u2_Display/n1745 ,\u2_Display/n1746 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c3 ),
    .fco(\u2_Display/lt61_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_6|u2_Display/lt61_5  (
    .a({\u2_Display/n1743 ,\u2_Display/n1744 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c5 ),
    .fco(\u2_Display/lt61_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_8|u2_Display/lt61_7  (
    .a({\u2_Display/n1741 ,\u2_Display/n1742 }),
    .b(2'b00),
    .fci(\u2_Display/lt61_c7 ),
    .fco(\u2_Display/lt61_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt61_0|u2_Display/lt61_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt61_cout|u2_Display/lt61_31  (
    .a({1'b0,\u2_Display/n1718 }),
    .b(2'b10),
    .fci(\u2_Display/lt61_c31 ),
    .f({\u2_Display/n1750 ,open_n59649}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_0|u2_Display/lt62_cin  (
    .a({\u2_Display/n1784 ,1'b0}),
    .b({1'b0,open_n59655}),
    .fco(\u2_Display/lt62_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_10|u2_Display/lt62_9  (
    .a({\u2_Display/n1774 ,\u2_Display/n1775 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c9 ),
    .fco(\u2_Display/lt62_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_12|u2_Display/lt62_11  (
    .a({\u2_Display/n1772 ,\u2_Display/n1773 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c11 ),
    .fco(\u2_Display/lt62_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_14|u2_Display/lt62_13  (
    .a({\u2_Display/n1770 ,\u2_Display/n1771 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c13 ),
    .fco(\u2_Display/lt62_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_16|u2_Display/lt62_15  (
    .a({\u2_Display/n1768 ,\u2_Display/n1769 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c15 ),
    .fco(\u2_Display/lt62_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_18|u2_Display/lt62_17  (
    .a({\u2_Display/n1766 ,\u2_Display/n1767 }),
    .b(2'b01),
    .fci(\u2_Display/lt62_c17 ),
    .fco(\u2_Display/lt62_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_20|u2_Display/lt62_19  (
    .a({\u2_Display/n1764 ,\u2_Display/n1765 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c19 ),
    .fco(\u2_Display/lt62_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_22|u2_Display/lt62_21  (
    .a({\u2_Display/n1762 ,\u2_Display/n1763 }),
    .b(2'b10),
    .fci(\u2_Display/lt62_c21 ),
    .fco(\u2_Display/lt62_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_24|u2_Display/lt62_23  (
    .a({\u2_Display/n1760 ,\u2_Display/n1761 }),
    .b(2'b11),
    .fci(\u2_Display/lt62_c23 ),
    .fco(\u2_Display/lt62_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_26|u2_Display/lt62_25  (
    .a({\u2_Display/n1758 ,\u2_Display/n1759 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c25 ),
    .fco(\u2_Display/lt62_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_28|u2_Display/lt62_27  (
    .a({\u2_Display/n1756 ,\u2_Display/n1757 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c27 ),
    .fco(\u2_Display/lt62_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_2|u2_Display/lt62_1  (
    .a({\u2_Display/n1782 ,\u2_Display/n1783 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c1 ),
    .fco(\u2_Display/lt62_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_30|u2_Display/lt62_29  (
    .a({\u2_Display/n1754 ,\u2_Display/n1755 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c29 ),
    .fco(\u2_Display/lt62_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_4|u2_Display/lt62_3  (
    .a({\u2_Display/n1780 ,\u2_Display/n1781 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c3 ),
    .fco(\u2_Display/lt62_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_6|u2_Display/lt62_5  (
    .a({\u2_Display/n1778 ,\u2_Display/n1779 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c5 ),
    .fco(\u2_Display/lt62_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_8|u2_Display/lt62_7  (
    .a({\u2_Display/n1776 ,\u2_Display/n1777 }),
    .b(2'b00),
    .fci(\u2_Display/lt62_c7 ),
    .fco(\u2_Display/lt62_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt62_0|u2_Display/lt62_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt62_cout|u2_Display/lt62_31  (
    .a({1'b0,\u2_Display/n1753 }),
    .b(2'b10),
    .fci(\u2_Display/lt62_c31 ),
    .f({\u2_Display/n1785 ,open_n60059}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_0|u2_Display/lt63_cin  (
    .a({\u2_Display/n1819 ,1'b0}),
    .b({1'b0,open_n60065}),
    .fco(\u2_Display/lt63_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_10|u2_Display/lt63_9  (
    .a({\u2_Display/n1809 ,\u2_Display/n1810 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c9 ),
    .fco(\u2_Display/lt63_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_12|u2_Display/lt63_11  (
    .a({\u2_Display/n1807 ,\u2_Display/n1808 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c11 ),
    .fco(\u2_Display/lt63_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_14|u2_Display/lt63_13  (
    .a({\u2_Display/n1805 ,\u2_Display/n1806 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c13 ),
    .fco(\u2_Display/lt63_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_16|u2_Display/lt63_15  (
    .a({\u2_Display/n1803 ,\u2_Display/n1804 }),
    .b(2'b10),
    .fci(\u2_Display/lt63_c15 ),
    .fco(\u2_Display/lt63_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_18|u2_Display/lt63_17  (
    .a({\u2_Display/n1801 ,\u2_Display/n1802 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c17 ),
    .fco(\u2_Display/lt63_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_20|u2_Display/lt63_19  (
    .a({\u2_Display/n1799 ,\u2_Display/n1800 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c19 ),
    .fco(\u2_Display/lt63_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_22|u2_Display/lt63_21  (
    .a({\u2_Display/n1797 ,\u2_Display/n1798 }),
    .b(2'b11),
    .fci(\u2_Display/lt63_c21 ),
    .fco(\u2_Display/lt63_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_24|u2_Display/lt63_23  (
    .a({\u2_Display/n1795 ,\u2_Display/n1796 }),
    .b(2'b01),
    .fci(\u2_Display/lt63_c23 ),
    .fco(\u2_Display/lt63_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_26|u2_Display/lt63_25  (
    .a({\u2_Display/n1793 ,\u2_Display/n1794 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c25 ),
    .fco(\u2_Display/lt63_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_28|u2_Display/lt63_27  (
    .a({\u2_Display/n1791 ,\u2_Display/n1792 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c27 ),
    .fco(\u2_Display/lt63_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_2|u2_Display/lt63_1  (
    .a({\u2_Display/n1817 ,\u2_Display/n1818 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c1 ),
    .fco(\u2_Display/lt63_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_30|u2_Display/lt63_29  (
    .a({\u2_Display/n1789 ,\u2_Display/n1790 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c29 ),
    .fco(\u2_Display/lt63_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_4|u2_Display/lt63_3  (
    .a({\u2_Display/n1815 ,\u2_Display/n1816 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c3 ),
    .fco(\u2_Display/lt63_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_6|u2_Display/lt63_5  (
    .a({\u2_Display/n1813 ,\u2_Display/n1814 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c5 ),
    .fco(\u2_Display/lt63_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_8|u2_Display/lt63_7  (
    .a({\u2_Display/n1811 ,\u2_Display/n1812 }),
    .b(2'b00),
    .fci(\u2_Display/lt63_c7 ),
    .fco(\u2_Display/lt63_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt63_0|u2_Display/lt63_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt63_cout|u2_Display/lt63_31  (
    .a({1'b0,\u2_Display/n1788 }),
    .b(2'b10),
    .fci(\u2_Display/lt63_c31 ),
    .f({\u2_Display/n1820 ,open_n60469}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_0|u2_Display/lt64_cin  (
    .a({\u2_Display/n1854 ,1'b0}),
    .b({1'b0,open_n60475}),
    .fco(\u2_Display/lt64_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_10|u2_Display/lt64_9  (
    .a({\u2_Display/n1844 ,\u2_Display/n1845 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c9 ),
    .fco(\u2_Display/lt64_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_12|u2_Display/lt64_11  (
    .a({\u2_Display/n1842 ,\u2_Display/n1843 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c11 ),
    .fco(\u2_Display/lt64_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_14|u2_Display/lt64_13  (
    .a({\u2_Display/n1840 ,\u2_Display/n1841 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c13 ),
    .fco(\u2_Display/lt64_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_16|u2_Display/lt64_15  (
    .a({\u2_Display/n1838 ,\u2_Display/n1839 }),
    .b(2'b01),
    .fci(\u2_Display/lt64_c15 ),
    .fco(\u2_Display/lt64_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_18|u2_Display/lt64_17  (
    .a({\u2_Display/n1836 ,\u2_Display/n1837 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c17 ),
    .fco(\u2_Display/lt64_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_20|u2_Display/lt64_19  (
    .a({\u2_Display/n1834 ,\u2_Display/n1835 }),
    .b(2'b10),
    .fci(\u2_Display/lt64_c19 ),
    .fco(\u2_Display/lt64_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_22|u2_Display/lt64_21  (
    .a({\u2_Display/n1832 ,\u2_Display/n1833 }),
    .b(2'b11),
    .fci(\u2_Display/lt64_c21 ),
    .fco(\u2_Display/lt64_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_24|u2_Display/lt64_23  (
    .a({\u2_Display/n1830 ,\u2_Display/n1831 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c23 ),
    .fco(\u2_Display/lt64_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_26|u2_Display/lt64_25  (
    .a({\u2_Display/n1828 ,\u2_Display/n1829 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c25 ),
    .fco(\u2_Display/lt64_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_28|u2_Display/lt64_27  (
    .a({\u2_Display/n1826 ,\u2_Display/n1827 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c27 ),
    .fco(\u2_Display/lt64_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_2|u2_Display/lt64_1  (
    .a({\u2_Display/n1852 ,\u2_Display/n1853 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c1 ),
    .fco(\u2_Display/lt64_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_30|u2_Display/lt64_29  (
    .a({\u2_Display/n1824 ,\u2_Display/n1825 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c29 ),
    .fco(\u2_Display/lt64_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_4|u2_Display/lt64_3  (
    .a({\u2_Display/n1850 ,\u2_Display/n1851 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c3 ),
    .fco(\u2_Display/lt64_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_6|u2_Display/lt64_5  (
    .a({\u2_Display/n1848 ,\u2_Display/n1849 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c5 ),
    .fco(\u2_Display/lt64_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_8|u2_Display/lt64_7  (
    .a({\u2_Display/n1846 ,\u2_Display/n1847 }),
    .b(2'b00),
    .fci(\u2_Display/lt64_c7 ),
    .fco(\u2_Display/lt64_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt64_0|u2_Display/lt64_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt64_cout|u2_Display/lt64_31  (
    .a({1'b0,\u2_Display/n1823 }),
    .b(2'b10),
    .fci(\u2_Display/lt64_c31 ),
    .f({\u2_Display/n1855 ,open_n60879}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_0|u2_Display/lt65_cin  (
    .a({\u2_Display/n1889 ,1'b0}),
    .b({1'b0,open_n60885}),
    .fco(\u2_Display/lt65_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_10|u2_Display/lt65_9  (
    .a({\u2_Display/n1879 ,\u2_Display/n1880 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c9 ),
    .fco(\u2_Display/lt65_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_12|u2_Display/lt65_11  (
    .a({\u2_Display/n1877 ,\u2_Display/n1878 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c11 ),
    .fco(\u2_Display/lt65_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_14|u2_Display/lt65_13  (
    .a({\u2_Display/n1875 ,\u2_Display/n1876 }),
    .b(2'b10),
    .fci(\u2_Display/lt65_c13 ),
    .fco(\u2_Display/lt65_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_16|u2_Display/lt65_15  (
    .a({\u2_Display/n1873 ,\u2_Display/n1874 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c15 ),
    .fco(\u2_Display/lt65_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_18|u2_Display/lt65_17  (
    .a({\u2_Display/n1871 ,\u2_Display/n1872 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c17 ),
    .fco(\u2_Display/lt65_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_20|u2_Display/lt65_19  (
    .a({\u2_Display/n1869 ,\u2_Display/n1870 }),
    .b(2'b11),
    .fci(\u2_Display/lt65_c19 ),
    .fco(\u2_Display/lt65_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_22|u2_Display/lt65_21  (
    .a({\u2_Display/n1867 ,\u2_Display/n1868 }),
    .b(2'b01),
    .fci(\u2_Display/lt65_c21 ),
    .fco(\u2_Display/lt65_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_24|u2_Display/lt65_23  (
    .a({\u2_Display/n1865 ,\u2_Display/n1866 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c23 ),
    .fco(\u2_Display/lt65_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_26|u2_Display/lt65_25  (
    .a({\u2_Display/n1863 ,\u2_Display/n1864 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c25 ),
    .fco(\u2_Display/lt65_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_28|u2_Display/lt65_27  (
    .a({\u2_Display/n1861 ,\u2_Display/n1862 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c27 ),
    .fco(\u2_Display/lt65_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_2|u2_Display/lt65_1  (
    .a({\u2_Display/n1887 ,\u2_Display/n1888 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c1 ),
    .fco(\u2_Display/lt65_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_30|u2_Display/lt65_29  (
    .a({\u2_Display/n1859 ,\u2_Display/n1860 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c29 ),
    .fco(\u2_Display/lt65_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_4|u2_Display/lt65_3  (
    .a({\u2_Display/n1885 ,\u2_Display/n1886 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c3 ),
    .fco(\u2_Display/lt65_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_6|u2_Display/lt65_5  (
    .a({\u2_Display/n1883 ,\u2_Display/n1884 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c5 ),
    .fco(\u2_Display/lt65_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_8|u2_Display/lt65_7  (
    .a({\u2_Display/n1881 ,\u2_Display/n1882 }),
    .b(2'b00),
    .fci(\u2_Display/lt65_c7 ),
    .fco(\u2_Display/lt65_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt65_0|u2_Display/lt65_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt65_cout|u2_Display/lt65_31  (
    .a({1'b0,\u2_Display/n1858 }),
    .b(2'b10),
    .fci(\u2_Display/lt65_c31 ),
    .f({\u2_Display/n1890 ,open_n61289}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_0|u2_Display/lt66_cin  (
    .a({\u2_Display/n1924 ,1'b0}),
    .b({1'b0,open_n61295}),
    .fco(\u2_Display/lt66_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_10|u2_Display/lt66_9  (
    .a({\u2_Display/n1914 ,\u2_Display/n1915 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c9 ),
    .fco(\u2_Display/lt66_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_12|u2_Display/lt66_11  (
    .a({\u2_Display/n1912 ,\u2_Display/n1913 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c11 ),
    .fco(\u2_Display/lt66_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_14|u2_Display/lt66_13  (
    .a({\u2_Display/n1910 ,\u2_Display/n1911 }),
    .b(2'b01),
    .fci(\u2_Display/lt66_c13 ),
    .fco(\u2_Display/lt66_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_16|u2_Display/lt66_15  (
    .a({\u2_Display/n1908 ,\u2_Display/n1909 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c15 ),
    .fco(\u2_Display/lt66_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_18|u2_Display/lt66_17  (
    .a({\u2_Display/n1906 ,\u2_Display/n1907 }),
    .b(2'b10),
    .fci(\u2_Display/lt66_c17 ),
    .fco(\u2_Display/lt66_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_20|u2_Display/lt66_19  (
    .a({\u2_Display/n1904 ,\u2_Display/n1905 }),
    .b(2'b11),
    .fci(\u2_Display/lt66_c19 ),
    .fco(\u2_Display/lt66_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_22|u2_Display/lt66_21  (
    .a({\u2_Display/n1902 ,\u2_Display/n1903 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c21 ),
    .fco(\u2_Display/lt66_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_24|u2_Display/lt66_23  (
    .a({\u2_Display/n1900 ,\u2_Display/n1901 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c23 ),
    .fco(\u2_Display/lt66_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_26|u2_Display/lt66_25  (
    .a({\u2_Display/n1898 ,\u2_Display/n1899 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c25 ),
    .fco(\u2_Display/lt66_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_28|u2_Display/lt66_27  (
    .a({\u2_Display/n1896 ,\u2_Display/n1897 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c27 ),
    .fco(\u2_Display/lt66_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_2|u2_Display/lt66_1  (
    .a({\u2_Display/n1922 ,\u2_Display/n1923 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c1 ),
    .fco(\u2_Display/lt66_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_30|u2_Display/lt66_29  (
    .a({\u2_Display/n1894 ,\u2_Display/n1895 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c29 ),
    .fco(\u2_Display/lt66_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_4|u2_Display/lt66_3  (
    .a({\u2_Display/n1920 ,\u2_Display/n1921 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c3 ),
    .fco(\u2_Display/lt66_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_6|u2_Display/lt66_5  (
    .a({\u2_Display/n1918 ,\u2_Display/n1919 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c5 ),
    .fco(\u2_Display/lt66_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_8|u2_Display/lt66_7  (
    .a({\u2_Display/n1916 ,\u2_Display/n1917 }),
    .b(2'b00),
    .fci(\u2_Display/lt66_c7 ),
    .fco(\u2_Display/lt66_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt66_0|u2_Display/lt66_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt66_cout|u2_Display/lt66_31  (
    .a({1'b0,\u2_Display/n1893 }),
    .b(2'b10),
    .fci(\u2_Display/lt66_c31 ),
    .f({\u2_Display/n1925 ,open_n61699}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_0|u2_Display/lt67_cin  (
    .a({\u2_Display/n1959 ,1'b0}),
    .b({1'b0,open_n61705}),
    .fco(\u2_Display/lt67_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_10|u2_Display/lt67_9  (
    .a({\u2_Display/n1949 ,\u2_Display/n1950 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c9 ),
    .fco(\u2_Display/lt67_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_12|u2_Display/lt67_11  (
    .a({\u2_Display/n1947 ,\u2_Display/n1948 }),
    .b(2'b10),
    .fci(\u2_Display/lt67_c11 ),
    .fco(\u2_Display/lt67_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_14|u2_Display/lt67_13  (
    .a({\u2_Display/n1945 ,\u2_Display/n1946 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c13 ),
    .fco(\u2_Display/lt67_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_16|u2_Display/lt67_15  (
    .a({\u2_Display/n1943 ,\u2_Display/n1944 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c15 ),
    .fco(\u2_Display/lt67_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_18|u2_Display/lt67_17  (
    .a({\u2_Display/n1941 ,\u2_Display/n1942 }),
    .b(2'b11),
    .fci(\u2_Display/lt67_c17 ),
    .fco(\u2_Display/lt67_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_20|u2_Display/lt67_19  (
    .a({\u2_Display/n1939 ,\u2_Display/n1940 }),
    .b(2'b01),
    .fci(\u2_Display/lt67_c19 ),
    .fco(\u2_Display/lt67_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_22|u2_Display/lt67_21  (
    .a({\u2_Display/n1937 ,\u2_Display/n1938 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c21 ),
    .fco(\u2_Display/lt67_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_24|u2_Display/lt67_23  (
    .a({\u2_Display/n1935 ,\u2_Display/n1936 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c23 ),
    .fco(\u2_Display/lt67_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_26|u2_Display/lt67_25  (
    .a({\u2_Display/n1933 ,\u2_Display/n1934 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c25 ),
    .fco(\u2_Display/lt67_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_28|u2_Display/lt67_27  (
    .a({\u2_Display/n1931 ,\u2_Display/n1932 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c27 ),
    .fco(\u2_Display/lt67_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_2|u2_Display/lt67_1  (
    .a({\u2_Display/n1957 ,\u2_Display/n1958 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c1 ),
    .fco(\u2_Display/lt67_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_30|u2_Display/lt67_29  (
    .a({\u2_Display/n1929 ,\u2_Display/n1930 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c29 ),
    .fco(\u2_Display/lt67_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_4|u2_Display/lt67_3  (
    .a({\u2_Display/n1955 ,\u2_Display/n1956 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c3 ),
    .fco(\u2_Display/lt67_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_6|u2_Display/lt67_5  (
    .a({\u2_Display/n1953 ,\u2_Display/n1954 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c5 ),
    .fco(\u2_Display/lt67_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_8|u2_Display/lt67_7  (
    .a({\u2_Display/n1951 ,\u2_Display/n1952 }),
    .b(2'b00),
    .fci(\u2_Display/lt67_c7 ),
    .fco(\u2_Display/lt67_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt67_0|u2_Display/lt67_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt67_cout|u2_Display/lt67_31  (
    .a({1'b0,\u2_Display/n1928 }),
    .b(2'b10),
    .fci(\u2_Display/lt67_c31 ),
    .f({\u2_Display/n1960 ,open_n62109}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_0|u2_Display/lt68_cin  (
    .a({\u2_Display/n1994 ,1'b0}),
    .b({1'b0,open_n62115}),
    .fco(\u2_Display/lt68_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_10|u2_Display/lt68_9  (
    .a({\u2_Display/n1984 ,\u2_Display/n1985 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c9 ),
    .fco(\u2_Display/lt68_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_12|u2_Display/lt68_11  (
    .a({\u2_Display/n1982 ,\u2_Display/n1983 }),
    .b(2'b01),
    .fci(\u2_Display/lt68_c11 ),
    .fco(\u2_Display/lt68_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_14|u2_Display/lt68_13  (
    .a({\u2_Display/n1980 ,\u2_Display/n1981 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c13 ),
    .fco(\u2_Display/lt68_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_16|u2_Display/lt68_15  (
    .a({\u2_Display/n1978 ,\u2_Display/n1979 }),
    .b(2'b10),
    .fci(\u2_Display/lt68_c15 ),
    .fco(\u2_Display/lt68_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_18|u2_Display/lt68_17  (
    .a({\u2_Display/n1976 ,\u2_Display/n1977 }),
    .b(2'b11),
    .fci(\u2_Display/lt68_c17 ),
    .fco(\u2_Display/lt68_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_20|u2_Display/lt68_19  (
    .a({\u2_Display/n1974 ,\u2_Display/n1975 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c19 ),
    .fco(\u2_Display/lt68_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_22|u2_Display/lt68_21  (
    .a({\u2_Display/n1972 ,\u2_Display/n1973 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c21 ),
    .fco(\u2_Display/lt68_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_24|u2_Display/lt68_23  (
    .a({\u2_Display/n1970 ,\u2_Display/n1971 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c23 ),
    .fco(\u2_Display/lt68_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_26|u2_Display/lt68_25  (
    .a({\u2_Display/n1968 ,\u2_Display/n1969 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c25 ),
    .fco(\u2_Display/lt68_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_28|u2_Display/lt68_27  (
    .a({\u2_Display/n1966 ,\u2_Display/n1967 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c27 ),
    .fco(\u2_Display/lt68_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_2|u2_Display/lt68_1  (
    .a({\u2_Display/n1992 ,\u2_Display/n1993 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c1 ),
    .fco(\u2_Display/lt68_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_30|u2_Display/lt68_29  (
    .a({\u2_Display/n1964 ,\u2_Display/n1965 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c29 ),
    .fco(\u2_Display/lt68_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_4|u2_Display/lt68_3  (
    .a({\u2_Display/n1990 ,\u2_Display/n1991 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c3 ),
    .fco(\u2_Display/lt68_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_6|u2_Display/lt68_5  (
    .a({\u2_Display/n1988 ,\u2_Display/n1989 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c5 ),
    .fco(\u2_Display/lt68_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_8|u2_Display/lt68_7  (
    .a({\u2_Display/n1986 ,\u2_Display/n1987 }),
    .b(2'b00),
    .fci(\u2_Display/lt68_c7 ),
    .fco(\u2_Display/lt68_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt68_0|u2_Display/lt68_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt68_cout|u2_Display/lt68_31  (
    .a({1'b0,\u2_Display/n1963 }),
    .b(2'b10),
    .fci(\u2_Display/lt68_c31 ),
    .f({\u2_Display/n1995 ,open_n62519}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_0|u2_Display/lt69_cin  (
    .a({\u2_Display/n2029 ,1'b0}),
    .b({1'b0,open_n62525}),
    .fco(\u2_Display/lt69_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_10|u2_Display/lt69_9  (
    .a({\u2_Display/n2019 ,\u2_Display/n2020 }),
    .b(2'b10),
    .fci(\u2_Display/lt69_c9 ),
    .fco(\u2_Display/lt69_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_12|u2_Display/lt69_11  (
    .a({\u2_Display/n2017 ,\u2_Display/n2018 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c11 ),
    .fco(\u2_Display/lt69_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_14|u2_Display/lt69_13  (
    .a({\u2_Display/n2015 ,\u2_Display/n2016 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c13 ),
    .fco(\u2_Display/lt69_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_16|u2_Display/lt69_15  (
    .a({\u2_Display/n2013 ,\u2_Display/n2014 }),
    .b(2'b11),
    .fci(\u2_Display/lt69_c15 ),
    .fco(\u2_Display/lt69_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_18|u2_Display/lt69_17  (
    .a({\u2_Display/n2011 ,\u2_Display/n2012 }),
    .b(2'b01),
    .fci(\u2_Display/lt69_c17 ),
    .fco(\u2_Display/lt69_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_20|u2_Display/lt69_19  (
    .a({\u2_Display/n2009 ,\u2_Display/n2010 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c19 ),
    .fco(\u2_Display/lt69_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_22|u2_Display/lt69_21  (
    .a({\u2_Display/n2007 ,\u2_Display/n2008 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c21 ),
    .fco(\u2_Display/lt69_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_24|u2_Display/lt69_23  (
    .a({\u2_Display/n2005 ,\u2_Display/n2006 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c23 ),
    .fco(\u2_Display/lt69_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_26|u2_Display/lt69_25  (
    .a({\u2_Display/n2003 ,\u2_Display/n2004 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c25 ),
    .fco(\u2_Display/lt69_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_28|u2_Display/lt69_27  (
    .a({\u2_Display/n2001 ,\u2_Display/n2002 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c27 ),
    .fco(\u2_Display/lt69_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_2|u2_Display/lt69_1  (
    .a({\u2_Display/n2027 ,\u2_Display/n2028 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c1 ),
    .fco(\u2_Display/lt69_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_30|u2_Display/lt69_29  (
    .a({\u2_Display/n1999 ,\u2_Display/n2000 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c29 ),
    .fco(\u2_Display/lt69_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_4|u2_Display/lt69_3  (
    .a({\u2_Display/n2025 ,\u2_Display/n2026 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c3 ),
    .fco(\u2_Display/lt69_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_6|u2_Display/lt69_5  (
    .a({\u2_Display/n2023 ,\u2_Display/n2024 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c5 ),
    .fco(\u2_Display/lt69_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_8|u2_Display/lt69_7  (
    .a({\u2_Display/n2021 ,\u2_Display/n2022 }),
    .b(2'b00),
    .fci(\u2_Display/lt69_c7 ),
    .fco(\u2_Display/lt69_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt69_0|u2_Display/lt69_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt69_cout|u2_Display/lt69_31  (
    .a({1'b0,\u2_Display/n1998 }),
    .b(2'b10),
    .fci(\u2_Display/lt69_c31 ),
    .f({\u2_Display/n2030 ,open_n62929}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_0|u2_Display/lt6_2_cin  (
    .a({lcd_ypos[0],1'b0}),
    .b({\u2_Display/j [0],open_n62935}),
    .fco(\u2_Display/lt6_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_10|u2_Display/lt6_2_9  (
    .a(lcd_ypos[10:9]),
    .b({\u2_Display/j [9],\u2_Display/n99 [0]}),
    .fci(\u2_Display/lt6_2_c9 ),
    .fco(\u2_Display/lt6_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_2|u2_Display/lt6_2_1  (
    .a(lcd_ypos[2:1]),
    .b(\u2_Display/j [2:1]),
    .fci(\u2_Display/lt6_2_c1 ),
    .fco(\u2_Display/lt6_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_4|u2_Display/lt6_2_3  (
    .a(lcd_ypos[4:3]),
    .b(\u2_Display/j [4:3]),
    .fci(\u2_Display/lt6_2_c3 ),
    .fco(\u2_Display/lt6_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_6|u2_Display/lt6_2_5  (
    .a(lcd_ypos[6:5]),
    .b(\u2_Display/j [6:5]),
    .fci(\u2_Display/lt6_2_c5 ),
    .fco(\u2_Display/lt6_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_8|u2_Display/lt6_2_7  (
    .a(lcd_ypos[8:7]),
    .b(\u2_Display/j [8:7]),
    .fci(\u2_Display/lt6_2_c7 ),
    .fco(\u2_Display/lt6_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt6_2_0|u2_Display/lt6_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt6_2_cout|u2_Display/lt6_2_11  (
    .a({1'b0,lcd_ypos[11]}),
    .b(2'b10),
    .fci(\u2_Display/lt6_2_c11 ),
    .f({\u2_Display/n100 ,open_n63099}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_0|u2_Display/lt70_cin  (
    .a({\u2_Display/n2064 ,1'b0}),
    .b({1'b0,open_n63105}),
    .fco(\u2_Display/lt70_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_10|u2_Display/lt70_9  (
    .a({\u2_Display/n2054 ,\u2_Display/n2055 }),
    .b(2'b01),
    .fci(\u2_Display/lt70_c9 ),
    .fco(\u2_Display/lt70_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_12|u2_Display/lt70_11  (
    .a({\u2_Display/n2052 ,\u2_Display/n2053 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c11 ),
    .fco(\u2_Display/lt70_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_14|u2_Display/lt70_13  (
    .a({\u2_Display/n2050 ,\u2_Display/n2051 }),
    .b(2'b10),
    .fci(\u2_Display/lt70_c13 ),
    .fco(\u2_Display/lt70_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_16|u2_Display/lt70_15  (
    .a({\u2_Display/n2048 ,\u2_Display/n2049 }),
    .b(2'b11),
    .fci(\u2_Display/lt70_c15 ),
    .fco(\u2_Display/lt70_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_18|u2_Display/lt70_17  (
    .a({\u2_Display/n2046 ,\u2_Display/n2047 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c17 ),
    .fco(\u2_Display/lt70_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_20|u2_Display/lt70_19  (
    .a({\u2_Display/n2044 ,\u2_Display/n2045 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c19 ),
    .fco(\u2_Display/lt70_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_22|u2_Display/lt70_21  (
    .a({\u2_Display/n2042 ,\u2_Display/n2043 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c21 ),
    .fco(\u2_Display/lt70_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_24|u2_Display/lt70_23  (
    .a({\u2_Display/n2040 ,\u2_Display/n2041 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c23 ),
    .fco(\u2_Display/lt70_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_26|u2_Display/lt70_25  (
    .a({\u2_Display/n2038 ,\u2_Display/n2039 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c25 ),
    .fco(\u2_Display/lt70_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_28|u2_Display/lt70_27  (
    .a({\u2_Display/n2036 ,\u2_Display/n2037 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c27 ),
    .fco(\u2_Display/lt70_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_2|u2_Display/lt70_1  (
    .a({\u2_Display/n2062 ,\u2_Display/n2063 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c1 ),
    .fco(\u2_Display/lt70_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_30|u2_Display/lt70_29  (
    .a({\u2_Display/n2034 ,\u2_Display/n2035 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c29 ),
    .fco(\u2_Display/lt70_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_4|u2_Display/lt70_3  (
    .a({\u2_Display/n2060 ,\u2_Display/n2061 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c3 ),
    .fco(\u2_Display/lt70_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_6|u2_Display/lt70_5  (
    .a({\u2_Display/n2058 ,\u2_Display/n2059 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c5 ),
    .fco(\u2_Display/lt70_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_8|u2_Display/lt70_7  (
    .a({\u2_Display/n2056 ,\u2_Display/n2057 }),
    .b(2'b00),
    .fci(\u2_Display/lt70_c7 ),
    .fco(\u2_Display/lt70_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt70_0|u2_Display/lt70_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt70_cout|u2_Display/lt70_31  (
    .a({1'b0,\u2_Display/n2033 }),
    .b(2'b10),
    .fci(\u2_Display/lt70_c31 ),
    .f({\u2_Display/n2065 ,open_n63509}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_0|u2_Display/lt71_cin  (
    .a({\u2_Display/n2099 ,1'b0}),
    .b({1'b0,open_n63515}),
    .fco(\u2_Display/lt71_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_10|u2_Display/lt71_9  (
    .a({\u2_Display/n2089 ,\u2_Display/n2090 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c9 ),
    .fco(\u2_Display/lt71_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_12|u2_Display/lt71_11  (
    .a({\u2_Display/n2087 ,\u2_Display/n2088 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c11 ),
    .fco(\u2_Display/lt71_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_14|u2_Display/lt71_13  (
    .a({\u2_Display/n2085 ,\u2_Display/n2086 }),
    .b(2'b11),
    .fci(\u2_Display/lt71_c13 ),
    .fco(\u2_Display/lt71_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_16|u2_Display/lt71_15  (
    .a({\u2_Display/n2083 ,\u2_Display/n2084 }),
    .b(2'b01),
    .fci(\u2_Display/lt71_c15 ),
    .fco(\u2_Display/lt71_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_18|u2_Display/lt71_17  (
    .a({\u2_Display/n2081 ,\u2_Display/n2082 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c17 ),
    .fco(\u2_Display/lt71_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_20|u2_Display/lt71_19  (
    .a({\u2_Display/n2079 ,\u2_Display/n2080 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c19 ),
    .fco(\u2_Display/lt71_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_22|u2_Display/lt71_21  (
    .a({\u2_Display/n2077 ,\u2_Display/n2078 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c21 ),
    .fco(\u2_Display/lt71_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_24|u2_Display/lt71_23  (
    .a({\u2_Display/n2075 ,\u2_Display/n2076 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c23 ),
    .fco(\u2_Display/lt71_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_26|u2_Display/lt71_25  (
    .a({\u2_Display/n2073 ,\u2_Display/n2074 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c25 ),
    .fco(\u2_Display/lt71_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_28|u2_Display/lt71_27  (
    .a({\u2_Display/n2071 ,\u2_Display/n2072 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c27 ),
    .fco(\u2_Display/lt71_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_2|u2_Display/lt71_1  (
    .a({\u2_Display/n2097 ,\u2_Display/n2098 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c1 ),
    .fco(\u2_Display/lt71_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_30|u2_Display/lt71_29  (
    .a({\u2_Display/n2069 ,\u2_Display/n2070 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c29 ),
    .fco(\u2_Display/lt71_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_4|u2_Display/lt71_3  (
    .a({\u2_Display/n2095 ,\u2_Display/n2096 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c3 ),
    .fco(\u2_Display/lt71_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_6|u2_Display/lt71_5  (
    .a({\u2_Display/n2093 ,\u2_Display/n2094 }),
    .b(2'b00),
    .fci(\u2_Display/lt71_c5 ),
    .fco(\u2_Display/lt71_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_8|u2_Display/lt71_7  (
    .a({\u2_Display/n2091 ,\u2_Display/n2092 }),
    .b(2'b10),
    .fci(\u2_Display/lt71_c7 ),
    .fco(\u2_Display/lt71_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt71_0|u2_Display/lt71_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt71_cout|u2_Display/lt71_31  (
    .a({1'b0,\u2_Display/n2068 }),
    .b(2'b10),
    .fci(\u2_Display/lt71_c31 ),
    .f({\u2_Display/n2100 ,open_n63919}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_0|u2_Display/lt72_cin  (
    .a({\u2_Display/n2134 ,1'b0}),
    .b({1'b0,open_n63925}),
    .fco(\u2_Display/lt72_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_10|u2_Display/lt72_9  (
    .a({\u2_Display/n2124 ,\u2_Display/n2125 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c9 ),
    .fco(\u2_Display/lt72_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_12|u2_Display/lt72_11  (
    .a({\u2_Display/n2122 ,\u2_Display/n2123 }),
    .b(2'b10),
    .fci(\u2_Display/lt72_c11 ),
    .fco(\u2_Display/lt72_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_14|u2_Display/lt72_13  (
    .a({\u2_Display/n2120 ,\u2_Display/n2121 }),
    .b(2'b11),
    .fci(\u2_Display/lt72_c13 ),
    .fco(\u2_Display/lt72_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_16|u2_Display/lt72_15  (
    .a({\u2_Display/n2118 ,\u2_Display/n2119 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c15 ),
    .fco(\u2_Display/lt72_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_18|u2_Display/lt72_17  (
    .a({\u2_Display/n2116 ,\u2_Display/n2117 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c17 ),
    .fco(\u2_Display/lt72_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_20|u2_Display/lt72_19  (
    .a({\u2_Display/n2114 ,\u2_Display/n2115 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c19 ),
    .fco(\u2_Display/lt72_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_22|u2_Display/lt72_21  (
    .a({\u2_Display/n2112 ,\u2_Display/n2113 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c21 ),
    .fco(\u2_Display/lt72_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_24|u2_Display/lt72_23  (
    .a({\u2_Display/n2110 ,\u2_Display/n2111 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c23 ),
    .fco(\u2_Display/lt72_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_26|u2_Display/lt72_25  (
    .a({\u2_Display/n2108 ,\u2_Display/n2109 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c25 ),
    .fco(\u2_Display/lt72_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_28|u2_Display/lt72_27  (
    .a({\u2_Display/n2106 ,\u2_Display/n2107 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c27 ),
    .fco(\u2_Display/lt72_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_2|u2_Display/lt72_1  (
    .a({\u2_Display/n2132 ,\u2_Display/n2133 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c1 ),
    .fco(\u2_Display/lt72_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_30|u2_Display/lt72_29  (
    .a({\u2_Display/n2104 ,\u2_Display/n2105 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c29 ),
    .fco(\u2_Display/lt72_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_4|u2_Display/lt72_3  (
    .a({\u2_Display/n2130 ,\u2_Display/n2131 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c3 ),
    .fco(\u2_Display/lt72_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_6|u2_Display/lt72_5  (
    .a({\u2_Display/n2128 ,\u2_Display/n2129 }),
    .b(2'b00),
    .fci(\u2_Display/lt72_c5 ),
    .fco(\u2_Display/lt72_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_8|u2_Display/lt72_7  (
    .a({\u2_Display/n2126 ,\u2_Display/n2127 }),
    .b(2'b01),
    .fci(\u2_Display/lt72_c7 ),
    .fco(\u2_Display/lt72_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt72_0|u2_Display/lt72_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt72_cout|u2_Display/lt72_31  (
    .a({1'b0,\u2_Display/n2103 }),
    .b(2'b10),
    .fci(\u2_Display/lt72_c31 ),
    .f({\u2_Display/n2135 ,open_n64329}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_0|u2_Display/lt73_cin  (
    .a({\u2_Display/n2169 ,1'b0}),
    .b({1'b0,open_n64335}),
    .fco(\u2_Display/lt73_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_10|u2_Display/lt73_9  (
    .a({\u2_Display/n2159 ,\u2_Display/n2160 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c9 ),
    .fco(\u2_Display/lt73_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_12|u2_Display/lt73_11  (
    .a({\u2_Display/n2157 ,\u2_Display/n2158 }),
    .b(2'b11),
    .fci(\u2_Display/lt73_c11 ),
    .fco(\u2_Display/lt73_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_14|u2_Display/lt73_13  (
    .a({\u2_Display/n2155 ,\u2_Display/n2156 }),
    .b(2'b01),
    .fci(\u2_Display/lt73_c13 ),
    .fco(\u2_Display/lt73_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_16|u2_Display/lt73_15  (
    .a({\u2_Display/n2153 ,\u2_Display/n2154 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c15 ),
    .fco(\u2_Display/lt73_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_18|u2_Display/lt73_17  (
    .a({\u2_Display/n2151 ,\u2_Display/n2152 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c17 ),
    .fco(\u2_Display/lt73_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_20|u2_Display/lt73_19  (
    .a({\u2_Display/n2149 ,\u2_Display/n2150 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c19 ),
    .fco(\u2_Display/lt73_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_22|u2_Display/lt73_21  (
    .a({\u2_Display/n2147 ,\u2_Display/n2148 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c21 ),
    .fco(\u2_Display/lt73_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_24|u2_Display/lt73_23  (
    .a({\u2_Display/n2145 ,\u2_Display/n2146 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c23 ),
    .fco(\u2_Display/lt73_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_26|u2_Display/lt73_25  (
    .a({\u2_Display/n2143 ,\u2_Display/n2144 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c25 ),
    .fco(\u2_Display/lt73_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_28|u2_Display/lt73_27  (
    .a({\u2_Display/n2141 ,\u2_Display/n2142 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c27 ),
    .fco(\u2_Display/lt73_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_2|u2_Display/lt73_1  (
    .a({\u2_Display/n2167 ,\u2_Display/n2168 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c1 ),
    .fco(\u2_Display/lt73_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_30|u2_Display/lt73_29  (
    .a({\u2_Display/n2139 ,\u2_Display/n2140 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c29 ),
    .fco(\u2_Display/lt73_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_4|u2_Display/lt73_3  (
    .a({\u2_Display/n2165 ,\u2_Display/n2166 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c3 ),
    .fco(\u2_Display/lt73_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_6|u2_Display/lt73_5  (
    .a({\u2_Display/n2163 ,\u2_Display/n2164 }),
    .b(2'b10),
    .fci(\u2_Display/lt73_c5 ),
    .fco(\u2_Display/lt73_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_8|u2_Display/lt73_7  (
    .a({\u2_Display/n2161 ,\u2_Display/n2162 }),
    .b(2'b00),
    .fci(\u2_Display/lt73_c7 ),
    .fco(\u2_Display/lt73_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt73_0|u2_Display/lt73_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt73_cout|u2_Display/lt73_31  (
    .a({1'b0,\u2_Display/n2138 }),
    .b(2'b10),
    .fci(\u2_Display/lt73_c31 ),
    .f({\u2_Display/n2170 ,open_n64739}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_0|u2_Display/lt74_cin  (
    .a({\u2_Display/n2204 ,1'b0}),
    .b({1'b0,open_n64745}),
    .fco(\u2_Display/lt74_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_10|u2_Display/lt74_9  (
    .a({\u2_Display/n2194 ,\u2_Display/n2195 }),
    .b(2'b10),
    .fci(\u2_Display/lt74_c9 ),
    .fco(\u2_Display/lt74_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_12|u2_Display/lt74_11  (
    .a({\u2_Display/n2192 ,\u2_Display/n2193 }),
    .b(2'b11),
    .fci(\u2_Display/lt74_c11 ),
    .fco(\u2_Display/lt74_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_14|u2_Display/lt74_13  (
    .a({\u2_Display/n2190 ,\u2_Display/n2191 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c13 ),
    .fco(\u2_Display/lt74_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_16|u2_Display/lt74_15  (
    .a({\u2_Display/n2188 ,\u2_Display/n2189 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c15 ),
    .fco(\u2_Display/lt74_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_18|u2_Display/lt74_17  (
    .a({\u2_Display/n2186 ,\u2_Display/n2187 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c17 ),
    .fco(\u2_Display/lt74_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_20|u2_Display/lt74_19  (
    .a({\u2_Display/n2184 ,\u2_Display/n2185 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c19 ),
    .fco(\u2_Display/lt74_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_22|u2_Display/lt74_21  (
    .a({\u2_Display/n2182 ,\u2_Display/n2183 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c21 ),
    .fco(\u2_Display/lt74_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_24|u2_Display/lt74_23  (
    .a({\u2_Display/n2180 ,\u2_Display/n2181 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c23 ),
    .fco(\u2_Display/lt74_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_26|u2_Display/lt74_25  (
    .a({\u2_Display/n2178 ,\u2_Display/n2179 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c25 ),
    .fco(\u2_Display/lt74_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_28|u2_Display/lt74_27  (
    .a({\u2_Display/n2176 ,\u2_Display/n2177 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c27 ),
    .fco(\u2_Display/lt74_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_2|u2_Display/lt74_1  (
    .a({\u2_Display/n2202 ,\u2_Display/n2203 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c1 ),
    .fco(\u2_Display/lt74_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_30|u2_Display/lt74_29  (
    .a({\u2_Display/n2174 ,\u2_Display/n2175 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c29 ),
    .fco(\u2_Display/lt74_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_4|u2_Display/lt74_3  (
    .a({\u2_Display/n2200 ,\u2_Display/n2201 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c3 ),
    .fco(\u2_Display/lt74_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_6|u2_Display/lt74_5  (
    .a({\u2_Display/n2198 ,\u2_Display/n2199 }),
    .b(2'b01),
    .fci(\u2_Display/lt74_c5 ),
    .fco(\u2_Display/lt74_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_8|u2_Display/lt74_7  (
    .a({\u2_Display/n2196 ,\u2_Display/n2197 }),
    .b(2'b00),
    .fci(\u2_Display/lt74_c7 ),
    .fco(\u2_Display/lt74_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt74_0|u2_Display/lt74_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt74_cout|u2_Display/lt74_31  (
    .a({1'b0,\u2_Display/n2173 }),
    .b(2'b10),
    .fci(\u2_Display/lt74_c31 ),
    .f({\u2_Display/n2205 ,open_n65149}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_0|u2_Display/lt75_cin  (
    .a({\u2_Display/n2239 ,1'b0}),
    .b({1'b0,open_n65155}),
    .fco(\u2_Display/lt75_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_10|u2_Display/lt75_9  (
    .a({\u2_Display/n2229 ,\u2_Display/n2230 }),
    .b(2'b11),
    .fci(\u2_Display/lt75_c9 ),
    .fco(\u2_Display/lt75_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_12|u2_Display/lt75_11  (
    .a({\u2_Display/n2227 ,\u2_Display/n2228 }),
    .b(2'b01),
    .fci(\u2_Display/lt75_c11 ),
    .fco(\u2_Display/lt75_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_14|u2_Display/lt75_13  (
    .a({\u2_Display/n2225 ,\u2_Display/n2226 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c13 ),
    .fco(\u2_Display/lt75_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_16|u2_Display/lt75_15  (
    .a({\u2_Display/n2223 ,\u2_Display/n2224 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c15 ),
    .fco(\u2_Display/lt75_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_18|u2_Display/lt75_17  (
    .a({\u2_Display/n2221 ,\u2_Display/n2222 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c17 ),
    .fco(\u2_Display/lt75_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_20|u2_Display/lt75_19  (
    .a({\u2_Display/n2219 ,\u2_Display/n2220 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c19 ),
    .fco(\u2_Display/lt75_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_22|u2_Display/lt75_21  (
    .a({\u2_Display/n2217 ,\u2_Display/n2218 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c21 ),
    .fco(\u2_Display/lt75_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_24|u2_Display/lt75_23  (
    .a({\u2_Display/n2215 ,\u2_Display/n2216 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c23 ),
    .fco(\u2_Display/lt75_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_26|u2_Display/lt75_25  (
    .a({\u2_Display/n2213 ,\u2_Display/n2214 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c25 ),
    .fco(\u2_Display/lt75_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_28|u2_Display/lt75_27  (
    .a({\u2_Display/n2211 ,\u2_Display/n2212 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c27 ),
    .fco(\u2_Display/lt75_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_2|u2_Display/lt75_1  (
    .a({\u2_Display/n2237 ,\u2_Display/n2238 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c1 ),
    .fco(\u2_Display/lt75_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_30|u2_Display/lt75_29  (
    .a({\u2_Display/n2209 ,\u2_Display/n2210 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c29 ),
    .fco(\u2_Display/lt75_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_4|u2_Display/lt75_3  (
    .a({\u2_Display/n2235 ,\u2_Display/n2236 }),
    .b(2'b10),
    .fci(\u2_Display/lt75_c3 ),
    .fco(\u2_Display/lt75_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_6|u2_Display/lt75_5  (
    .a({\u2_Display/n2233 ,\u2_Display/n2234 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c5 ),
    .fco(\u2_Display/lt75_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_8|u2_Display/lt75_7  (
    .a({\u2_Display/n2231 ,\u2_Display/n2232 }),
    .b(2'b00),
    .fci(\u2_Display/lt75_c7 ),
    .fco(\u2_Display/lt75_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt75_0|u2_Display/lt75_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt75_cout|u2_Display/lt75_31  (
    .a({1'b0,\u2_Display/n2208 }),
    .b(2'b10),
    .fci(\u2_Display/lt75_c31 ),
    .f({\u2_Display/n2240 ,open_n65559}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_0|u2_Display/lt76_cin  (
    .a({\u2_Display/n2274 ,1'b0}),
    .b({1'b0,open_n65565}),
    .fco(\u2_Display/lt76_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_10|u2_Display/lt76_9  (
    .a({\u2_Display/n2264 ,\u2_Display/n2265 }),
    .b(2'b11),
    .fci(\u2_Display/lt76_c9 ),
    .fco(\u2_Display/lt76_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_12|u2_Display/lt76_11  (
    .a({\u2_Display/n2262 ,\u2_Display/n2263 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c11 ),
    .fco(\u2_Display/lt76_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_14|u2_Display/lt76_13  (
    .a({\u2_Display/n2260 ,\u2_Display/n2261 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c13 ),
    .fco(\u2_Display/lt76_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_16|u2_Display/lt76_15  (
    .a({\u2_Display/n2258 ,\u2_Display/n2259 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c15 ),
    .fco(\u2_Display/lt76_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_18|u2_Display/lt76_17  (
    .a({\u2_Display/n2256 ,\u2_Display/n2257 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c17 ),
    .fco(\u2_Display/lt76_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_20|u2_Display/lt76_19  (
    .a({\u2_Display/n2254 ,\u2_Display/n2255 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c19 ),
    .fco(\u2_Display/lt76_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_22|u2_Display/lt76_21  (
    .a({\u2_Display/n2252 ,\u2_Display/n2253 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c21 ),
    .fco(\u2_Display/lt76_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_24|u2_Display/lt76_23  (
    .a({\u2_Display/n2250 ,\u2_Display/n2251 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c23 ),
    .fco(\u2_Display/lt76_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_26|u2_Display/lt76_25  (
    .a({\u2_Display/n2248 ,\u2_Display/n2249 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c25 ),
    .fco(\u2_Display/lt76_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_28|u2_Display/lt76_27  (
    .a({\u2_Display/n2246 ,\u2_Display/n2247 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c27 ),
    .fco(\u2_Display/lt76_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_2|u2_Display/lt76_1  (
    .a({\u2_Display/n2272 ,\u2_Display/n2273 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c1 ),
    .fco(\u2_Display/lt76_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_30|u2_Display/lt76_29  (
    .a({\u2_Display/n2244 ,\u2_Display/n2245 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c29 ),
    .fco(\u2_Display/lt76_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_4|u2_Display/lt76_3  (
    .a({\u2_Display/n2270 ,\u2_Display/n2271 }),
    .b(2'b01),
    .fci(\u2_Display/lt76_c3 ),
    .fco(\u2_Display/lt76_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_6|u2_Display/lt76_5  (
    .a({\u2_Display/n2268 ,\u2_Display/n2269 }),
    .b(2'b00),
    .fci(\u2_Display/lt76_c5 ),
    .fco(\u2_Display/lt76_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_8|u2_Display/lt76_7  (
    .a({\u2_Display/n2266 ,\u2_Display/n2267 }),
    .b(2'b10),
    .fci(\u2_Display/lt76_c7 ),
    .fco(\u2_Display/lt76_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt76_0|u2_Display/lt76_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt76_cout|u2_Display/lt76_31  (
    .a({1'b0,\u2_Display/n2243 }),
    .b(2'b10),
    .fci(\u2_Display/lt76_c31 ),
    .f({\u2_Display/n2275 ,open_n65969}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_0|u2_Display/lt77_cin  (
    .a({\u2_Display/n2309 ,1'b0}),
    .b({1'b0,open_n65975}),
    .fco(\u2_Display/lt77_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_10|u2_Display/lt77_9  (
    .a({\u2_Display/n2299 ,\u2_Display/n2300 }),
    .b(2'b01),
    .fci(\u2_Display/lt77_c9 ),
    .fco(\u2_Display/lt77_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_12|u2_Display/lt77_11  (
    .a({\u2_Display/n2297 ,\u2_Display/n2298 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c11 ),
    .fco(\u2_Display/lt77_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_14|u2_Display/lt77_13  (
    .a({\u2_Display/n2295 ,\u2_Display/n2296 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c13 ),
    .fco(\u2_Display/lt77_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_16|u2_Display/lt77_15  (
    .a({\u2_Display/n2293 ,\u2_Display/n2294 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c15 ),
    .fco(\u2_Display/lt77_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_18|u2_Display/lt77_17  (
    .a({\u2_Display/n2291 ,\u2_Display/n2292 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c17 ),
    .fco(\u2_Display/lt77_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_20|u2_Display/lt77_19  (
    .a({\u2_Display/n2289 ,\u2_Display/n2290 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c19 ),
    .fco(\u2_Display/lt77_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_22|u2_Display/lt77_21  (
    .a({\u2_Display/n2287 ,\u2_Display/n2288 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c21 ),
    .fco(\u2_Display/lt77_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_24|u2_Display/lt77_23  (
    .a({\u2_Display/n2285 ,\u2_Display/n2286 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c23 ),
    .fco(\u2_Display/lt77_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_26|u2_Display/lt77_25  (
    .a({\u2_Display/n2283 ,\u2_Display/n2284 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c25 ),
    .fco(\u2_Display/lt77_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_28|u2_Display/lt77_27  (
    .a({\u2_Display/n2281 ,\u2_Display/n2282 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c27 ),
    .fco(\u2_Display/lt77_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_2|u2_Display/lt77_1  (
    .a({\u2_Display/n2307 ,\u2_Display/n2308 }),
    .b(2'b10),
    .fci(\u2_Display/lt77_c1 ),
    .fco(\u2_Display/lt77_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_30|u2_Display/lt77_29  (
    .a({\u2_Display/n2279 ,\u2_Display/n2280 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c29 ),
    .fco(\u2_Display/lt77_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_4|u2_Display/lt77_3  (
    .a({\u2_Display/n2305 ,\u2_Display/n2306 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c3 ),
    .fco(\u2_Display/lt77_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_6|u2_Display/lt77_5  (
    .a({\u2_Display/n2303 ,\u2_Display/n2304 }),
    .b(2'b00),
    .fci(\u2_Display/lt77_c5 ),
    .fco(\u2_Display/lt77_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_8|u2_Display/lt77_7  (
    .a({\u2_Display/n2301 ,\u2_Display/n2302 }),
    .b(2'b11),
    .fci(\u2_Display/lt77_c7 ),
    .fco(\u2_Display/lt77_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt77_0|u2_Display/lt77_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt77_cout|u2_Display/lt77_31  (
    .a({1'b0,\u2_Display/n2278 }),
    .b(2'b10),
    .fci(\u2_Display/lt77_c31 ),
    .f({\u2_Display/n2310 ,open_n66379}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_0|u2_Display/lt7_2_cin  (
    .a({\u2_Display/n102 [0],1'b0}),
    .b({lcd_ypos[0],open_n66385}),
    .fco(\u2_Display/lt7_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_10|u2_Display/lt7_2_9  (
    .a({\u2_Display/n102 [31],\u2_Display/n102 [9]}),
    .b(lcd_ypos[10:9]),
    .fci(\u2_Display/lt7_2_c9 ),
    .fco(\u2_Display/lt7_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_12|u2_Display/lt7_2_11  (
    .a({\u2_Display/n102 [31],\u2_Display/n102 [31]}),
    .b({1'b0,lcd_ypos[11]}),
    .fci(\u2_Display/lt7_2_c11 ),
    .fco(\u2_Display/lt7_2_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_2|u2_Display/lt7_2_1  (
    .a(\u2_Display/n102 [2:1]),
    .b(lcd_ypos[2:1]),
    .fci(\u2_Display/lt7_2_c1 ),
    .fco(\u2_Display/lt7_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_4|u2_Display/lt7_2_3  (
    .a(\u2_Display/n102 [4:3]),
    .b(lcd_ypos[4:3]),
    .fci(\u2_Display/lt7_2_c3 ),
    .fco(\u2_Display/lt7_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_6|u2_Display/lt7_2_5  (
    .a(\u2_Display/n102 [6:5]),
    .b(lcd_ypos[6:5]),
    .fci(\u2_Display/lt7_2_c5 ),
    .fco(\u2_Display/lt7_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_8|u2_Display/lt7_2_7  (
    .a(\u2_Display/n102 [8:7]),
    .b(lcd_ypos[8:7]),
    .fci(\u2_Display/lt7_2_c7 ),
    .fco(\u2_Display/lt7_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt7_2_0|u2_Display/lt7_2_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt7_2_cout_al_u5062  (
    .a({open_n66555,1'b0}),
    .b({open_n66556,1'b1}),
    .fci(\u2_Display/lt7_2_c13 ),
    .f({open_n66575,\u2_Display/n103 }));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_0|u2_Display/lt88_cin  (
    .a({\u2_Display/counta [0],1'b0}),
    .b({1'b0,open_n66581}),
    .fco(\u2_Display/lt88_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_10|u2_Display/lt88_9  (
    .a(\u2_Display/counta [10:9]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c9 ),
    .fco(\u2_Display/lt88_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_12|u2_Display/lt88_11  (
    .a(\u2_Display/counta [12:11]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c11 ),
    .fco(\u2_Display/lt88_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_14|u2_Display/lt88_13  (
    .a(\u2_Display/counta [14:13]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c13 ),
    .fco(\u2_Display/lt88_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_16|u2_Display/lt88_15  (
    .a(\u2_Display/counta [16:15]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c15 ),
    .fco(\u2_Display/lt88_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_18|u2_Display/lt88_17  (
    .a(\u2_Display/counta [18:17]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c17 ),
    .fco(\u2_Display/lt88_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_20|u2_Display/lt88_19  (
    .a(\u2_Display/counta [20:19]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c19 ),
    .fco(\u2_Display/lt88_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_22|u2_Display/lt88_21  (
    .a(\u2_Display/counta [22:21]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c21 ),
    .fco(\u2_Display/lt88_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_24|u2_Display/lt88_23  (
    .a(\u2_Display/counta [24:23]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c23 ),
    .fco(\u2_Display/lt88_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_26|u2_Display/lt88_25  (
    .a(\u2_Display/counta [26:25]),
    .b(2'b11),
    .fci(\u2_Display/lt88_c25 ),
    .fco(\u2_Display/lt88_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_28|u2_Display/lt88_27  (
    .a(\u2_Display/counta [28:27]),
    .b(2'b10),
    .fci(\u2_Display/lt88_c27 ),
    .fco(\u2_Display/lt88_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_2|u2_Display/lt88_1  (
    .a(\u2_Display/counta [2:1]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c1 ),
    .fco(\u2_Display/lt88_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_30|u2_Display/lt88_29  (
    .a(\u2_Display/counta [30:29]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c29 ),
    .fco(\u2_Display/lt88_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_4|u2_Display/lt88_3  (
    .a(\u2_Display/counta [4:3]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c3 ),
    .fco(\u2_Display/lt88_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_6|u2_Display/lt88_5  (
    .a(\u2_Display/counta [6:5]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c5 ),
    .fco(\u2_Display/lt88_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_8|u2_Display/lt88_7  (
    .a(\u2_Display/counta [8:7]),
    .b(2'b00),
    .fci(\u2_Display/lt88_c7 ),
    .fco(\u2_Display/lt88_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt88_0|u2_Display/lt88_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt88_cout|u2_Display/lt88_31  (
    .a({1'b0,\u2_Display/counta [31]}),
    .b(2'b11),
    .fci(\u2_Display/lt88_c31 ),
    .f({\u2_Display/n2663 ,open_n66985}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_0|u2_Display/lt89_cin  (
    .a({\u2_Display/n2697 ,1'b0}),
    .b({1'b0,open_n66991}),
    .fco(\u2_Display/lt89_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_10|u2_Display/lt89_9  (
    .a({\u2_Display/n2687 ,\u2_Display/n2688 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c9 ),
    .fco(\u2_Display/lt89_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_12|u2_Display/lt89_11  (
    .a({\u2_Display/n2685 ,\u2_Display/n2686 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c11 ),
    .fco(\u2_Display/lt89_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_14|u2_Display/lt89_13  (
    .a({\u2_Display/n2683 ,\u2_Display/n2684 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c13 ),
    .fco(\u2_Display/lt89_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_16|u2_Display/lt89_15  (
    .a({\u2_Display/n2681 ,\u2_Display/n2682 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c15 ),
    .fco(\u2_Display/lt89_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_18|u2_Display/lt89_17  (
    .a({\u2_Display/n2679 ,\u2_Display/n2680 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c17 ),
    .fco(\u2_Display/lt89_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_20|u2_Display/lt89_19  (
    .a({\u2_Display/n2677 ,\u2_Display/n2678 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c19 ),
    .fco(\u2_Display/lt89_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_22|u2_Display/lt89_21  (
    .a({\u2_Display/n2675 ,\u2_Display/n2676 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c21 ),
    .fco(\u2_Display/lt89_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_24|u2_Display/lt89_23  (
    .a({\u2_Display/n2673 ,\u2_Display/n2674 }),
    .b(2'b10),
    .fci(\u2_Display/lt89_c23 ),
    .fco(\u2_Display/lt89_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_26|u2_Display/lt89_25  (
    .a({\u2_Display/n2671 ,\u2_Display/n2672 }),
    .b(2'b01),
    .fci(\u2_Display/lt89_c25 ),
    .fco(\u2_Display/lt89_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_28|u2_Display/lt89_27  (
    .a({\u2_Display/n2669 ,\u2_Display/n2670 }),
    .b(2'b01),
    .fci(\u2_Display/lt89_c27 ),
    .fco(\u2_Display/lt89_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_2|u2_Display/lt89_1  (
    .a({\u2_Display/n2695 ,\u2_Display/n2696 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c1 ),
    .fco(\u2_Display/lt89_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_30|u2_Display/lt89_29  (
    .a({\u2_Display/n2667 ,\u2_Display/n2668 }),
    .b(2'b10),
    .fci(\u2_Display/lt89_c29 ),
    .fco(\u2_Display/lt89_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_4|u2_Display/lt89_3  (
    .a({\u2_Display/n2693 ,\u2_Display/n2694 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c3 ),
    .fco(\u2_Display/lt89_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_6|u2_Display/lt89_5  (
    .a({\u2_Display/n2691 ,\u2_Display/n2692 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c5 ),
    .fco(\u2_Display/lt89_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_8|u2_Display/lt89_7  (
    .a({\u2_Display/n2689 ,\u2_Display/n2690 }),
    .b(2'b00),
    .fci(\u2_Display/lt89_c7 ),
    .fco(\u2_Display/lt89_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt89_0|u2_Display/lt89_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt89_cout|u2_Display/lt89_31  (
    .a({1'b0,\u2_Display/n2666 }),
    .b(2'b10),
    .fci(\u2_Display/lt89_c31 ),
    .f({\u2_Display/n2698 ,open_n67395}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_0|u2_Display/lt8_2_cin  (
    .a({lcd_xpos[0],1'b0}),
    .b({\u2_Display/j [0],open_n67401}),
    .fco(\u2_Display/lt8_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_10|u2_Display/lt8_2_9  (
    .a(lcd_xpos[10:9]),
    .b({\u2_Display/add6_2_co ,\u2_Display/n135 [2]}),
    .fci(\u2_Display/lt8_2_c9 ),
    .fco(\u2_Display/lt8_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_2|u2_Display/lt8_2_1  (
    .a(lcd_xpos[2:1]),
    .b(\u2_Display/j [2:1]),
    .fci(\u2_Display/lt8_2_c1 ),
    .fco(\u2_Display/lt8_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_4|u2_Display/lt8_2_3  (
    .a(lcd_xpos[4:3]),
    .b(\u2_Display/j [4:3]),
    .fci(\u2_Display/lt8_2_c3 ),
    .fco(\u2_Display/lt8_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_6|u2_Display/lt8_2_5  (
    .a(lcd_xpos[6:5]),
    .b(\u2_Display/j [6:5]),
    .fci(\u2_Display/lt8_2_c5 ),
    .fco(\u2_Display/lt8_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_8|u2_Display/lt8_2_7  (
    .a(lcd_xpos[8:7]),
    .b(\u2_Display/n135 [1:0]),
    .fci(\u2_Display/lt8_2_c7 ),
    .fco(\u2_Display/lt8_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt8_2_0|u2_Display/lt8_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt8_2_cout|u2_Display/lt8_2_11  (
    .a({1'b0,lcd_xpos[11]}),
    .b(2'b10),
    .fci(\u2_Display/lt8_2_c11 ),
    .f({\u2_Display/n136 ,open_n67565}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_0|u2_Display/lt90_cin  (
    .a({\u2_Display/n2732 ,1'b0}),
    .b({1'b0,open_n67571}),
    .fco(\u2_Display/lt90_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_10|u2_Display/lt90_9  (
    .a({\u2_Display/n2722 ,\u2_Display/n2723 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c9 ),
    .fco(\u2_Display/lt90_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_12|u2_Display/lt90_11  (
    .a({\u2_Display/n2720 ,\u2_Display/n2721 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c11 ),
    .fco(\u2_Display/lt90_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_14|u2_Display/lt90_13  (
    .a({\u2_Display/n2718 ,\u2_Display/n2719 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c13 ),
    .fco(\u2_Display/lt90_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_16|u2_Display/lt90_15  (
    .a({\u2_Display/n2716 ,\u2_Display/n2717 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c15 ),
    .fco(\u2_Display/lt90_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_18|u2_Display/lt90_17  (
    .a({\u2_Display/n2714 ,\u2_Display/n2715 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c17 ),
    .fco(\u2_Display/lt90_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_20|u2_Display/lt90_19  (
    .a({\u2_Display/n2712 ,\u2_Display/n2713 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c19 ),
    .fco(\u2_Display/lt90_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_22|u2_Display/lt90_21  (
    .a({\u2_Display/n2710 ,\u2_Display/n2711 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c21 ),
    .fco(\u2_Display/lt90_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_24|u2_Display/lt90_23  (
    .a({\u2_Display/n2708 ,\u2_Display/n2709 }),
    .b(2'b11),
    .fci(\u2_Display/lt90_c23 ),
    .fco(\u2_Display/lt90_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_26|u2_Display/lt90_25  (
    .a({\u2_Display/n2706 ,\u2_Display/n2707 }),
    .b(2'b10),
    .fci(\u2_Display/lt90_c25 ),
    .fco(\u2_Display/lt90_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_28|u2_Display/lt90_27  (
    .a({\u2_Display/n2704 ,\u2_Display/n2705 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c27 ),
    .fco(\u2_Display/lt90_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_2|u2_Display/lt90_1  (
    .a({\u2_Display/n2730 ,\u2_Display/n2731 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c1 ),
    .fco(\u2_Display/lt90_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_30|u2_Display/lt90_29  (
    .a({\u2_Display/n2702 ,\u2_Display/n2703 }),
    .b(2'b01),
    .fci(\u2_Display/lt90_c29 ),
    .fco(\u2_Display/lt90_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_4|u2_Display/lt90_3  (
    .a({\u2_Display/n2728 ,\u2_Display/n2729 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c3 ),
    .fco(\u2_Display/lt90_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_6|u2_Display/lt90_5  (
    .a({\u2_Display/n2726 ,\u2_Display/n2727 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c5 ),
    .fco(\u2_Display/lt90_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_8|u2_Display/lt90_7  (
    .a({\u2_Display/n2724 ,\u2_Display/n2725 }),
    .b(2'b00),
    .fci(\u2_Display/lt90_c7 ),
    .fco(\u2_Display/lt90_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt90_0|u2_Display/lt90_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt90_cout|u2_Display/lt90_31  (
    .a({1'b0,\u2_Display/n2701 }),
    .b(2'b10),
    .fci(\u2_Display/lt90_c31 ),
    .f({\u2_Display/n2733 ,open_n67975}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_0|u2_Display/lt91_cin  (
    .a({\u2_Display/n2767 ,1'b0}),
    .b({1'b0,open_n67981}),
    .fco(\u2_Display/lt91_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_10|u2_Display/lt91_9  (
    .a({\u2_Display/n2757 ,\u2_Display/n2758 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c9 ),
    .fco(\u2_Display/lt91_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_12|u2_Display/lt91_11  (
    .a({\u2_Display/n2755 ,\u2_Display/n2756 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c11 ),
    .fco(\u2_Display/lt91_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_14|u2_Display/lt91_13  (
    .a({\u2_Display/n2753 ,\u2_Display/n2754 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c13 ),
    .fco(\u2_Display/lt91_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_16|u2_Display/lt91_15  (
    .a({\u2_Display/n2751 ,\u2_Display/n2752 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c15 ),
    .fco(\u2_Display/lt91_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_18|u2_Display/lt91_17  (
    .a({\u2_Display/n2749 ,\u2_Display/n2750 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c17 ),
    .fco(\u2_Display/lt91_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_20|u2_Display/lt91_19  (
    .a({\u2_Display/n2747 ,\u2_Display/n2748 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c19 ),
    .fco(\u2_Display/lt91_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_22|u2_Display/lt91_21  (
    .a({\u2_Display/n2745 ,\u2_Display/n2746 }),
    .b(2'b10),
    .fci(\u2_Display/lt91_c21 ),
    .fco(\u2_Display/lt91_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_24|u2_Display/lt91_23  (
    .a({\u2_Display/n2743 ,\u2_Display/n2744 }),
    .b(2'b01),
    .fci(\u2_Display/lt91_c23 ),
    .fco(\u2_Display/lt91_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_26|u2_Display/lt91_25  (
    .a({\u2_Display/n2741 ,\u2_Display/n2742 }),
    .b(2'b01),
    .fci(\u2_Display/lt91_c25 ),
    .fco(\u2_Display/lt91_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_28|u2_Display/lt91_27  (
    .a({\u2_Display/n2739 ,\u2_Display/n2740 }),
    .b(2'b10),
    .fci(\u2_Display/lt91_c27 ),
    .fco(\u2_Display/lt91_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_2|u2_Display/lt91_1  (
    .a({\u2_Display/n2765 ,\u2_Display/n2766 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c1 ),
    .fco(\u2_Display/lt91_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_30|u2_Display/lt91_29  (
    .a({\u2_Display/n2737 ,\u2_Display/n2738 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c29 ),
    .fco(\u2_Display/lt91_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_4|u2_Display/lt91_3  (
    .a({\u2_Display/n2763 ,\u2_Display/n2764 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c3 ),
    .fco(\u2_Display/lt91_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_6|u2_Display/lt91_5  (
    .a({\u2_Display/n2761 ,\u2_Display/n2762 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c5 ),
    .fco(\u2_Display/lt91_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_8|u2_Display/lt91_7  (
    .a({\u2_Display/n2759 ,\u2_Display/n2760 }),
    .b(2'b00),
    .fci(\u2_Display/lt91_c7 ),
    .fco(\u2_Display/lt91_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt91_0|u2_Display/lt91_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt91_cout|u2_Display/lt91_31  (
    .a({1'b0,\u2_Display/n2736 }),
    .b(2'b10),
    .fci(\u2_Display/lt91_c31 ),
    .f({\u2_Display/n2768 ,open_n68385}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_0|u2_Display/lt92_cin  (
    .a({\u2_Display/n2802 ,1'b0}),
    .b({1'b0,open_n68391}),
    .fco(\u2_Display/lt92_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_10|u2_Display/lt92_9  (
    .a({\u2_Display/n2792 ,\u2_Display/n2793 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c9 ),
    .fco(\u2_Display/lt92_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_12|u2_Display/lt92_11  (
    .a({\u2_Display/n2790 ,\u2_Display/n2791 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c11 ),
    .fco(\u2_Display/lt92_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_14|u2_Display/lt92_13  (
    .a({\u2_Display/n2788 ,\u2_Display/n2789 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c13 ),
    .fco(\u2_Display/lt92_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_16|u2_Display/lt92_15  (
    .a({\u2_Display/n2786 ,\u2_Display/n2787 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c15 ),
    .fco(\u2_Display/lt92_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_18|u2_Display/lt92_17  (
    .a({\u2_Display/n2784 ,\u2_Display/n2785 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c17 ),
    .fco(\u2_Display/lt92_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_20|u2_Display/lt92_19  (
    .a({\u2_Display/n2782 ,\u2_Display/n2783 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c19 ),
    .fco(\u2_Display/lt92_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_22|u2_Display/lt92_21  (
    .a({\u2_Display/n2780 ,\u2_Display/n2781 }),
    .b(2'b11),
    .fci(\u2_Display/lt92_c21 ),
    .fco(\u2_Display/lt92_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_24|u2_Display/lt92_23  (
    .a({\u2_Display/n2778 ,\u2_Display/n2779 }),
    .b(2'b10),
    .fci(\u2_Display/lt92_c23 ),
    .fco(\u2_Display/lt92_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_26|u2_Display/lt92_25  (
    .a({\u2_Display/n2776 ,\u2_Display/n2777 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c25 ),
    .fco(\u2_Display/lt92_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_28|u2_Display/lt92_27  (
    .a({\u2_Display/n2774 ,\u2_Display/n2775 }),
    .b(2'b01),
    .fci(\u2_Display/lt92_c27 ),
    .fco(\u2_Display/lt92_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_2|u2_Display/lt92_1  (
    .a({\u2_Display/n2800 ,\u2_Display/n2801 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c1 ),
    .fco(\u2_Display/lt92_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_30|u2_Display/lt92_29  (
    .a({\u2_Display/n2772 ,\u2_Display/n2773 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c29 ),
    .fco(\u2_Display/lt92_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_4|u2_Display/lt92_3  (
    .a({\u2_Display/n2798 ,\u2_Display/n2799 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c3 ),
    .fco(\u2_Display/lt92_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_6|u2_Display/lt92_5  (
    .a({\u2_Display/n2796 ,\u2_Display/n2797 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c5 ),
    .fco(\u2_Display/lt92_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_8|u2_Display/lt92_7  (
    .a({\u2_Display/n2794 ,\u2_Display/n2795 }),
    .b(2'b00),
    .fci(\u2_Display/lt92_c7 ),
    .fco(\u2_Display/lt92_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt92_0|u2_Display/lt92_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt92_cout|u2_Display/lt92_31  (
    .a({1'b0,\u2_Display/n2771 }),
    .b(2'b10),
    .fci(\u2_Display/lt92_c31 ),
    .f({\u2_Display/n2803 ,open_n68795}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_0|u2_Display/lt93_cin  (
    .a({\u2_Display/n2837 ,1'b0}),
    .b({1'b0,open_n68801}),
    .fco(\u2_Display/lt93_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_10|u2_Display/lt93_9  (
    .a({\u2_Display/n2827 ,\u2_Display/n2828 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c9 ),
    .fco(\u2_Display/lt93_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_12|u2_Display/lt93_11  (
    .a({\u2_Display/n2825 ,\u2_Display/n2826 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c11 ),
    .fco(\u2_Display/lt93_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_14|u2_Display/lt93_13  (
    .a({\u2_Display/n2823 ,\u2_Display/n2824 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c13 ),
    .fco(\u2_Display/lt93_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_16|u2_Display/lt93_15  (
    .a({\u2_Display/n2821 ,\u2_Display/n2822 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c15 ),
    .fco(\u2_Display/lt93_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_18|u2_Display/lt93_17  (
    .a({\u2_Display/n2819 ,\u2_Display/n2820 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c17 ),
    .fco(\u2_Display/lt93_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_20|u2_Display/lt93_19  (
    .a({\u2_Display/n2817 ,\u2_Display/n2818 }),
    .b(2'b10),
    .fci(\u2_Display/lt93_c19 ),
    .fco(\u2_Display/lt93_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_22|u2_Display/lt93_21  (
    .a({\u2_Display/n2815 ,\u2_Display/n2816 }),
    .b(2'b01),
    .fci(\u2_Display/lt93_c21 ),
    .fco(\u2_Display/lt93_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_24|u2_Display/lt93_23  (
    .a({\u2_Display/n2813 ,\u2_Display/n2814 }),
    .b(2'b01),
    .fci(\u2_Display/lt93_c23 ),
    .fco(\u2_Display/lt93_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_26|u2_Display/lt93_25  (
    .a({\u2_Display/n2811 ,\u2_Display/n2812 }),
    .b(2'b10),
    .fci(\u2_Display/lt93_c25 ),
    .fco(\u2_Display/lt93_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_28|u2_Display/lt93_27  (
    .a({\u2_Display/n2809 ,\u2_Display/n2810 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c27 ),
    .fco(\u2_Display/lt93_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_2|u2_Display/lt93_1  (
    .a({\u2_Display/n2835 ,\u2_Display/n2836 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c1 ),
    .fco(\u2_Display/lt93_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_30|u2_Display/lt93_29  (
    .a({\u2_Display/n2807 ,\u2_Display/n2808 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c29 ),
    .fco(\u2_Display/lt93_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_4|u2_Display/lt93_3  (
    .a({\u2_Display/n2833 ,\u2_Display/n2834 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c3 ),
    .fco(\u2_Display/lt93_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_6|u2_Display/lt93_5  (
    .a({\u2_Display/n2831 ,\u2_Display/n2832 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c5 ),
    .fco(\u2_Display/lt93_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_8|u2_Display/lt93_7  (
    .a({\u2_Display/n2829 ,\u2_Display/n2830 }),
    .b(2'b00),
    .fci(\u2_Display/lt93_c7 ),
    .fco(\u2_Display/lt93_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt93_0|u2_Display/lt93_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt93_cout|u2_Display/lt93_31  (
    .a({1'b0,\u2_Display/n2806 }),
    .b(2'b10),
    .fci(\u2_Display/lt93_c31 ),
    .f({\u2_Display/n2838 ,open_n69205}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_0|u2_Display/lt94_cin  (
    .a({\u2_Display/n2872 ,1'b0}),
    .b({1'b0,open_n69211}),
    .fco(\u2_Display/lt94_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_10|u2_Display/lt94_9  (
    .a({\u2_Display/n2862 ,\u2_Display/n2863 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c9 ),
    .fco(\u2_Display/lt94_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_12|u2_Display/lt94_11  (
    .a({\u2_Display/n2860 ,\u2_Display/n2861 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c11 ),
    .fco(\u2_Display/lt94_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_14|u2_Display/lt94_13  (
    .a({\u2_Display/n2858 ,\u2_Display/n2859 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c13 ),
    .fco(\u2_Display/lt94_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_16|u2_Display/lt94_15  (
    .a({\u2_Display/n2856 ,\u2_Display/n2857 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c15 ),
    .fco(\u2_Display/lt94_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_18|u2_Display/lt94_17  (
    .a({\u2_Display/n2854 ,\u2_Display/n2855 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c17 ),
    .fco(\u2_Display/lt94_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_20|u2_Display/lt94_19  (
    .a({\u2_Display/n2852 ,\u2_Display/n2853 }),
    .b(2'b11),
    .fci(\u2_Display/lt94_c19 ),
    .fco(\u2_Display/lt94_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_22|u2_Display/lt94_21  (
    .a({\u2_Display/n2850 ,\u2_Display/n2851 }),
    .b(2'b10),
    .fci(\u2_Display/lt94_c21 ),
    .fco(\u2_Display/lt94_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_24|u2_Display/lt94_23  (
    .a({\u2_Display/n2848 ,\u2_Display/n2849 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c23 ),
    .fco(\u2_Display/lt94_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_26|u2_Display/lt94_25  (
    .a({\u2_Display/n2846 ,\u2_Display/n2847 }),
    .b(2'b01),
    .fci(\u2_Display/lt94_c25 ),
    .fco(\u2_Display/lt94_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_28|u2_Display/lt94_27  (
    .a({\u2_Display/n2844 ,\u2_Display/n2845 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c27 ),
    .fco(\u2_Display/lt94_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_2|u2_Display/lt94_1  (
    .a({\u2_Display/n2870 ,\u2_Display/n2871 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c1 ),
    .fco(\u2_Display/lt94_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_30|u2_Display/lt94_29  (
    .a({\u2_Display/n2842 ,\u2_Display/n2843 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c29 ),
    .fco(\u2_Display/lt94_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_4|u2_Display/lt94_3  (
    .a({\u2_Display/n2868 ,\u2_Display/n2869 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c3 ),
    .fco(\u2_Display/lt94_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_6|u2_Display/lt94_5  (
    .a({\u2_Display/n2866 ,\u2_Display/n2867 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c5 ),
    .fco(\u2_Display/lt94_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_8|u2_Display/lt94_7  (
    .a({\u2_Display/n2864 ,\u2_Display/n2865 }),
    .b(2'b00),
    .fci(\u2_Display/lt94_c7 ),
    .fco(\u2_Display/lt94_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt94_0|u2_Display/lt94_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt94_cout|u2_Display/lt94_31  (
    .a({1'b0,\u2_Display/n2841 }),
    .b(2'b10),
    .fci(\u2_Display/lt94_c31 ),
    .f({\u2_Display/n2873 ,open_n69615}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_0|u2_Display/lt95_cin  (
    .a({\u2_Display/n2907 ,1'b0}),
    .b({1'b0,open_n69621}),
    .fco(\u2_Display/lt95_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_10|u2_Display/lt95_9  (
    .a({\u2_Display/n2897 ,\u2_Display/n2898 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c9 ),
    .fco(\u2_Display/lt95_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_12|u2_Display/lt95_11  (
    .a({\u2_Display/n2895 ,\u2_Display/n2896 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c11 ),
    .fco(\u2_Display/lt95_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_14|u2_Display/lt95_13  (
    .a({\u2_Display/n2893 ,\u2_Display/n2894 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c13 ),
    .fco(\u2_Display/lt95_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_16|u2_Display/lt95_15  (
    .a({\u2_Display/n2891 ,\u2_Display/n2892 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c15 ),
    .fco(\u2_Display/lt95_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_18|u2_Display/lt95_17  (
    .a({\u2_Display/n2889 ,\u2_Display/n2890 }),
    .b(2'b10),
    .fci(\u2_Display/lt95_c17 ),
    .fco(\u2_Display/lt95_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_20|u2_Display/lt95_19  (
    .a({\u2_Display/n2887 ,\u2_Display/n2888 }),
    .b(2'b01),
    .fci(\u2_Display/lt95_c19 ),
    .fco(\u2_Display/lt95_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_22|u2_Display/lt95_21  (
    .a({\u2_Display/n2885 ,\u2_Display/n2886 }),
    .b(2'b01),
    .fci(\u2_Display/lt95_c21 ),
    .fco(\u2_Display/lt95_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_24|u2_Display/lt95_23  (
    .a({\u2_Display/n2883 ,\u2_Display/n2884 }),
    .b(2'b10),
    .fci(\u2_Display/lt95_c23 ),
    .fco(\u2_Display/lt95_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_26|u2_Display/lt95_25  (
    .a({\u2_Display/n2881 ,\u2_Display/n2882 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c25 ),
    .fco(\u2_Display/lt95_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_28|u2_Display/lt95_27  (
    .a({\u2_Display/n2879 ,\u2_Display/n2880 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c27 ),
    .fco(\u2_Display/lt95_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_2|u2_Display/lt95_1  (
    .a({\u2_Display/n2905 ,\u2_Display/n2906 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c1 ),
    .fco(\u2_Display/lt95_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_30|u2_Display/lt95_29  (
    .a({\u2_Display/n2877 ,\u2_Display/n2878 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c29 ),
    .fco(\u2_Display/lt95_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_4|u2_Display/lt95_3  (
    .a({\u2_Display/n2903 ,\u2_Display/n2904 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c3 ),
    .fco(\u2_Display/lt95_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_6|u2_Display/lt95_5  (
    .a({\u2_Display/n2901 ,\u2_Display/n2902 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c5 ),
    .fco(\u2_Display/lt95_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_8|u2_Display/lt95_7  (
    .a({\u2_Display/n2899 ,\u2_Display/n2900 }),
    .b(2'b00),
    .fci(\u2_Display/lt95_c7 ),
    .fco(\u2_Display/lt95_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt95_0|u2_Display/lt95_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt95_cout|u2_Display/lt95_31  (
    .a({1'b0,\u2_Display/n2876 }),
    .b(2'b10),
    .fci(\u2_Display/lt95_c31 ),
    .f({\u2_Display/n2908 ,open_n70025}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_0|u2_Display/lt96_cin  (
    .a({\u2_Display/n2942 ,1'b0}),
    .b({1'b0,open_n70031}),
    .fco(\u2_Display/lt96_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_10|u2_Display/lt96_9  (
    .a({\u2_Display/n2932 ,\u2_Display/n2933 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c9 ),
    .fco(\u2_Display/lt96_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_12|u2_Display/lt96_11  (
    .a({\u2_Display/n2930 ,\u2_Display/n2931 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c11 ),
    .fco(\u2_Display/lt96_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_14|u2_Display/lt96_13  (
    .a({\u2_Display/n2928 ,\u2_Display/n2929 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c13 ),
    .fco(\u2_Display/lt96_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_16|u2_Display/lt96_15  (
    .a({\u2_Display/n2926 ,\u2_Display/n2927 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c15 ),
    .fco(\u2_Display/lt96_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_18|u2_Display/lt96_17  (
    .a({\u2_Display/n2924 ,\u2_Display/n2925 }),
    .b(2'b11),
    .fci(\u2_Display/lt96_c17 ),
    .fco(\u2_Display/lt96_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_20|u2_Display/lt96_19  (
    .a({\u2_Display/n2922 ,\u2_Display/n2923 }),
    .b(2'b10),
    .fci(\u2_Display/lt96_c19 ),
    .fco(\u2_Display/lt96_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_22|u2_Display/lt96_21  (
    .a({\u2_Display/n2920 ,\u2_Display/n2921 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c21 ),
    .fco(\u2_Display/lt96_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_24|u2_Display/lt96_23  (
    .a({\u2_Display/n2918 ,\u2_Display/n2919 }),
    .b(2'b01),
    .fci(\u2_Display/lt96_c23 ),
    .fco(\u2_Display/lt96_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_26|u2_Display/lt96_25  (
    .a({\u2_Display/n2916 ,\u2_Display/n2917 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c25 ),
    .fco(\u2_Display/lt96_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_28|u2_Display/lt96_27  (
    .a({\u2_Display/n2914 ,\u2_Display/n2915 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c27 ),
    .fco(\u2_Display/lt96_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_2|u2_Display/lt96_1  (
    .a({\u2_Display/n2940 ,\u2_Display/n2941 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c1 ),
    .fco(\u2_Display/lt96_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_30|u2_Display/lt96_29  (
    .a({\u2_Display/n2912 ,\u2_Display/n2913 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c29 ),
    .fco(\u2_Display/lt96_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_4|u2_Display/lt96_3  (
    .a({\u2_Display/n2938 ,\u2_Display/n2939 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c3 ),
    .fco(\u2_Display/lt96_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_6|u2_Display/lt96_5  (
    .a({\u2_Display/n2936 ,\u2_Display/n2937 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c5 ),
    .fco(\u2_Display/lt96_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_8|u2_Display/lt96_7  (
    .a({\u2_Display/n2934 ,\u2_Display/n2935 }),
    .b(2'b00),
    .fci(\u2_Display/lt96_c7 ),
    .fco(\u2_Display/lt96_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt96_0|u2_Display/lt96_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt96_cout|u2_Display/lt96_31  (
    .a({1'b0,\u2_Display/n2911 }),
    .b(2'b10),
    .fci(\u2_Display/lt96_c31 ),
    .f({\u2_Display/n2943 ,open_n70435}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_0|u2_Display/lt97_cin  (
    .a({\u2_Display/n2977 ,1'b0}),
    .b({1'b0,open_n70441}),
    .fco(\u2_Display/lt97_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_10|u2_Display/lt97_9  (
    .a({\u2_Display/n2967 ,\u2_Display/n2968 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c9 ),
    .fco(\u2_Display/lt97_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_12|u2_Display/lt97_11  (
    .a({\u2_Display/n2965 ,\u2_Display/n2966 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c11 ),
    .fco(\u2_Display/lt97_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_14|u2_Display/lt97_13  (
    .a({\u2_Display/n2963 ,\u2_Display/n2964 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c13 ),
    .fco(\u2_Display/lt97_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_16|u2_Display/lt97_15  (
    .a({\u2_Display/n2961 ,\u2_Display/n2962 }),
    .b(2'b10),
    .fci(\u2_Display/lt97_c15 ),
    .fco(\u2_Display/lt97_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_18|u2_Display/lt97_17  (
    .a({\u2_Display/n2959 ,\u2_Display/n2960 }),
    .b(2'b01),
    .fci(\u2_Display/lt97_c17 ),
    .fco(\u2_Display/lt97_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_20|u2_Display/lt97_19  (
    .a({\u2_Display/n2957 ,\u2_Display/n2958 }),
    .b(2'b01),
    .fci(\u2_Display/lt97_c19 ),
    .fco(\u2_Display/lt97_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_22|u2_Display/lt97_21  (
    .a({\u2_Display/n2955 ,\u2_Display/n2956 }),
    .b(2'b10),
    .fci(\u2_Display/lt97_c21 ),
    .fco(\u2_Display/lt97_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_24|u2_Display/lt97_23  (
    .a({\u2_Display/n2953 ,\u2_Display/n2954 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c23 ),
    .fco(\u2_Display/lt97_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_26|u2_Display/lt97_25  (
    .a({\u2_Display/n2951 ,\u2_Display/n2952 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c25 ),
    .fco(\u2_Display/lt97_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_28|u2_Display/lt97_27  (
    .a({\u2_Display/n2949 ,\u2_Display/n2950 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c27 ),
    .fco(\u2_Display/lt97_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_2|u2_Display/lt97_1  (
    .a({\u2_Display/n2975 ,\u2_Display/n2976 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c1 ),
    .fco(\u2_Display/lt97_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_30|u2_Display/lt97_29  (
    .a({\u2_Display/n2947 ,\u2_Display/n2948 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c29 ),
    .fco(\u2_Display/lt97_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_4|u2_Display/lt97_3  (
    .a({\u2_Display/n2973 ,\u2_Display/n2974 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c3 ),
    .fco(\u2_Display/lt97_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_6|u2_Display/lt97_5  (
    .a({\u2_Display/n2971 ,\u2_Display/n2972 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c5 ),
    .fco(\u2_Display/lt97_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_8|u2_Display/lt97_7  (
    .a({\u2_Display/n2969 ,\u2_Display/n2970 }),
    .b(2'b00),
    .fci(\u2_Display/lt97_c7 ),
    .fco(\u2_Display/lt97_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt97_0|u2_Display/lt97_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt97_cout|u2_Display/lt97_31  (
    .a({1'b0,\u2_Display/n2946 }),
    .b(2'b10),
    .fci(\u2_Display/lt97_c31 ),
    .f({\u2_Display/n2978 ,open_n70845}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_0|u2_Display/lt98_cin  (
    .a({\u2_Display/n3012 ,1'b0}),
    .b({1'b0,open_n70851}),
    .fco(\u2_Display/lt98_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_10|u2_Display/lt98_9  (
    .a({\u2_Display/n3002 ,\u2_Display/n3003 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c9 ),
    .fco(\u2_Display/lt98_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_12|u2_Display/lt98_11  (
    .a({\u2_Display/n3000 ,\u2_Display/n3001 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c11 ),
    .fco(\u2_Display/lt98_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_14|u2_Display/lt98_13  (
    .a({\u2_Display/n2998 ,\u2_Display/n2999 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c13 ),
    .fco(\u2_Display/lt98_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_16|u2_Display/lt98_15  (
    .a({\u2_Display/n2996 ,\u2_Display/n2997 }),
    .b(2'b11),
    .fci(\u2_Display/lt98_c15 ),
    .fco(\u2_Display/lt98_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_18|u2_Display/lt98_17  (
    .a({\u2_Display/n2994 ,\u2_Display/n2995 }),
    .b(2'b10),
    .fci(\u2_Display/lt98_c17 ),
    .fco(\u2_Display/lt98_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_20|u2_Display/lt98_19  (
    .a({\u2_Display/n2992 ,\u2_Display/n2993 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c19 ),
    .fco(\u2_Display/lt98_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_22|u2_Display/lt98_21  (
    .a({\u2_Display/n2990 ,\u2_Display/n2991 }),
    .b(2'b01),
    .fci(\u2_Display/lt98_c21 ),
    .fco(\u2_Display/lt98_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_24|u2_Display/lt98_23  (
    .a({\u2_Display/n2988 ,\u2_Display/n2989 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c23 ),
    .fco(\u2_Display/lt98_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_26|u2_Display/lt98_25  (
    .a({\u2_Display/n2986 ,\u2_Display/n2987 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c25 ),
    .fco(\u2_Display/lt98_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_28|u2_Display/lt98_27  (
    .a({\u2_Display/n2984 ,\u2_Display/n2985 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c27 ),
    .fco(\u2_Display/lt98_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_2|u2_Display/lt98_1  (
    .a({\u2_Display/n3010 ,\u2_Display/n3011 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c1 ),
    .fco(\u2_Display/lt98_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_30|u2_Display/lt98_29  (
    .a({\u2_Display/n2982 ,\u2_Display/n2983 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c29 ),
    .fco(\u2_Display/lt98_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_4|u2_Display/lt98_3  (
    .a({\u2_Display/n3008 ,\u2_Display/n3009 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c3 ),
    .fco(\u2_Display/lt98_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_6|u2_Display/lt98_5  (
    .a({\u2_Display/n3006 ,\u2_Display/n3007 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c5 ),
    .fco(\u2_Display/lt98_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_8|u2_Display/lt98_7  (
    .a({\u2_Display/n3004 ,\u2_Display/n3005 }),
    .b(2'b00),
    .fci(\u2_Display/lt98_c7 ),
    .fco(\u2_Display/lt98_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt98_0|u2_Display/lt98_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt98_cout|u2_Display/lt98_31  (
    .a({1'b0,\u2_Display/n2981 }),
    .b(2'b10),
    .fci(\u2_Display/lt98_c31 ),
    .f({\u2_Display/n3013 ,open_n71255}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_0|u2_Display/lt99_cin  (
    .a({\u2_Display/n3047 ,1'b0}),
    .b({1'b0,open_n71261}),
    .fco(\u2_Display/lt99_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_10|u2_Display/lt99_9  (
    .a({\u2_Display/n3037 ,\u2_Display/n3038 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c9 ),
    .fco(\u2_Display/lt99_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_12|u2_Display/lt99_11  (
    .a({\u2_Display/n3035 ,\u2_Display/n3036 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c11 ),
    .fco(\u2_Display/lt99_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_14|u2_Display/lt99_13  (
    .a({\u2_Display/n3033 ,\u2_Display/n3034 }),
    .b(2'b10),
    .fci(\u2_Display/lt99_c13 ),
    .fco(\u2_Display/lt99_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_16|u2_Display/lt99_15  (
    .a({\u2_Display/n3031 ,\u2_Display/n3032 }),
    .b(2'b01),
    .fci(\u2_Display/lt99_c15 ),
    .fco(\u2_Display/lt99_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_18|u2_Display/lt99_17  (
    .a({\u2_Display/n3029 ,\u2_Display/n3030 }),
    .b(2'b01),
    .fci(\u2_Display/lt99_c17 ),
    .fco(\u2_Display/lt99_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_20|u2_Display/lt99_19  (
    .a({\u2_Display/n3027 ,\u2_Display/n3028 }),
    .b(2'b10),
    .fci(\u2_Display/lt99_c19 ),
    .fco(\u2_Display/lt99_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_22|u2_Display/lt99_21  (
    .a({\u2_Display/n3025 ,\u2_Display/n3026 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c21 ),
    .fco(\u2_Display/lt99_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_24|u2_Display/lt99_23  (
    .a({\u2_Display/n3023 ,\u2_Display/n3024 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c23 ),
    .fco(\u2_Display/lt99_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_26|u2_Display/lt99_25  (
    .a({\u2_Display/n3021 ,\u2_Display/n3022 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c25 ),
    .fco(\u2_Display/lt99_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_28|u2_Display/lt99_27  (
    .a({\u2_Display/n3019 ,\u2_Display/n3020 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c27 ),
    .fco(\u2_Display/lt99_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_2|u2_Display/lt99_1  (
    .a({\u2_Display/n3045 ,\u2_Display/n3046 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c1 ),
    .fco(\u2_Display/lt99_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_30|u2_Display/lt99_29  (
    .a({\u2_Display/n3017 ,\u2_Display/n3018 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c29 ),
    .fco(\u2_Display/lt99_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_4|u2_Display/lt99_3  (
    .a({\u2_Display/n3043 ,\u2_Display/n3044 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c3 ),
    .fco(\u2_Display/lt99_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_6|u2_Display/lt99_5  (
    .a({\u2_Display/n3041 ,\u2_Display/n3042 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c5 ),
    .fco(\u2_Display/lt99_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_8|u2_Display/lt99_7  (
    .a({\u2_Display/n3039 ,\u2_Display/n3040 }),
    .b(2'b00),
    .fci(\u2_Display/lt99_c7 ),
    .fco(\u2_Display/lt99_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt99_0|u2_Display/lt99_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt99_cout|u2_Display/lt99_31  (
    .a({1'b0,\u2_Display/n3016 }),
    .b(2'b10),
    .fci(\u2_Display/lt99_c31 ),
    .f({\u2_Display/n3048 ,open_n71665}));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_0|u2_Display/lt9_2_cin  (
    .a({\u2_Display/n137 [0],1'b0}),
    .b({lcd_xpos[0],open_n71671}),
    .fco(\u2_Display/lt9_2_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_10|u2_Display/lt9_2_9  (
    .a({\u2_Display/n137 [31],\u2_Display/n137 [9]}),
    .b(lcd_xpos[10:9]),
    .fci(\u2_Display/lt9_2_c9 ),
    .fco(\u2_Display/lt9_2_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_12|u2_Display/lt9_2_11  (
    .a({\u2_Display/n137 [31],\u2_Display/n137 [31]}),
    .b({1'b0,lcd_xpos[11]}),
    .fci(\u2_Display/lt9_2_c11 ),
    .fco(\u2_Display/lt9_2_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_2|u2_Display/lt9_2_1  (
    .a(\u2_Display/n137 [2:1]),
    .b(lcd_xpos[2:1]),
    .fci(\u2_Display/lt9_2_c1 ),
    .fco(\u2_Display/lt9_2_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_4|u2_Display/lt9_2_3  (
    .a(\u2_Display/n137 [4:3]),
    .b(lcd_xpos[4:3]),
    .fci(\u2_Display/lt9_2_c3 ),
    .fco(\u2_Display/lt9_2_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_6|u2_Display/lt9_2_5  (
    .a(\u2_Display/n137 [6:5]),
    .b(lcd_xpos[6:5]),
    .fci(\u2_Display/lt9_2_c5 ),
    .fco(\u2_Display/lt9_2_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_8|u2_Display/lt9_2_7  (
    .a(\u2_Display/n137 [8:7]),
    .b(lcd_xpos[8:7]),
    .fci(\u2_Display/lt9_2_c7 ),
    .fco(\u2_Display/lt9_2_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u2_Display/lt9_2_0|u2_Display/lt9_2_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u2_Display/lt9_2_cout_al_u5063  (
    .a({open_n71841,1'b0}),
    .b({open_n71842,1'b1}),
    .fci(\u2_Display/lt9_2_c13 ),
    .f({open_n71861,\u2_Display/n138 }));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b0  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [0]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [0]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b1  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [1]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [1]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b10  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [10]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [10]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b11  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [11]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [11]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b12  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [12]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [12]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b13  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [13]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [13]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b14  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [14]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [14]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b15  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [15]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [15]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b16  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [16]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [16]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b17  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [17]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [17]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b18  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [18]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [18]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b19  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [19]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [19]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b2  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [2]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [2]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b20  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [20]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [20]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b21  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [21]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [21]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b22  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [22]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [22]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b23  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [23]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [23]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b24  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [24]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [24]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b25  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [25]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [25]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b26  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [26]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [26]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b27  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [27]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [27]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b28  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [28]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [28]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b29  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [29]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [29]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b3  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [3]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [3]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b30  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [30]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [30]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b4  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [4]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [4]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b5  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [5]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [5]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b6  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [6]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [6]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b7  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [7]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [7]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b8  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [8]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [8]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u2_Display/reg0_b9  (
    .clk(clk_vga),
    .d(\u2_Display/n37 [9]),
    .sr(\u2_Display/n35 ),
    .q(\u2_Display/n [9]));  // source/rtl/Display.v(61)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u2_Display/reg1_b0  (
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n240 [0]),
    .sr(rst_n_pad),
    .q(lcd_data[23]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b0  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [0]),
    .q(\u2_Display/counta [0]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b1  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [1]),
    .q(\u2_Display/counta [1]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b10  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [10]),
    .q(\u2_Display/counta [10]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b11  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [11]),
    .q(\u2_Display/counta [11]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b12  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [12]),
    .q(\u2_Display/counta [12]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b13  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [13]),
    .q(\u2_Display/counta [13]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b14  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [14]),
    .q(\u2_Display/counta [14]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b15  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [15]),
    .q(\u2_Display/counta [15]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b16  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [16]),
    .q(\u2_Display/counta [16]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b17  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [17]),
    .q(\u2_Display/counta [17]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b18  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [18]),
    .q(\u2_Display/counta [18]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b19  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [19]),
    .q(\u2_Display/counta [19]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b2  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [2]),
    .q(\u2_Display/counta [2]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b20  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [20]),
    .q(\u2_Display/counta [20]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b21  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [21]),
    .q(\u2_Display/counta [21]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b22  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [22]),
    .q(\u2_Display/counta [22]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b23  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [23]),
    .q(\u2_Display/counta [23]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b24  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [24]),
    .q(\u2_Display/counta [24]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b25  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [25]),
    .q(\u2_Display/counta [25]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b26  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [26]),
    .q(\u2_Display/counta [26]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b27  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [27]),
    .q(\u2_Display/counta [27]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b28  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [28]),
    .q(\u2_Display/counta [28]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b29  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [29]),
    .q(\u2_Display/counta [29]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b3  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [3]),
    .q(\u2_Display/counta [3]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b30  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [30]),
    .q(\u2_Display/counta [30]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b31  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [31]),
    .q(\u2_Display/counta [31]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b4  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [4]),
    .q(\u2_Display/counta [4]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b5  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [5]),
    .q(\u2_Display/counta [5]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b6  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [6]),
    .q(\u2_Display/counta [6]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b7  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [7]),
    .q(\u2_Display/counta [7]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b8  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [8]),
    .q(\u2_Display/counta [8]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg2_b9  (
    .ce(\u2_Display/mux21_b0_sel_is_0_o ),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n41 [9]),
    .q(\u2_Display/counta [9]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b0  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [0]),
    .q(\u2_Display/i [0]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b1  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [1]),
    .q(\u2_Display/i [1]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b10  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [10]),
    .q(\u2_Display/i [10]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b2  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [2]),
    .q(\u2_Display/i [2]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b3  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [3]),
    .q(\u2_Display/i [3]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b4  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [4]),
    .q(\u2_Display/i [4]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b5  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [5]),
    .q(\u2_Display/i [5]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b6  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [6]),
    .q(\u2_Display/i [6]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b7  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [7]),
    .q(\u2_Display/i [7]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b8  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [8]),
    .q(\u2_Display/i [8]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg3_b9  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n238 [9]),
    .q(\u2_Display/i [9]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b0  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [0]),
    .q(\u2_Display/j [0]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b1  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [1]),
    .q(\u2_Display/j [1]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b2  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [2]),
    .q(\u2_Display/j [2]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b3  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [3]),
    .q(\u2_Display/j [3]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b4  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [4]),
    .q(\u2_Display/j [4]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b5  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [5]),
    .q(\u2_Display/j [5]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b6  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [6]),
    .q(\u2_Display/j [6]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b7  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [7]),
    .q(\u2_Display/j [7]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b8  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [8]),
    .q(\u2_Display/j [8]));  // source/rtl/Display.v(252)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u2_Display/reg4_b9  (
    .ce(rst_n_pad),
    .clk(\u2_Display/clk1s ),
    .d(\u2_Display/n239 [9]),
    .q(\u2_Display/j [9]));  // source/rtl/Display.v(252)
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub0_2/ucin_al_u5029"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub0_2/u3_al_u5030  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/i [5],\u2_Display/i [3]}),
    .e({\u2_Display/i [6],\u2_Display/i [4]}),
    .fci(\u2_Display/sub0_2/c3 ),
    .f({\u2_Display/n96 [5],\u2_Display/n96 [3]}),
    .fco(\u2_Display/sub0_2/c7 ),
    .fx({\u2_Display/n96 [6],\u2_Display/n96 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub0_2/ucin_al_u5029"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub0_2/u7_al_u5031  (
    .a(2'b11),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/i [9],\u2_Display/i [7]}),
    .e({\u2_Display/i [10],\u2_Display/i [8]}),
    .fci(\u2_Display/sub0_2/c7 ),
    .f({\u2_Display/n96 [9],\u2_Display/n96 [7]}),
    .fco(\u2_Display/sub0_2/c11 ),
    .fx({\u2_Display/n96 [10],\u2_Display/n96 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub0_2/ucin_al_u5029"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub0_2/ucin_al_u5029  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/i [1],1'b1}),
    .e({\u2_Display/i [2],\u2_Display/i [0]}),
    .f({\u2_Display/n96 [1],open_n72005}),
    .fco(\u2_Display/sub0_2/c3 ),
    .fx({\u2_Display/n96 [2],\u2_Display/n96 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub0_2/ucin_al_u5029"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub0_2/ucout_al_u5032  (
    .c(2'b11),
    .fci(\u2_Display/sub0_2/c11 ),
    .f({open_n72032,\u2_Display/n96 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub1_2/ucin_al_u5037"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub1_2/u3_al_u5038  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/j [5],\u2_Display/j [3]}),
    .e({\u2_Display/j [6],\u2_Display/j [4]}),
    .fci(\u2_Display/sub1_2/c3 ),
    .f({\u2_Display/n102 [5],\u2_Display/n102 [3]}),
    .fco(\u2_Display/sub1_2/c7 ),
    .fx({\u2_Display/n102 [6],\u2_Display/n102 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub1_2/ucin_al_u5037"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub1_2/u7_al_u5039  (
    .a(2'b10),
    .b({open_n72056,1'b0}),
    .c(2'b11),
    .d({\u2_Display/j [9],\u2_Display/j [7]}),
    .e({open_n72059,\u2_Display/j [8]}),
    .fci(\u2_Display/sub1_2/c7 ),
    .f({\u2_Display/n102 [9],\u2_Display/n102 [7]}),
    .fx({\u2_Display/n102 [31],\u2_Display/n102 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub1_2/ucin_al_u5037"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub1_2/ucin_al_u5037  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/j [1],1'b1}),
    .e({\u2_Display/j [2],\u2_Display/j [0]}),
    .f({\u2_Display/n102 [1],open_n72094}),
    .fco(\u2_Display/sub1_2/c3 ),
    .fx({\u2_Display/n102 [2],\u2_Display/n102 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub2_2/ucin_al_u5040"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub2_2/u3_al_u5041  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/j [5],\u2_Display/j [3]}),
    .e({\u2_Display/j [6],\u2_Display/j [4]}),
    .fci(\u2_Display/sub2_2/c3 ),
    .f({\u2_Display/n137 [5],\u2_Display/n137 [3]}),
    .fco(\u2_Display/sub2_2/c7 ),
    .fx({\u2_Display/n137 [6],\u2_Display/n137 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub2_2/ucin_al_u5040"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub2_2/u7_al_u5042  (
    .a(2'b11),
    .b({open_n72115,1'b0}),
    .c(2'b11),
    .d({\u2_Display/j [9],\u2_Display/j [7]}),
    .e({open_n72118,\u2_Display/j [8]}),
    .fci(\u2_Display/sub2_2/c7 ),
    .f({\u2_Display/n137 [9],\u2_Display/n137 [7]}),
    .fx({\u2_Display/n137 [31],\u2_Display/n137 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub2_2/ucin_al_u5040"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub2_2/ucin_al_u5040  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/j [1],1'b1}),
    .e({\u2_Display/j [2],\u2_Display/j [0]}),
    .f({\u2_Display/n137 [1],open_n72153}),
    .fco(\u2_Display/sub2_2/c3 ),
    .fx({\u2_Display/n137 [2],\u2_Display/n137 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub3_2/ucin_al_u5033"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub3_2/u3_al_u5034  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/i [5],\u2_Display/i [3]}),
    .e({\u2_Display/i [6],\u2_Display/i [4]}),
    .fci(\u2_Display/sub3_2/c3 ),
    .f({\u2_Display/n143 [5],\u2_Display/n143 [3]}),
    .fco(\u2_Display/sub3_2/c7 ),
    .fx({\u2_Display/n143 [6],\u2_Display/n143 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub3_2/ucin_al_u5033"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub3_2/u7_al_u5035  (
    .a(2'b10),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/i [9],\u2_Display/i [7]}),
    .e({\u2_Display/i [10],\u2_Display/i [8]}),
    .fci(\u2_Display/sub3_2/c7 ),
    .f({\u2_Display/n143 [9],\u2_Display/n143 [7]}),
    .fco(\u2_Display/sub3_2/c11 ),
    .fx({\u2_Display/n143 [10],\u2_Display/n143 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub3_2/ucin_al_u5033"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub3_2/ucin_al_u5033  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({\u2_Display/i [1],1'b1}),
    .e({\u2_Display/i [2],\u2_Display/i [0]}),
    .f({\u2_Display/n143 [1],open_n72209}),
    .fco(\u2_Display/sub3_2/c3 ),
    .fx({\u2_Display/n143 [2],\u2_Display/n143 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2_Display/sub3_2/ucin_al_u5033"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2_Display/sub3_2/ucout_al_u5036  (
    .c(2'b11),
    .fci(\u2_Display/sub3_2/c11 ),
    .f({open_n72236,\u2_Display/n143 [31]}));

endmodule 

